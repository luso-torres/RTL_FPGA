// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Thu Jul 24 12:29:56 2025
//
// Verilog Description of module matrix_inv
//

module matrix_inv (clk, reset, a, b, c, d, a_inv, b_inv, c_inv, 
            d_inv, error) /* synthesis syn_module_defined=1 */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(8[8:18])
    input clk;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[20:23])
    input reset;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[25:30])
    input [15:0]a;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    input [15:0]b;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    input [15:0]c;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    input [15:0]d;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    output [15:0]a_inv;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    output [15:0]b_inv;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    output [15:0]c_inv;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    output [15:0]d_inv;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    output error;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(19[26:31])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[20:23])
    
    wire GND_net, VCC_net, reset_c, a_c_15, a_c_14, a_c_13, a_c_12, 
        a_c_11, a_c_10, a_c_9, a_c_8, a_c_7, a_c_6, a_c_5, a_c_4, 
        a_c_3, a_c_2, a_c_1, a_c_0, b_c_15, b_c_14, b_c_13, b_c_12, 
        b_c_11, b_c_10, b_c_9, b_c_8, b_c_7, b_c_6, b_c_5, b_c_4, 
        b_c_3, b_c_2, b_c_1, b_c_0, c_c_15, c_c_14, c_c_13, c_c_12, 
        c_c_11, c_c_10, c_c_9, c_c_8, c_c_7, c_c_6, c_c_5, c_c_4, 
        c_c_3, c_c_2, c_c_1, c_c_0, d_c_15, d_c_14, d_c_13, d_c_12, 
        d_c_11, d_c_10, d_c_9, d_c_8, d_c_7, d_c_6, d_c_5, d_c_4, 
        d_c_3, d_c_2, d_c_1, d_c_0, a_inv_c_15, a_inv_c_14, a_inv_c_13, 
        a_inv_c_12, a_inv_c_11, a_inv_c_10, a_inv_c_9, a_inv_c_8, 
        a_inv_c_7, a_inv_c_6, a_inv_c_5, a_inv_c_4, a_inv_c_3, a_inv_c_2, 
        a_inv_c_1, a_inv_c_0, b_inv_c_15, b_inv_c_14, b_inv_c_13, 
        b_inv_c_12, b_inv_c_11, b_inv_c_10, b_inv_c_9, b_inv_c_8, 
        b_inv_c_7, b_inv_c_6, b_inv_c_5, b_inv_c_4, b_inv_c_3, b_inv_c_2, 
        b_inv_c_1, b_inv_c_0, c_inv_c_15, c_inv_c_14, c_inv_c_13, 
        c_inv_c_12, c_inv_c_11, c_inv_c_10, c_inv_c_9, c_inv_c_8, 
        c_inv_c_7, c_inv_c_6, c_inv_c_5, c_inv_c_4, c_inv_c_3, c_inv_c_2, 
        c_inv_c_1, c_inv_c_0, d_inv_c_15, d_inv_c_14, d_inv_c_13, 
        d_inv_c_12, d_inv_c_11, d_inv_c_10, d_inv_c_9, d_inv_c_8, 
        d_inv_c_7, d_inv_c_6, d_inv_c_5, d_inv_c_4, d_inv_c_3, d_inv_c_2, 
        d_inv_c_1, d_inv_c_0, error_c;
    wire [31:0]det_q4_28;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(31[34:43])
    wire [15:0]a1_reg;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(32[34:40])
    wire [15:0]b1_reg;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(32[42:48])
    wire [15:0]c1_reg;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(32[50:56])
    wire [15:0]d1_reg;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(32[58:64])
    
    wire det_zero_reg, n10808, n11140, n10817, n11124, n10807, n11139, 
        n10818, n11125, n11138, n11126, n11137, n11127, n11136, 
        n11128;
    wire [15:0]b2_reg;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(36[42:48])
    wire [15:0]c2_reg;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(36[50:56])
    
    wire n11135, n11129, n11134, n11130, n11133, n11131, n11132, 
        n10700, n10701, n10702, n10703, n10704, n10705, n10706, 
        n10707, n10708, det_zero_stage2, n10903, n10535, n10904, 
        n10534, n10905, n10533, n10906, n10532, n10907, n10391, 
        n10390, n10389, n10388, n10387, n10386, n10385, n10384, 
        n10383, n10382, n10381, n10380, n10379, n10378, n10377, 
        n10568, n10567, n10566, error_recip, n10531, n10709, n10710, 
        n10819, n11368, n10530, n11369, n10529, n11370, n10528, 
        n11371, n10376, n10375, n10374, n10711;
    wire [31:0]b_s;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[24:27])
    
    wire n10373, n10372, n10371, n10370, n10369, n10368, n10367, 
        n10366, n10365, n10364, n10363, n10362, n10667, n10666;
    wire [31:0]c_s;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[24:27])
    wire [47:0]prod_a;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[35:41])
    wire [47:0]prod_b;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[35:41])
    
    wire n10712, n10800, n10549;
    wire [47:0]prod_c;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[35:41])
    
    wire n10548, n10806, n10547, n64, n63, n62, n61, n60, n59, 
        n58, n57, n56;
    wire [47:0]prod_d;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[35:41])
    
    wire n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, 
        n45, n44, n43;
    wire [31:0]det_q4_28_31__N_97;
    wire [31:0]det_q4_28_31__N_129;
    wire [31:0]det_q4_28_31__N_65;
    
    wire det_zero_reg_N_162;
    wire [47:0]a_inv_15__N_1;
    wire [47:0]b_inv_15__N_17;
    wire [47:0]c_inv_15__N_33;
    wire [47:0]d_inv_15__N_49;
    
    wire n1412, n1413, n10546, n10527, n10545, n10526, n10544, 
        n10525, n10543, n10524, n10542, n10523, n10541, n10522, 
        n10540, n10521, n10539, n10520, n10538, n10519, n10537, 
        n10518, n10536, n10517, n10361, n10516, n10360, n10515, 
        n10359, n10514, n10358, n10513, n10357, inv_det_31__N_227, 
        n1415, n1414, n1411, n1410, n1416, n1417, n1418, n1419, 
        n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
        n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
        n1436, n1437, n1438, n1439, n1440, n1441, n42, n1444, 
        n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
        n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
        n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
        n1469, n1470, n1471, n1472, n1473, n1474, n1475, n10658, 
        n10657, n10656, n10655, n10654, n10653, n10652, n10651, 
        n10650, n10649, n10648, n10647, n10646, n10645, n10644, 
        n10643, n10642, n10641, n10640, n10639, n10638, n10637, 
        n10636, n10635, n10356, n10355, n10354, n10353, n10352, 
        n10351, n10350, n10349, n10348, n10347, n10346, n10345, 
        n10344, n10343, n10342, n10341, n130, n11307, n128, n11306, 
        n126, n11305, n124, n11304, n122, n11303, n120, n11302, 
        n118, n11301, n116, n11300, n114, n11299, n112, n11298, 
        n110, n11297, n108, n41, n11296, n106, n11295, n104, 
        n11294, n102, n11293, n11260, n11292, n11261, n11291, 
        n11262, n11290, n11263, n11289, n11264, n11288, n11265, 
        n11287, n11266, n11286, n11267, n11268, n11269, n40, n68, 
        n10668, n11259, n10669, n11258, n10670, n11257, n10671, 
        n11256, n10672, n11255, n10673, n11254, n10674, n11253, 
        n10675, n11252, n10676, n11251, n10677, n11250, n10678, 
        n39, n11249, n10679, n11248, n10680, n11247, n10681, n11246, 
        n10682, n11245, n10683, n11244, n10684, n11243, n10685, 
        n11242, n10686, n11241, n10687, n11240, n10688, n11239, 
        n10689, n11238, n10690, n11237, n10691, n11236, n10692, 
        n11235, n10693, n11234, n38, n10694, n11233, n10695, n11232, 
        n10696, n11231, n10697, n11230, n10698, n11229, n10699, 
        n11228, n10512, n11164, n10511, n11165, n10510, n11166, 
        n10509, n11167, n10508, n11168, n10507, n11169, n10506, 
        n11170, n10505, n11171, n10504, n11172, n10503, n37, n1813, 
        n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
        n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
        n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
        n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1846, 
        n36, n11173, n10502, n11174, n10501, n11175, n10500, n11176, 
        n10499, n11177, n10498, n11178, n11179, n11180, n11181, 
        n11182, n11183, n11184, n11185, n11186, n11187, n11188, 
        n11189, n11190, n11191, n11192, n11193, n11194, n11195, 
        n11196, n11197, n11198, n11199, n11200, n11201, n11202, 
        n11203, n11204, n11205, n11206, n11207, n11208, n11209, 
        n11210, n11211, n10497, n11212, n10496, n11213, n10495, 
        n11214, n10494, n11215, n10493, n11216, n10492, n11217, 
        n10491, n11218, n10490, n11219, n10489, n11220, n10488, 
        n10665, n11221, n10487, n11222, n10486, n11223, n10485, 
        n11224, n10484, n11225, n10483, n11226, n10482, n11227, 
        n10340, n10339, n10338, n10337, n10336, n10335, n10334, 
        n10333, n10332, n10331, n10330, n10329, n10328, n10327, 
        n10326, n10634, n10633, n10632, n10664, n10631, n10630, 
        n10629, n10628, n10627, n10626, n10625, n10624, n10623, 
        n10622, n10621, n10620, n10619, n10618, n10617, n10616, 
        n10615, n10614, n10613, n10612, n10611, n10610, n10609, 
        n10608, n10607, n10606, n10605, n10604, n10603, n10602, 
        n10325, n10663, n10324, n10323, n10322, n10321, n10320, 
        n10319, n10318, n10317, n10316, n10315, n10314, n10313, 
        n10312, n10311, n10310, n11100, n11163, n11101, n11162, 
        n11102, n11161, n11103, n11160, n11104, n11159, n11105, 
        n11158, n11106, n11157, n11107, n11156, n10662, n11108, 
        n11155, n11109, n11154, n11110, n11153, n11111, n11152, 
        n11112, n11151, n11113, n11150, n11114, n11149, n11115, 
        n11148, n11116, n11147, n11117, n11146, n11118, n11145, 
        n11119, n11144, n11120, n11143, n11121, n11142, n11122, 
        n11141, n11123, n10661, n10713, n10714, n10715, n10716, 
        n10717, n10718, n10719, n10720, n10721, n10722, n10723, 
        n10724, n10725, n10726, n10727, n10728, n10729, n10730, 
        n10731, n10481, n11004, n10480, n11005, n10479, n11006, 
        n10478, n11007, n10477, n11008, n10476, n11009, n10660, 
        n10475, n11010, n10474, n11011, n10473, n11012, n10472, 
        n11013, n10471, n11014, n10470, n11015, n10469, n11016, 
        n10468, n11017, n10467, n11018, n11019, n11020, n11021, 
        n11022, n11023, n11024, n11025, n11026, n11027, n11028, 
        n11029, n11030, n11031, n35, n2349, n2350, n2351, n2352, 
        n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
        n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, 
        n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
        n2377, n2378, n2379, n2380, n2382, n34, n11032, n11033, 
        n11099, n11098, n11097, n11096, n11095, n11094, n11093, 
        n11092, n11091, n11090, n11089, n11088, n11087, n11086, 
        n11085, n11084, n11083, n11082, n11081, n11080, n11079, 
        n11078, n11077, n11076, n11075, n11074, n11073, n11072, 
        n11071, n11070, n2449, n10659, n11069, n11068, n11034, 
        n11035, n11036, n11037, n11038, n11039, n11040, n11041, 
        n11042, n11043, n11044, n11045, n11046, n11047, n11048, 
        n11049, n11050, n11051, n10466, n11052, n10465, n11053, 
        n10464, n11054, n10463, n11055, n10462, n11056, n10461, 
        n11057, n2516, n10460, n10459, n11058, n10908, n10909, 
        n10926, n10927, n10928, n10929, n10930, n10931, n10932, 
        n10933, n10934, n10935, n10936, n10937, n2583, n10938, 
        n10939, n10458, n11059, n10457, n11060, n10456, n11061, 
        n10455, n11062, n10454, n11063, n10453, n11064, n10452, 
        n11065, n10451, n11066, n10450, n11067, n10309, n10308, 
        n10307, n10306, n10305, n10304, n10303, n10302, n10301, 
        n10300, n10299, n10449, n2617, n2618, n2619, n2620, n2621, 
        n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
        n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
        n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, 
        n2646, n2647, n2648, n2650, n33, n10298, n10297, n10296, 
        n10295, n10294, n10293, n10292, n10291, n10290, n10289, 
        n10288, n10287, n10286, n10285, n10284, n10283, n10282, 
        n10281, n10280, n10279, n10278, n10277, n10276, n10275, 
        n10274, n10273, n10272, n10271, n10270, n10269, n10268, 
        n10267, n10266, n10265, n10264, n10263, n10601, n10600, 
        n10599, n10598, n10597, n10596, n10595, n10594, n10593, 
        n10592, n10591, n10590, n10589, n10588, n10587, n10586, 
        n10585, n10584, n10583, n10582, n10581, n10580, n10579, 
        n10578, n10577, n10576, n10575, n10574, n10573, n10572, 
        n10571, n10570, n10569, n10262, n10261, n10260, n10259, 
        n10258, n10257, n10256, n10255, n10254, n10253, n10252, 
        n10251, n10250, n10249, n10248, n10247, n10940, n11003, 
        n10941, n11002, n10942, n11001, n10943, n11000, n10944, 
        n106_adj_230, n10999, n10945, n10998, n10946, n10997, n10947, 
        n10996, n10948, n10995, n10949, n10994, n10950, n10993, 
        n10951, n10992, n10952, n10991, n10953, n10990, n10954, 
        n10989, n10955, n10988, n10956, n10987, n10957, n10986, 
        n10958, n10985, n10959, n10984, n10960, n10983, n10961, 
        n10982, n10246, n10245, n10244, n10243, n10242, n10241, 
        n10240, n10239, n10238, n10237, n10236, n130_adj_231, n10843, 
        n128_adj_232, n10842, n126_adj_233, n10841, n124_adj_234, 
        n10840, n122_adj_235, n10839, n120_adj_236, n10838, n118_adj_237, 
        n10837, n116_adj_238, n10836, n114_adj_239, n10835, n112_adj_240, 
        n10834, n110_adj_241, n10962, n10981, n10963, n10980, n10964, 
        n10979, n10965, n10978, n10448, n10824, n10966, n10801, 
        n10977, n10967, n10976, n10968, n10975, n10969, n10974, 
        n10970, n10973, n10971, n10972, n10732, n10733, n10734, 
        n10735, n10736, n10737, n10738, n10739, n10740, n10741, 
        n10742, n10743, n10744, n10745, n10746, n10747, n10748, 
        n10749, n10750, n10751, n10752, n10832, n10753, n10833, 
        n108_adj_242, n10754, n3421, n3422, n3423, n3424, n3425, 
        n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
        n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
        n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
        n3450, n3451, n3452, n3454, n10755, n10830, n10447, n10446, 
        n10756, n10445, n3488, n3489, n3490, n3491, n3492, n3493, 
        n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
        n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, 
        n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
        n3518, n3519, n13837, n10757, n10821, n12390, n12389, 
        n12388, n12387, n12386, n12385, n12384, n12383, n12382, 
        n12381, n12380, n12379, n12378, n12377, n12376, n12375, 
        n12374, n10758, n10804, n10759, n10820, n10760, n10805, 
        n10444, n10443, n10442, n10441, n10440, n10439, n10438, 
        n10437, n10436, n10435, n10434, n10433, n10432, n10431, 
        n10430, n10429, n10428, n10427, n10426, n10425, n10424, 
        n10423, n10422, n10421, n10420, n10419, n10761, n10825, 
        n10762, n10799, n10803, n10763, n10822, n10418, n10802, 
        n10844, n10831, n10417, n104_adj_243, n10845, n102_adj_244, 
        n10416, n10829, n10846, n10796, n10415, n10828, n10847, 
        n10797, n10414, n10827, n10848, n10798, n10413, n10826, 
        n10849, n10823, n10412, n10411, n10410, n10409, n10408, 
        n10407, n10406, n10405, n10404, n10403, n10402, n10401, 
        n10400, n10399, n10398, n10397, n10396, n10395, n10850, 
        n10394, n10816, n10851, n10809, n10393, n10815, n10852, 
        n10810, n10392, n10814, n10853, n10811, n10235, n10813, 
        n10854, n68_adj_245, n10234, n10812, n10855, n10795, n10233, 
        n10794, n10856, n10793, n10232, n10792, n10857, n10791, 
        n10231, n10790, n10858, n10789, n10859, n10788, n10860, 
        n10787, n10861, n10786, n10862, n10785, n10863, n10784, 
        n10864, n10783, n10865, n10782, n10866, n10781, n10867, 
        n10780, n10868, n10779, n10869, n10778, n10870, n10777, 
        n10871, n10776, n10872, n10775, n10873, n10774, n10874, 
        n10773, n10875, n10772, n10876, n10771, n10877, n10770, 
        n10878, n10769, n10879, n10768, n10880, n10767, n10881, 
        n10766, n10882, n10765, n10883, n10764, n10884, n10885, 
        n10886, n10887, n10888, n10889, n10890, n10891, n10230, 
        n10892, n10229, n10893, n10228, n10894, n10227, n10895, 
        n10226, n10896, n10225, n10897, n10224, n10898, n10223, 
        n10899, n10222, n10900, n10221, n10901, n10220, n10902, 
        n10219, n10218, n11367, n10217, n11366, n10216, n11365, 
        n10215, n11364, n10214, n11363, n10213, n11362, n10212, 
        n11361, n10211, n11360, n10210, n11359, n10209, n11358, 
        n10208, n11357, n10207, n11356, n10206, n11355, n11354, 
        n11353, n11352, n11351, n11350, n11349, n11348, n11347, 
        n11346, n11345, n11344, n11343, n11342, n11341, n11340, 
        n11339, n11338, n11337, n11336, n11335, n11334, n11333, 
        n11332, n11331, n11330, n11329, n11328, n11327, n11326, 
        n11325, n11324, n11323, n11322, n11321, n11320, n11319, 
        n11318, n11317, n11316, n11315, n11314, n11313, n11312, 
        n11311, n11310, n11309, n11308, n11372, n11373, n11374, 
        n11375, n11376, n11377, n11378, n11379, n11380, n11381, 
        n11382, n11383, n11384, n11385, n11386, n11387, n11388, 
        n11389, n11390, n11391, n11392, n11393, n11394, n11395, 
        n11396, n11397, n11398, n11399, n11400, n11401, n11402, 
        n11403, n11404, n11405, n11406, n11407, n11408, n11409, 
        n11410, n11411, n11412, n11413, n11414, n11415, n11416, 
        n11417, n11418, n11419, n11420, n11421, n11422, n11423, 
        n11424, n11425, n11426, n11427, n11428, n11429, n11430, 
        n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
        n11438, n11439, n11440, n11441, n11442, n11443, n11444, 
        n11445, n11446, n11447, n11448, n11449, n11450, n11451, 
        n11452, n11453, n11454, n11455, n11456, n11457, n11458, 
        n11459, n11460, n11461, n11462, n11463, n11464, n11465, 
        n11466, n11467, n11468, n11469, n11470, n11471, n11472, 
        n11473, n11474, n11475, n11476, n11477, n11478, n11479, 
        n11480, n11481, n11482, n11483, n11484, n11485, n11486, 
        n11487, n11488, n11489, n11490, n11491, n11492, n11493, 
        n11494, n11495, n11496, n11497, n11498, n11499, n11500, 
        n11501, n11502, n11503, n11504, n11505, n11506, n11507, 
        n11508, n11509, n11510, n11511, n11512, n11513, n11514, 
        n11515, n11516, n11517, n11518, n11519, n11520, n11521, 
        n11522, n11523, n11524, n11525, n11526, n11527, n11528, 
        n11529, n11530, n11531, n11532, n11533, n11534, n11535, 
        n11536, n11537, n11538, n11539, n11540, n11541, n11542, 
        n11543, n11544, n11545, n11546, n11547, n11548, n11549, 
        n11550, n11551, n11552, n11553, n11554, n11555, n11556, 
        n11557, n11558, n11559, n11560, n11561, n11562, n11563, 
        n11564, n11565, n11566, n11567, n11568, n11569, n11570, 
        n11571, n11572, n11573, n11574, n11575, n11576, n11577, 
        n11578, n11579, n11580, n11581, n11582, n11583, n11584, 
        n11585, n11586, n11587, n11588, n11589, n11590, n11591, 
        n11592, n11593, n11594, n11595, n11596, n11597, n11598, 
        n11599, n11600, n11601, n11602, n11603, n11604, n11605, 
        n11606, n11607, n11608, n11609, n11610, n11611, n11612, 
        n11613, n11614, n11615, n11616, n11617, n11618, n11619, 
        n11620, n11621, n11622, n11623, n11624, n11625, n11626, 
        n11627, n11628, n11629, n71, n74, n77, n80, n83, n86, 
        n89, n92, n95, n98, n101, n104_adj_246, n107, n110_adj_247, 
        n113, n116_adj_248, n119, n122_adj_249, n125, n128_adj_250, 
        n131, n134, n137, n140, n143, n146, n149, n152, n155, 
        n158, n161, n68_adj_251, n71_adj_252, n74_adj_253, n77_adj_254, 
        n80_adj_255, n83_adj_256, n86_adj_257, n89_adj_258, n92_adj_259, 
        n95_adj_260, n98_adj_261, n101_adj_262, n104_adj_263, n107_adj_264, 
        n110_adj_265, n113_adj_266, n116_adj_267, n119_adj_268, n122_adj_269, 
        n125_adj_270, n128_adj_271, n131_adj_272, n134_adj_273, n137_adj_274, 
        n140_adj_275, n143_adj_276, n146_adj_277, n149_adj_278, n152_adj_279, 
        n155_adj_280, n158_adj_281, n161_adj_282, n68_adj_283, n71_adj_284, 
        n74_adj_285, n77_adj_286, n80_adj_287, n83_adj_288, n86_adj_289, 
        n89_adj_290, n92_adj_291, n95_adj_292, n98_adj_293, n101_adj_294, 
        n104_adj_295, n107_adj_296, n110_adj_297, n113_adj_298, n116_adj_299, 
        n119_adj_300, n122_adj_301, n125_adj_302, n128_adj_303, n131_adj_304, 
        n134_adj_305, n137_adj_306, n140_adj_307, n143_adj_308, n146_adj_309, 
        n149_adj_310, n152_adj_311, n155_adj_312, n158_adj_313, n161_adj_314, 
        n68_adj_315, n71_adj_316, n74_adj_317, n77_adj_318, n80_adj_319, 
        n83_adj_320, n86_adj_321, n89_adj_322, n92_adj_323, n95_adj_324, 
        n98_adj_325, n101_adj_326, n104_adj_327, n107_adj_328, n110_adj_329, 
        n113_adj_330, n116_adj_331, n119_adj_332, n122_adj_333, n125_adj_334, 
        n128_adj_335, n131_adj_336, n134_adj_337, n137_adj_338, n140_adj_339, 
        n143_adj_340, n146_adj_341, n149_adj_342, n152_adj_343, n155_adj_344, 
        n158_adj_345, n161_adj_346, n68_adj_347, n71_adj_348, n74_adj_349, 
        n77_adj_350, n80_adj_351, n83_adj_352, n86_adj_353, n89_adj_354, 
        n92_adj_355, n95_adj_356, n98_adj_357, n101_adj_358, n104_adj_359, 
        n107_adj_360, n110_adj_361, n113_adj_362, n116_adj_363, n119_adj_364, 
        n122_adj_365, n125_adj_366, n128_adj_367, n131_adj_368, n134_adj_369, 
        n137_adj_370, n140_adj_371, n143_adj_372, n146_adj_373, n149_adj_374, 
        n152_adj_375, n155_adj_376, n158_adj_377, n161_adj_378, n68_adj_379, 
        n71_adj_380, n74_adj_381, n77_adj_382, n80_adj_383, n83_adj_384, 
        n86_adj_385, n89_adj_386, n92_adj_387, n95_adj_388, n98_adj_389, 
        n101_adj_390, n104_adj_391, n107_adj_392, n110_adj_393, n113_adj_394, 
        n116_adj_395, n119_adj_396, n122_adj_397, n125_adj_398, n128_adj_399, 
        n131_adj_400, n134_adj_401, n137_adj_402, n140_adj_403, n143_adj_404, 
        n146_adj_405, n149_adj_406, n152_adj_407, n155_adj_408, n158_adj_409, 
        n161_adj_410, n71_adj_411, n74_adj_412, n77_adj_413, n80_adj_414, 
        n83_adj_415, n86_adj_416, n89_adj_417, n92_adj_418, n95_adj_419, 
        n98_adj_420, n101_adj_421, n104_adj_422, n107_adj_423, n110_adj_424, 
        n113_adj_425, n116_adj_426, n119_adj_427, n122_adj_428, n125_adj_429, 
        n128_adj_430, n131_adj_431, n134_adj_432, n137_adj_433, n140_adj_434, 
        n143_adj_435, n146_adj_436, n149_adj_437, n152_adj_438, n155_adj_439, 
        n158_adj_440, n161_adj_441, n68_adj_442, n71_adj_443, n74_adj_444, 
        n77_adj_445, n80_adj_446, n83_adj_447, n86_adj_448, n89_adj_449, 
        n92_adj_450, n95_adj_451, n98_adj_452, n101_adj_453, n104_adj_454, 
        n107_adj_455, n110_adj_456, n113_adj_457, n116_adj_458, n119_adj_459, 
        n122_adj_460, n125_adj_461, n128_adj_462, n131_adj_463, n134_adj_464, 
        n137_adj_465, n140_adj_466, n143_adj_467, n146_adj_468, n149_adj_469, 
        n152_adj_470, n155_adj_471, n158_adj_472, n161_adj_473, n68_adj_474, 
        n71_adj_475, n74_adj_476, n77_adj_477, n80_adj_478, n83_adj_479, 
        n86_adj_480, n89_adj_481, n92_adj_482, n95_adj_483, n98_adj_484, 
        n101_adj_485, n104_adj_486, n107_adj_487, n110_adj_488, n113_adj_489, 
        n116_adj_490, n119_adj_491, n122_adj_492, n125_adj_493, n128_adj_494, 
        n131_adj_495, n134_adj_496, n137_adj_497, n140_adj_498, n143_adj_499, 
        n146_adj_500, n149_adj_501, n152_adj_502, n155_adj_503, n158_adj_504, 
        n161_adj_505, n68_adj_506, n71_adj_507, n74_adj_508, n77_adj_509, 
        n80_adj_510, n83_adj_511, n86_adj_512, n89_adj_513, n92_adj_514, 
        n95_adj_515, n98_adj_516, n101_adj_517, n104_adj_518, n107_adj_519, 
        n110_adj_520, n113_adj_521, n116_adj_522, n119_adj_523, n122_adj_524, 
        n125_adj_525, n128_adj_526, n131_adj_527, n134_adj_528, n137_adj_529, 
        n140_adj_530, n143_adj_531, n146_adj_532, n149_adj_533, n152_adj_534, 
        n155_adj_535, n158_adj_536, n161_adj_537, n68_adj_538, n71_adj_539, 
        n74_adj_540, n77_adj_541, n80_adj_542, n83_adj_543, n86_adj_544, 
        n89_adj_545, n92_adj_546, n95_adj_547, n98_adj_548, n101_adj_549, 
        n104_adj_550, n107_adj_551, n110_adj_552, n113_adj_553, n116_adj_554, 
        n119_adj_555, n122_adj_556, n125_adj_557, n128_adj_558, n131_adj_559, 
        n134_adj_560, n137_adj_561, n140_adj_562, n143_adj_563, n146_adj_564, 
        n149_adj_565, n152_adj_566, n155_adj_567, n158_adj_568, n161_adj_569, 
        n68_adj_570, n71_adj_571, n74_adj_572, n77_adj_573, n80_adj_574, 
        n83_adj_575, n86_adj_576, n89_adj_577, n92_adj_578, n95_adj_579, 
        n98_adj_580, n101_adj_581, n104_adj_582, n107_adj_583, n110_adj_584, 
        n113_adj_585, n116_adj_586, n119_adj_587, n122_adj_588, n125_adj_589, 
        n128_adj_590, n131_adj_591, n134_adj_592, n137_adj_593, n140_adj_594, 
        n143_adj_595, n146_adj_596, n149_adj_597, n152_adj_598, n155_adj_599, 
        n158_adj_600, n161_adj_601, n68_adj_602, n71_adj_603, n74_adj_604, 
        n77_adj_605, n80_adj_606, n83_adj_607, n86_adj_608, n89_adj_609, 
        n92_adj_610, n95_adj_611, n98_adj_612, n101_adj_613, n104_adj_614, 
        n107_adj_615, n110_adj_616, n113_adj_617, n116_adj_618, n119_adj_619, 
        n122_adj_620, n125_adj_621, n128_adj_622, n131_adj_623, n134_adj_624, 
        n137_adj_625, n140_adj_626, n143_adj_627, n146_adj_628, n149_adj_629, 
        n152_adj_630, n155_adj_631, n158_adj_632, n161_adj_633, n68_adj_634, 
        n71_adj_635, n74_adj_636, n77_adj_637, n80_adj_638, n83_adj_639, 
        n86_adj_640, n89_adj_641, n92_adj_642, n95_adj_643, n98_adj_644, 
        n101_adj_645, n104_adj_646, n107_adj_647, n110_adj_648, n113_adj_649, 
        n116_adj_650, n119_adj_651, n122_adj_652, n125_adj_653, n128_adj_654, 
        n131_adj_655, n134_adj_656, n137_adj_657, n140_adj_658, n143_adj_659, 
        n146_adj_660, n149_adj_661, n152_adj_662, n155_adj_663, n158_adj_664, 
        n161_adj_665, n68_adj_666, n71_adj_667, n74_adj_668, n77_adj_669, 
        n80_adj_670, n83_adj_671, n86_adj_672, n89_adj_673, n92_adj_674, 
        n95_adj_675, n98_adj_676, n101_adj_677, n104_adj_678, n107_adj_679, 
        n110_adj_680, n113_adj_681, n116_adj_682, n119_adj_683, n122_adj_684, 
        n125_adj_685, n128_adj_686, n131_adj_687, n134_adj_688, n137_adj_689, 
        n140_adj_690, n143_adj_691, n146_adj_692, n149_adj_693, n152_adj_694, 
        n155_adj_695, n158_adj_696, n161_adj_697, n68_adj_698, n71_adj_699, 
        n74_adj_700, n77_adj_701, n80_adj_702, n83_adj_703, n86_adj_704, 
        n89_adj_705, n92_adj_706, n95_adj_707, n98_adj_708, n101_adj_709, 
        n104_adj_710, n107_adj_711, n110_adj_712, n113_adj_713, n116_adj_714, 
        n119_adj_715, n122_adj_716, n125_adj_717, n128_adj_718, n131_adj_719, 
        n134_adj_720, n137_adj_721, n140_adj_722, n143_adj_723, n146_adj_724, 
        n149_adj_725, n152_adj_726, n155_adj_727, n158_adj_728, n161_adj_729, 
        n68_adj_730, n71_adj_731, n74_adj_732, n77_adj_733, n80_adj_734, 
        n83_adj_735, n86_adj_736, n89_adj_737, n92_adj_738, n95_adj_739, 
        n98_adj_740, n101_adj_741, n104_adj_742, n107_adj_743, n110_adj_744, 
        n113_adj_745, n116_adj_746, n119_adj_747, n122_adj_748, n125_adj_749, 
        n128_adj_750, n131_adj_751, n134_adj_752, n137_adj_753, n140_adj_754, 
        n143_adj_755, n146_adj_756, n149_adj_757, n152_adj_758, n155_adj_759, 
        n158_adj_760, n161_adj_761, n68_adj_762, n71_adj_763, n74_adj_764, 
        n77_adj_765, n80_adj_766, n83_adj_767, n86_adj_768, n89_adj_769, 
        n92_adj_770, n95_adj_771, n98_adj_772, n101_adj_773, n104_adj_774, 
        n107_adj_775, n110_adj_776, n113_adj_777, n116_adj_778, n119_adj_779, 
        n122_adj_780, n125_adj_781, n128_adj_782, n131_adj_783, n134_adj_784, 
        n137_adj_785, n140_adj_786, n143_adj_787, n146_adj_788, n149_adj_789, 
        n152_adj_790, n155_adj_791, n158_adj_792, n161_adj_793, n68_adj_794, 
        n71_adj_795, n74_adj_796, n77_adj_797, n80_adj_798, n83_adj_799, 
        n86_adj_800, n89_adj_801, n92_adj_802, n95_adj_803, n98_adj_804, 
        n101_adj_805, n104_adj_806, n107_adj_807, n110_adj_808, n113_adj_809, 
        n116_adj_810, n119_adj_811, n122_adj_812, n125_adj_813, n128_adj_814, 
        n131_adj_815, n134_adj_816, n137_adj_817, n140_adj_818, n143_adj_819, 
        n146_adj_820, n149_adj_821, n152_adj_822, n155_adj_823, n158_adj_824, 
        n161_adj_825, n68_adj_826, n71_adj_827, n74_adj_828, n77_adj_829, 
        n80_adj_830, n83_adj_831, n86_adj_832, n89_adj_833, n92_adj_834, 
        n95_adj_835, n98_adj_836, n101_adj_837, n104_adj_838, n107_adj_839, 
        n110_adj_840, n113_adj_841, n116_adj_842, n119_adj_843, n122_adj_844, 
        n125_adj_845, n128_adj_846, n131_adj_847, n134_adj_848, n137_adj_849, 
        n140_adj_850, n143_adj_851, n146_adj_852, n149_adj_853, n152_adj_854, 
        n155_adj_855, n158_adj_856, n161_adj_857, n68_adj_858, n71_adj_859, 
        n74_adj_860, n77_adj_861, n80_adj_862, n83_adj_863, n86_adj_864, 
        n89_adj_865, n92_adj_866, n95_adj_867, n98_adj_868, n101_adj_869, 
        n104_adj_870, n107_adj_871, n110_adj_872, n113_adj_873, n116_adj_874, 
        n119_adj_875, n122_adj_876, n125_adj_877, n128_adj_878, n131_adj_879, 
        n134_adj_880, n137_adj_881, n140_adj_882, n143_adj_883, n146_adj_884, 
        n149_adj_885, n152_adj_886, n155_adj_887, n158_adj_888, n161_adj_889, 
        n68_adj_890, n71_adj_891, n74_adj_892, n77_adj_893, n80_adj_894, 
        n83_adj_895, n86_adj_896, n89_adj_897, n92_adj_898, n95_adj_899, 
        n98_adj_900, n101_adj_901, n104_adj_902, n107_adj_903, n110_adj_904, 
        n113_adj_905, n116_adj_906, n119_adj_907, n122_adj_908, n125_adj_909, 
        n128_adj_910, n131_adj_911, n134_adj_912, n137_adj_913, n140_adj_914, 
        n143_adj_915, n146_adj_916, n149_adj_917, n152_adj_918, n155_adj_919, 
        n158_adj_920, n161_adj_921, n68_adj_922, n71_adj_923, n74_adj_924, 
        n77_adj_925, n80_adj_926, n83_adj_927, n86_adj_928, n89_adj_929, 
        n92_adj_930, n95_adj_931, n98_adj_932, n101_adj_933, n104_adj_934, 
        n107_adj_935, n110_adj_936, n113_adj_937, n116_adj_938, n119_adj_939, 
        n122_adj_940, n125_adj_941, n128_adj_942, n131_adj_943, n134_adj_944, 
        n137_adj_945, n140_adj_946, n143_adj_947, n146_adj_948, n149_adj_949, 
        n152_adj_950, n155_adj_951, n158_adj_952, n161_adj_953, n68_adj_954, 
        n71_adj_955, n74_adj_956, n77_adj_957, n80_adj_958, n83_adj_959, 
        n86_adj_960, n89_adj_961, n92_adj_962, n95_adj_963, n98_adj_964, 
        n101_adj_965, n104_adj_966, n107_adj_967, n110_adj_968, n113_adj_969, 
        n116_adj_970, n119_adj_971, n122_adj_972, n125_adj_973, n128_adj_974, 
        n131_adj_975, n134_adj_976, n137_adj_977, n140_adj_978, n143_adj_979, 
        n146_adj_980, n149_adj_981, n152_adj_982, n155_adj_983, n158_adj_984, 
        n161_adj_985, n68_adj_986, n71_adj_987, n74_adj_988, n77_adj_989, 
        n80_adj_990, n83_adj_991, n86_adj_992, n89_adj_993, n92_adj_994, 
        n95_adj_995, n98_adj_996, n101_adj_997, n104_adj_998, n107_adj_999, 
        n110_adj_1000, n113_adj_1001, n116_adj_1002, n119_adj_1003, 
        n122_adj_1004, n125_adj_1005, n128_adj_1006, n131_adj_1007, 
        n134_adj_1008, n137_adj_1009, n140_adj_1010, n143_adj_1011, 
        n146_adj_1012, n149_adj_1013, n152_adj_1014, n155_adj_1015, 
        n158_adj_1016, n161_adj_1017, n68_adj_1018, n71_adj_1019, n74_adj_1020, 
        n77_adj_1021, n80_adj_1022, n83_adj_1023, n86_adj_1024, n89_adj_1025, 
        n92_adj_1026, n95_adj_1027, n98_adj_1028, n101_adj_1029, n104_adj_1030, 
        n107_adj_1031, n110_adj_1032, n113_adj_1033, n116_adj_1034, 
        n119_adj_1035, n122_adj_1036, n125_adj_1037, n128_adj_1038, 
        n131_adj_1039, n134_adj_1040, n137_adj_1041, n140_adj_1042, 
        n143_adj_1043, n146_adj_1044, n149_adj_1045, n152_adj_1046, 
        n155_adj_1047, n158_adj_1048, n161_adj_1049, n68_adj_1050, n71_adj_1051, 
        n74_adj_1052, n77_adj_1053, n80_adj_1054, n83_adj_1055, n86_adj_1056, 
        n89_adj_1057, n92_adj_1058, n95_adj_1059, n98_adj_1060, n101_adj_1061, 
        n104_adj_1062, n107_adj_1063, n110_adj_1064, n113_adj_1065, 
        n116_adj_1066, n119_adj_1067, n122_adj_1068, n125_adj_1069, 
        n128_adj_1070, n131_adj_1071, n134_adj_1072, n137_adj_1073, 
        n140_adj_1074, n143_adj_1075, n146_adj_1076, n149_adj_1077, 
        n152_adj_1078, n155_adj_1079, n158_adj_1080, n161_adj_1081, 
        n68_adj_1082, n71_adj_1083, n74_adj_1084, n77_adj_1085, n80_adj_1086, 
        n83_adj_1087, n86_adj_1088, n89_adj_1089, n92_adj_1090, n95_adj_1091, 
        n98_adj_1092, n101_adj_1093, n104_adj_1094, n107_adj_1095, n110_adj_1096, 
        n113_adj_1097, n116_adj_1098, n119_adj_1099, n122_adj_1100, 
        n125_adj_1101, n128_adj_1102, n131_adj_1103, n134_adj_1104, 
        n137_adj_1105, n140_adj_1106, n143_adj_1107, n146_adj_1108, 
        n149_adj_1109, n152_adj_1110, n155_adj_1111, n158_adj_1112, 
        n161_adj_1113, n68_adj_1114, n71_adj_1115, n74_adj_1116, n77_adj_1117, 
        n80_adj_1118, n83_adj_1119, n86_adj_1120, n89_adj_1121, n92_adj_1122, 
        n95_adj_1123, n98_adj_1124, n101_adj_1125, n104_adj_1126, n107_adj_1127, 
        n110_adj_1128, n113_adj_1129, n116_adj_1130, n119_adj_1131, 
        n122_adj_1132, n125_adj_1133, n128_adj_1134, n131_adj_1135, 
        n134_adj_1136, n137_adj_1137, n140_adj_1138, n143_adj_1139, 
        n146_adj_1140, n149_adj_1141, n152_adj_1142, n155_adj_1143, 
        n158_adj_1144, n161_adj_1145, n68_adj_1146, n71_adj_1147, n74_adj_1148, 
        n77_adj_1149, n80_adj_1150, n83_adj_1151, n86_adj_1152, n89_adj_1153, 
        n92_adj_1154, n95_adj_1155, n98_adj_1156, n101_adj_1157, n104_adj_1158, 
        n107_adj_1159, n110_adj_1160, n113_adj_1161, n116_adj_1162, 
        n119_adj_1163, n122_adj_1164, n125_adj_1165, n128_adj_1166, 
        n131_adj_1167, n134_adj_1168, n137_adj_1169, n140_adj_1170, 
        n143_adj_1171, n146_adj_1172, n149_adj_1173, n152_adj_1174, 
        n155_adj_1175, n158_adj_1176, n161_adj_1177, n71_adj_1178, n74_adj_1179, 
        n77_adj_1180, n80_adj_1181, n83_adj_1182, n86_adj_1183, n89_adj_1184, 
        n92_adj_1185, n95_adj_1186, n98_adj_1187, n101_adj_1188, n104_adj_1189, 
        n107_adj_1190, n110_adj_1191, n113_adj_1192, n116_adj_1193, 
        n119_adj_1194, n122_adj_1195, n125_adj_1196, n128_adj_1197, 
        n131_adj_1198, n134_adj_1199, n137_adj_1200, n140_adj_1201, 
        n143_adj_1202, n146_adj_1203, n149_adj_1204, n152_adj_1205, 
        n155_adj_1206, n158_adj_1207, n161_adj_1208, n68_adj_1209, n71_adj_1210, 
        n74_adj_1211, n77_adj_1212, n80_adj_1213, n83_adj_1214, n86_adj_1215, 
        n89_adj_1216, n92_adj_1217, n95_adj_1218, n98_adj_1219, n101_adj_1220, 
        n104_adj_1221, n107_adj_1222, n110_adj_1223, n113_adj_1224, 
        n116_adj_1225, n119_adj_1226, n122_adj_1227, n125_adj_1228, 
        n128_adj_1229, n131_adj_1230, n134_adj_1231, n137_adj_1232, 
        n140_adj_1233, n143_adj_1234, n146_adj_1235, n149_adj_1236, 
        n152_adj_1237, n155_adj_1238, n158_adj_1239, n161_adj_1240, 
        n68_adj_1241, n71_adj_1242, n74_adj_1243, n77_adj_1244, n80_adj_1245, 
        n83_adj_1246, n86_adj_1247, n89_adj_1248, n92_adj_1249, n95_adj_1250, 
        n98_adj_1251, n101_adj_1252, n104_adj_1253, n107_adj_1254, n110_adj_1255, 
        n113_adj_1256, n116_adj_1257, n119_adj_1258, n122_adj_1259, 
        n125_adj_1260, n128_adj_1261, n131_adj_1262, n134_adj_1263, 
        n137_adj_1264, n140_adj_1265, n143_adj_1266, n146_adj_1267, 
        n149_adj_1268, n152_adj_1269, n155_adj_1270, n158_adj_1271, 
        n161_adj_1272, n71_adj_1273, n74_adj_1274, n77_adj_1275, n80_adj_1276, 
        n83_adj_1277, n86_adj_1278, n89_adj_1279, n92_adj_1280, n95_adj_1281, 
        n98_adj_1282, n101_adj_1283, n104_adj_1284, n107_adj_1285, n110_adj_1286, 
        n113_adj_1287, n116_adj_1288, n119_adj_1289, n122_adj_1290, 
        n125_adj_1291, n128_adj_1292, n131_adj_1293, n134_adj_1294, 
        n137_adj_1295, n140_adj_1296, n143_adj_1297, n146_adj_1298, 
        n149_adj_1299, n152_adj_1300, n155_adj_1301, n158_adj_1302, 
        n161_adj_1303, n68_adj_1304, n71_adj_1305, n74_adj_1306, n77_adj_1307, 
        n80_adj_1308, n83_adj_1309, n86_adj_1310, n89_adj_1311, n92_adj_1312, 
        n95_adj_1313, n98_adj_1314, n101_adj_1315, n104_adj_1316, n107_adj_1317, 
        n110_adj_1318, n113_adj_1319, n116_adj_1320, n119_adj_1321, 
        n122_adj_1322, n125_adj_1323, n128_adj_1324, n131_adj_1325, 
        n134_adj_1326, n137_adj_1327, n140_adj_1328, n143_adj_1329, 
        n146_adj_1330, n149_adj_1331, n152_adj_1332, n155_adj_1333, 
        n158_adj_1334, n68_adj_1335, n71_adj_1336, n74_adj_1337, n77_adj_1338, 
        n80_adj_1339, n83_adj_1340, n86_adj_1341, n89_adj_1342, n92_adj_1343, 
        n95_adj_1344, n98_adj_1345, n101_adj_1346, n104_adj_1347, n107_adj_1348, 
        n110_adj_1349, n113_adj_1350, n116_adj_1351, n119_adj_1352, 
        n122_adj_1353, n125_adj_1354, n128_adj_1355, n131_adj_1356, 
        n134_adj_1357, n137_adj_1358, n140_adj_1359, n143_adj_1360, 
        n146_adj_1361, n149_adj_1362, n152_adj_1363, n155_adj_1364, 
        n158_adj_1365, n161_adj_1366, n68_adj_1367, n71_adj_1368, n74_adj_1369, 
        n77_adj_1370, n80_adj_1371, n83_adj_1372, n86_adj_1373, n89_adj_1374, 
        n92_adj_1375, n95_adj_1376, n98_adj_1377, n101_adj_1378, n104_adj_1379, 
        n107_adj_1380, n110_adj_1381, n113_adj_1382, n116_adj_1383, 
        n119_adj_1384, n122_adj_1385, n125_adj_1386, n128_adj_1387, 
        n131_adj_1388, n134_adj_1389, n137_adj_1390, n140_adj_1391, 
        n143_adj_1392, n146_adj_1393, n149_adj_1394, n152_adj_1395, 
        n155_adj_1396, n158_adj_1397, n68_adj_1398, n71_adj_1399, n74_adj_1400, 
        n77_adj_1401, n80_adj_1402, n83_adj_1403, n86_adj_1404, n89_adj_1405, 
        n92_adj_1406, n95_adj_1407, n98_adj_1408, n101_adj_1409, n104_adj_1410, 
        n107_adj_1411, n110_adj_1412, n113_adj_1413, n116_adj_1414, 
        n119_adj_1415, n122_adj_1416, n125_adj_1417, n128_adj_1418, 
        n131_adj_1419, n134_adj_1420, n137_adj_1421, n140_adj_1422, 
        n143_adj_1423, n146_adj_1424, n149_adj_1425, n152_adj_1426, 
        n155_adj_1427, n158_adj_1428, n161_adj_1429, n68_adj_1430, n71_adj_1431, 
        n74_adj_1432, n77_adj_1433, n80_adj_1434, n83_adj_1435, n86_adj_1436, 
        n89_adj_1437, n92_adj_1438, n95_adj_1439, n98_adj_1440, n101_adj_1441, 
        n104_adj_1442, n107_adj_1443, n110_adj_1444, n113_adj_1445, 
        n116_adj_1446, n119_adj_1447, n122_adj_1448, n125_adj_1449, 
        n128_adj_1450, n131_adj_1451, n134_adj_1452, n137_adj_1453, 
        n140_adj_1454, n143_adj_1455, n146_adj_1456, n149_adj_1457, 
        n152_adj_1458, n155_adj_1459, n158_adj_1460, n161_adj_1461, 
        n68_adj_1462, n71_adj_1463, n74_adj_1464, n77_adj_1465, n80_adj_1466, 
        n83_adj_1467, n86_adj_1468, n89_adj_1469, n92_adj_1470, n95_adj_1471, 
        n98_adj_1472, n101_adj_1473, n104_adj_1474, n107_adj_1475, n110_adj_1476, 
        n113_adj_1477, n116_adj_1478, n119_adj_1479, n122_adj_1480, 
        n125_adj_1481, n128_adj_1482, n131_adj_1483, n134_adj_1484, 
        n137_adj_1485, n140_adj_1486, n143_adj_1487, n146_adj_1488, 
        n149_adj_1489, n152_adj_1490, n155_adj_1491, n158_adj_1492, 
        n161_adj_1493, n68_adj_1494, n71_adj_1495, n74_adj_1496, n77_adj_1497, 
        n80_adj_1498, n83_adj_1499, n86_adj_1500, n89_adj_1501, n92_adj_1502, 
        n95_adj_1503, n98_adj_1504, n101_adj_1505, n104_adj_1506, n107_adj_1507, 
        n110_adj_1508, n113_adj_1509, n116_adj_1510, n119_adj_1511, 
        n122_adj_1512, n125_adj_1513, n128_adj_1514, n131_adj_1515, 
        n134_adj_1516, n137_adj_1517, n140_adj_1518, n143_adj_1519, 
        n146_adj_1520, n149_adj_1521, n152_adj_1522, n155_adj_1523, 
        n158_adj_1524, n71_adj_1525, n74_adj_1526, n77_adj_1527, n80_adj_1528, 
        n83_adj_1529, n86_adj_1530, n89_adj_1531, n92_adj_1532, n95_adj_1533, 
        n98_adj_1534, n101_adj_1535, n104_adj_1536, n107_adj_1537, n110_adj_1538, 
        n113_adj_1539, n116_adj_1540, n119_adj_1541, n122_adj_1542, 
        n125_adj_1543, n128_adj_1544, n131_adj_1545, n134_adj_1546, 
        n137_adj_1547, n140_adj_1548, n143_adj_1549, n146_adj_1550, 
        n149_adj_1551, n152_adj_1552, n155_adj_1553, n158_adj_1554, 
        n161_adj_1555, n68_adj_1556, n71_adj_1557, n74_adj_1558, n77_adj_1559, 
        n80_adj_1560, n83_adj_1561, n86_adj_1562, n89_adj_1563, n92_adj_1564, 
        n95_adj_1565, n98_adj_1566, n101_adj_1567, n104_adj_1568, n107_adj_1569, 
        n110_adj_1570, n113_adj_1571, n116_adj_1572, n119_adj_1573, 
        n122_adj_1574, n125_adj_1575, n128_adj_1576, n131_adj_1577, 
        n134_adj_1578, n137_adj_1579, n140_adj_1580, n143_adj_1581, 
        n146_adj_1582, n149_adj_1583, n152_adj_1584, n155_adj_1585, 
        n158_adj_1586, n161_adj_1587, n68_adj_1588, n71_adj_1589, n74_adj_1590, 
        n77_adj_1591, n80_adj_1592, n83_adj_1593, n86_adj_1594, n89_adj_1595, 
        n92_adj_1596, n95_adj_1597, n98_adj_1598, n101_adj_1599, n104_adj_1600, 
        n107_adj_1601, n110_adj_1602, n113_adj_1603, n116_adj_1604, 
        n119_adj_1605, n122_adj_1606, n125_adj_1607, n128_adj_1608, 
        n131_adj_1609, n134_adj_1610, n137_adj_1611, n140_adj_1612, 
        n143_adj_1613, n146_adj_1614, n149_adj_1615, n152_adj_1616, 
        n155_adj_1617, n158_adj_1618, n161_adj_1619, n68_adj_1620, n71_adj_1621, 
        n74_adj_1622, n77_adj_1623, n80_adj_1624, n83_adj_1625, n86_adj_1626, 
        n89_adj_1627, n92_adj_1628, n95_adj_1629, n98_adj_1630, n101_adj_1631, 
        n104_adj_1632, n107_adj_1633, n110_adj_1634, n113_adj_1635, 
        n116_adj_1636, n119_adj_1637, n122_adj_1638, n125_adj_1639, 
        n128_adj_1640, n131_adj_1641, n134_adj_1642, n137_adj_1643, 
        n140_adj_1644, n143_adj_1645, n146_adj_1646, n149_adj_1647, 
        n152_adj_1648, n155_adj_1649, n158_adj_1650, n161_adj_1651, 
        n68_adj_1652, n68_adj_1653, n71_adj_1654, n74_adj_1655, n77_adj_1656, 
        n80_adj_1657, n83_adj_1658, n86_adj_1659, n89_adj_1660, n92_adj_1661, 
        n95_adj_1662, n98_adj_1663, n101_adj_1664, n104_adj_1665, n107_adj_1666, 
        n110_adj_1667, n113_adj_1668, n116_adj_1669, n119_adj_1670, 
        n122_adj_1671, n125_adj_1672, n128_adj_1673, n131_adj_1674, 
        n134_adj_1675, n137_adj_1676, n140_adj_1677, n143_adj_1678, 
        n146_adj_1679, n149_adj_1680, n152_adj_1681, n155_adj_1682, 
        n158_adj_1683, n161_adj_1684, n68_adj_1685, n71_adj_1686, n74_adj_1687, 
        n77_adj_1688, n80_adj_1689, n83_adj_1690, n86_adj_1691, n89_adj_1692, 
        n92_adj_1693, n95_adj_1694, n98_adj_1695, n101_adj_1696, n104_adj_1697, 
        n107_adj_1698, n110_adj_1699, n113_adj_1700, n116_adj_1701, 
        n119_adj_1702, n122_adj_1703, n125_adj_1704, n128_adj_1705, 
        n131_adj_1706, n134_adj_1707, n137_adj_1708, n140_adj_1709, 
        n143_adj_1710, n146_adj_1711, n149_adj_1712, n152_adj_1713, 
        n155_adj_1714, n158_adj_1715, n161_adj_1716, n13565, n13564, 
        n13563, n13562, n13561, n13560, n13559, n13558, n13557, 
        n13556, n13555, n13554, n13553, n13552, n13551, n13550, 
        n13549, n13548, n13547, n13546, n13545, n13544, n13543, 
        n13542, n13541, n13540, n13539, n13538, n13537, n13536, 
        n13535, n13534, n13533, n13532, n13531, n13530, n13529, 
        n13528, n13527, n13526, n13525, n13524, n13523, n13522, 
        n13521, n13520, n13519, n13518, n13517, n68_adj_1717, n13516, 
        n71_adj_1718, n13515, n74_adj_1719, n13514, n77_adj_1720, 
        n13513, n80_adj_1721, n13512, n83_adj_1722, n13511, n86_adj_1723, 
        n13510, n89_adj_1724, n13509, n92_adj_1725, n13508, n95_adj_1726, 
        n13507, n98_adj_1727, n13506, n101_adj_1728, n13505, n104_adj_1729, 
        n13504, n107_adj_1730, n13503, n110_adj_1731, n13502, n113_adj_1732, 
        n13501, n116_adj_1733, n13500, n119_adj_1734, n13499, n122_adj_1735, 
        n13498, n125_adj_1736, n13497, n128_adj_1737, n13496, n131_adj_1738, 
        n13495, n134_adj_1739, n13494, n137_adj_1740, n13493, n140_adj_1741, 
        n13492, n143_adj_1742, n13491, n146_adj_1743, n13490, n149_adj_1744, 
        n13489, n152_adj_1745, n13488, n155_adj_1746, n13487, n158_adj_1747, 
        n13486, n161_adj_1748, n13485, n13484, n13483, n13482, n13481, 
        n13480, n13479, n13478, n13477, n13476, n13475, n13474, 
        n13473, n13472, n13471, n13469, n13468, n13467, n13466, 
        n13465, n13464, n13463, n13462, n13461, n13460, n13459, 
        n13458, n13457, n13456, n13455, n13454, n13450, n13449, 
        n13448, n13447, n13446, n13445, n13444, n13443, n13442, 
        n13441, n13440, n13439, n13438, n13437, n13436, n13435, 
        n13434, n13433, n13432, n13431, n13430, n13429, n13428, 
        n13427, n13426, n13425, n13424, n13423, n13422, n13421, 
        n13420, n68_adj_1749, n13419, n71_adj_1750, n74_adj_1751, 
        n13417, n77_adj_1752, n13416, n80_adj_1753, n13415, n83_adj_1754, 
        n13414, n86_adj_1755, n13413, n89_adj_1756, n13412, n92_adj_1757, 
        n13411, n95_adj_1758, n13410, n98_adj_1759, n101_adj_1760, 
        n13408, n104_adj_1761, n13407, n107_adj_1762, n13406, n110_adj_1763, 
        n13405, n113_adj_1764, n13404, n116_adj_1765, n13403, n119_adj_1766, 
        n13402, n122_adj_1767, n13401, n125_adj_1768, n13400, n128_adj_1769, 
        n13399, n131_adj_1770, n13398, n134_adj_1771, n13397, n137_adj_1772, 
        n13396, n140_adj_1773, n13395, n143_adj_1774, n13394, n146_adj_1775, 
        n13392, n149_adj_1776, n13391, n152_adj_1777, n13390, n155_adj_1778, 
        n13389, n158_adj_1779, n13388, n13387, n13386, n13385, n13384, 
        n13383, n13382, n13381, n13380, n13379, n13378, n13377, 
        n13376, n13375, n13374, n13373, n13372, n13371, n13370, 
        n13369, n13368, n13367, n13366, n13365, n13364, n13363, 
        n13362, n13361, n13360, n13359, n13358, n13357, n13356, 
        n13355, n13354, n13353, n13352, n13351, n13350, n13349, 
        n13348, n13347, n13346, n13345, n13344, n13343, n13342, 
        n13341, n13340, n13339, n13338, n13337, n13336, n13335, 
        n13334, n13333, n13332, n13331, n13330, n13329, n13328, 
        n13327, n13326, n13325, n13324, n13323, n13322, n68_adj_1780, 
        n13321, n71_adj_1781, n13320, n74_adj_1782, n13319, n77_adj_1783, 
        n13318, n80_adj_1784, n13317, n83_adj_1785, n13316, n86_adj_1786, 
        n13315, n89_adj_1787, n13314, n92_adj_1788, n13313, n95_adj_1789, 
        n98_adj_1790, n13311, n101_adj_1791, n13310, n104_adj_1792, 
        n13309, n107_adj_1793, n13308, n110_adj_1794, n13307, n113_adj_1795, 
        n13306, n116_adj_1796, n13305, n119_adj_1797, n13304, n122_adj_1798, 
        n13303, n125_adj_1799, n13302, n128_adj_1800, n13301, n131_adj_1801, 
        n13300, n134_adj_1802, n13299, n137_adj_1803, n13298, n140_adj_1804, 
        n13297, n143_adj_1805, n13295, n146_adj_1806, n13294, n149_adj_1807, 
        n13293, n152_adj_1808, n13292, n155_adj_1809, n13291, n158_adj_1810, 
        n13290, n161_adj_1811, n13289, n13288, n13287, n13286, n13285, 
        n13284, n13283, n13282, n13281, n13280, n13279, n13278, 
        n13277, n13276, n13275, n13274, n13273, n13272, n13271, 
        n13270, n13269, n13268, n13267, n13266, n13265, n13264, 
        n13263, n13262, n13261, n13260, n13259, n13258, n13257, 
        n13256, n13255, n13254, n13253, n13252, n13251, n13250, 
        n13249, n13248, n13246, n13245, n13244, n13243, n13242, 
        n13241, n13240, n13239, n13238, n13237, n13236, n13235, 
        n13234, n13233, n13232, n13231, n13230, n13229, n13228, 
        n13227, n13226, n13225, n13224, n68_adj_1812, n13223, n71_adj_1813, 
        n13222, n74_adj_1814, n13221, n77_adj_1815, n13220, n80_adj_1816, 
        n13219, n83_adj_1817, n13218, n86_adj_1818, n13217, n89_adj_1819, 
        n13216, n92_adj_1820, n13215, n95_adj_1821, n13214, n98_adj_1822, 
        n13213, n101_adj_1823, n13212, n104_adj_1824, n13211, n107_adj_1825, 
        n13210, n110_adj_1826, n13209, n113_adj_1827, n13208, n116_adj_1828, 
        n13207, n119_adj_1829, n13206, n122_adj_1830, n13205, n125_adj_1831, 
        n13204, n128_adj_1832, n13203, n131_adj_1833, n13202, n134_adj_1834, 
        n13201, n137_adj_1835, n13200, n140_adj_1836, n13199, n143_adj_1837, 
        n13198, n146_adj_1838, n13197, n149_adj_1839, n13196, n152_adj_1840, 
        n13195, n155_adj_1841, n13194, n158_adj_1842, n13193, n161_adj_1843, 
        n13192, n13191, n13190, n13189, n13188, n13187, n13186, 
        n13185, n13184, n13182, n13181, n13180, n13179, n13178, 
        n13177, n13176, n13175, n13174, n13173, n13172, n13171, 
        n13170, n13169, n13168, n13167, n13162, n13161, n13160, 
        n13159, n13158, n13157, n13156, n13155, n13154, n13153, 
        n13152, n13151, n13150, n13149, n13148, n13145, n13144, 
        n13143, n13142, n13141, n13140, n13139, n13138, n13137, 
        n13136, n13135, n13134, n13133, n13132, n13131, n13130, 
        n13129, n13128, n13127, n13126, n13125, n68_adj_1844, n13124, 
        n71_adj_1845, n13123, n74_adj_1846, n13122, n77_adj_1847, 
        n13121, n80_adj_1848, n13120, n83_adj_1849, n13119, n86_adj_1850, 
        n13118, n89_adj_1851, n13117, n92_adj_1852, n13116, n95_adj_1853, 
        n13115, n98_adj_1854, n13114, n101_adj_1855, n13113, n104_adj_1856, 
        n13112, n107_adj_1857, n13111, n110_adj_1858, n13110, n113_adj_1859, 
        n13109, n116_adj_1860, n13108, n119_adj_1861, n13107, n122_adj_1862, 
        n13106, n125_adj_1863, n13105, n128_adj_1864, n13104, n131_adj_1865, 
        n13103, n134_adj_1866, n13102, n137_adj_1867, n13101, n140_adj_1868, 
        n13100, n143_adj_1869, n13099, n146_adj_1870, n13098, n149_adj_1871, 
        n13097, n152_adj_1872, n13096, n155_adj_1873, n13095, n158_adj_1874, 
        n13094, n161_adj_1875, n13093, n13092, n13091, n13090, n13088, 
        n13087, n13086, n13085, n13084, n13083, n13082, n13081, 
        n13080, n13079, n13078, n13077, n13076, n13075, n13074, 
        n13071, n13070, n13069, n13068, n13067, n13066, n13065, 
        n13064, n13063, n13062, n13061, n13060, n13059, n13058, 
        n13057, n13054, n13053, n13052, n13051, n13050, n13049, 
        n13048, n13047, n13046, n13045, n13044, n13043, n13042, 
        n13041, n13040, n13037, n13036, n13035, n13034, n13033, 
        n13032, n13031, n13030, n13029, n13028, n13027, n13026, 
        n13025, n68_adj_1876, n13024, n71_adj_1877, n13023, n74_adj_1878, 
        n13022, n77_adj_1879, n80_adj_1880, n83_adj_1881, n86_adj_1882, 
        n13017, n89_adj_1883, n13016, n92_adj_1884, n13015, n95_adj_1885, 
        n13014, n98_adj_1886, n13013, n101_adj_1887, n13012, n104_adj_1888, 
        n13011, n107_adj_1889, n13010, n110_adj_1890, n13009, n113_adj_1891, 
        n13008, n116_adj_1892, n13007, n119_adj_1893, n13006, n122_adj_1894, 
        n13005, n125_adj_1895, n13004, n128_adj_1896, n13003, n131_adj_1897, 
        n134_adj_1898, n13000, n137_adj_1899, n12999, n140_adj_1900, 
        n12998, n143_adj_1901, n12997, n146_adj_1902, n12996, n149_adj_1903, 
        n12995, n152_adj_1904, n12994, n155_adj_1905, n12993, n158_adj_1906, 
        n12992, n161_adj_1907, n12991, n12990, n12989, n12988, n12987, 
        n12986, n12985, n12980, n12979, n12978, n12977, n12976, 
        n12975, n12974, n12973, n12972, n12971, n12970, n12969, 
        n12968, n12967, n12966, n12964, n12963, n12962, n12961, 
        n12960, n12959, n12958, n12957, n12956, n12955, n12954, 
        n12953, n12952, n12951, n12950, n12948, n12947, n12946, 
        n12945, n12944, n12943, n12942, n12941, n12940, n12939, 
        n12938, n12937, n12936, n12935, n12934, n12932, n12931, 
        n12930, n12929, n12928, n12927, n12926, n12925, n68_adj_1908, 
        n12924, n71_adj_1909, n12923, n74_adj_1910, n12922, n77_adj_1911, 
        n12921, n80_adj_1912, n12920, n83_adj_1913, n12919, n86_adj_1914, 
        n12918, n89_adj_1915, n12917, n92_adj_1916, n12916, n95_adj_1917, 
        n12915, n98_adj_1918, n12914, n101_adj_1919, n12913, n104_adj_1920, 
        n12912, n107_adj_1921, n12911, n110_adj_1922, n12910, n113_adj_1923, 
        n12909, n116_adj_1924, n12908, n119_adj_1925, n12907, n122_adj_1926, 
        n12906, n125_adj_1927, n12905, n128_adj_1928, n12904, n131_adj_1929, 
        n12903, n134_adj_1930, n12902, n137_adj_1931, n140_adj_1932, 
        n12900, n143_adj_1933, n12899, n146_adj_1934, n12898, n149_adj_1935, 
        n12897, n152_adj_1936, n12896, n155_adj_1937, n12895, n158_adj_1938, 
        n12894, n161_adj_1939, n12893, n12892, n12891, n12890, n12889, 
        n12888, n12887, n12886, n12885, n12881, n12880, n12879, 
        n12878, n12877, n12876, n12875, n12874, n12873, n12872, 
        n12871, n12870, n12869, n12868, n12867, n12866, n12865, 
        n12864, n12863, n12862, n12861, n12860, n12859, n12858, 
        n12857, n12856, n12855, n12854, n12853, n12852, n12851, 
        n12850, n12849, n12848, n12847, n12846, n12845, n12844, 
        n12843, n12842, n12841, n12840, n12839, n12838, n12837, 
        n12836, n12835, n12834, n12833, n12832, n12831, n12830, 
        n12829, n12828, n12827, n68_adj_1940, n12826, n71_adj_1941, 
        n12825, n74_adj_1942, n12824, n77_adj_1943, n12823, n80_adj_1944, 
        n12822, n83_adj_1945, n12821, n86_adj_1946, n12820, n89_adj_1947, 
        n12819, n92_adj_1948, n12818, n95_adj_1949, n12817, n98_adj_1950, 
        n12816, n101_adj_1951, n12815, n104_adj_1952, n12814, n107_adj_1953, 
        n12813, n110_adj_1954, n12812, n113_adj_1955, n12811, n116_adj_1956, 
        n12810, n119_adj_1957, n12809, n122_adj_1958, n12808, n125_adj_1959, 
        n12807, n128_adj_1960, n12806, n131_adj_1961, n12805, n134_adj_1962, 
        n12804, n137_adj_1963, n12803, n140_adj_1964, n12802, n143_adj_1965, 
        n12801, n146_adj_1966, n12800, n149_adj_1967, n12799, n152_adj_1968, 
        n12798, n155_adj_1969, n12797, n158_adj_1970, n12796, n12795, 
        n12794, n12793, n12792, n12791, n12790, n12789, n12788, 
        n12787, n12786, n12785, n12784, n12783, n12782, n12781, 
        n12780, n12779, n12778, n12777, n12776, n12775, n12774, 
        n12773, n12772, n12771, n12770, n12769, n12768, n12767, 
        n12766, n12765, n12764, n12763, n12762, n12761, n12760, 
        n12759, n12758, n12757, n12756, n12755, n12754, n12753, 
        n12752, n12751, n12750, n12749, n12748, n12747, n12746, 
        n12745, n12744, n12743, n12742, n12741, n12740, n12739, 
        n12738, n12737, n12736, n12735, n12734, n12733, n12732, 
        n12731, n12730, n12729, n12728, n12727, n12726, n12725, 
        n12724, n12723, n12722, n12721, n12720, n12719, n12718, 
        n12717, n12716, n12715, n12714, n12713, n12712, n12711, 
        n12710, n12709, n12708, n12707, n12706, n12705, n12704, 
        n12703, n12702, n12701, n12700, n12699, n12698, n12697, 
        n12696, n68_adj_1971, n12695, n71_adj_1972, n12694, n74_adj_1973, 
        n12693, n77_adj_1974, n12692, n80_adj_1975, n12691, n83_adj_1976, 
        n12690, n86_adj_1977, n12689, n89_adj_1978, n12688, n92_adj_1979, 
        n12687, n95_adj_1980, n12686, n98_adj_1981, n12685, n101_adj_1982, 
        n12684, n104_adj_1983, n12683, n107_adj_1984, n12682, n110_adj_1985, 
        n12681, n113_adj_1986, n12680, n116_adj_1987, n12679, n119_adj_1988, 
        n12678, n122_adj_1989, n12677, n125_adj_1990, n12676, n128_adj_1991, 
        n12675, n131_adj_1992, n12674, n134_adj_1993, n12673, n137_adj_1994, 
        n12672, n140_adj_1995, n12671, n143_adj_1996, n12670, n146_adj_1997, 
        n12669, n149_adj_1998, n12668, n152_adj_1999, n12667, n155_adj_2000, 
        n12666, n158_adj_2001, n12665, n161_adj_2002, n12664, n12663, 
        n12662, n12661, n12660, n12659, n12658, n12657, n12656, 
        n12655, n12654, n12653, n12652, n12651, n12650, n12649, 
        n12648, n12647, n12646, n12645, n12644, n12643, n12642, 
        n12641, n12640, n12639, n12638, n12637, n12636, n12635, 
        n12634, n12633, n12632, n12631, n12630, n12629, n12628, 
        n12627, n12626, n12625, n12624, n12623, n12622, n12621, 
        n12620, n12619, n12618, n12617, n12616, n12615, n12614, 
        n12613, n12612, n12611, n12610, n12609, n12608, n12607, 
        n12606, n12605, n12604, n12603, n12602, n12601, n12600, 
        n12599, n68_adj_2003, n12598, n71_adj_2004, n12597, n74_adj_2005, 
        n12596, n77_adj_2006, n12595, n80_adj_2007, n12594, n83_adj_2008, 
        n86_adj_2009, n12592, n89_adj_2010, n12591, n92_adj_2011, 
        n12590, n95_adj_2012, n12589, n98_adj_2013, n12588, n101_adj_2014, 
        n12587, n104_adj_2015, n12586, n107_adj_2016, n12585, n110_adj_2017, 
        n12584, n113_adj_2018, n12583, n116_adj_2019, n12582, n119_adj_2020, 
        n12581, n122_adj_2021, n12580, n125_adj_2022, n12579, n128_adj_2023, 
        n12578, n131_adj_2024, n12577, n134_adj_2025, n137_adj_2026, 
        n140_adj_2027, n12573, n143_adj_2028, n12572, n146_adj_2029, 
        n12571, n149_adj_2030, n12570, n152_adj_2031, n12569, n155_adj_2032, 
        n12568, n158_adj_2033, n12567, n161_adj_2034, n12566, n12565, 
        n12564, n12563, n12562, n12561, n12560, n12559, n12558, 
        n12557, n12556, n12555, n12554, n12553, n12552, n12551, 
        n12550, n12549, n12548, n12547, n12546, n12545, n12544, 
        n12543, n12542, n12541, n12540, n12539, n12538, n12537, 
        n12536, n12535, n12534, n12533, n12532, n12531, n12530, 
        n12529, n12528, n12527, n12526, n12524, n12523, n12522, 
        n12521, n12520, n12519, n12518, n12517, n12516, n12515, 
        n12514, n12513, n12512, n12511, n12510, n12509, n12505, 
        n12504, n12503, n12502, n12501, n12500, n12499, n71_adj_2035, 
        n12498, n74_adj_2036, n12497, n77_adj_2037, n12496, n80_adj_2038, 
        n12495, n83_adj_2039, n12494, n86_adj_2040, n12493, n89_adj_2041, 
        n12492, n92_adj_2042, n12491, n95_adj_2043, n12490, n98_adj_2044, 
        n12489, n101_adj_2045, n12488, n104_adj_2046, n12487, n107_adj_2047, 
        n12486, n110_adj_2048, n12485, n113_adj_2049, n12484, n116_adj_2050, 
        n12483, n119_adj_2051, n12482, n122_adj_2052, n12481, n125_adj_2053, 
        n12480, n128_adj_2054, n12479, n131_adj_2055, n12478, n134_adj_2056, 
        n12477, n137_adj_2057, n12476, n140_adj_2058, n12475, n143_adj_2059, 
        n12474, n146_adj_2060, n12473, n149_adj_2061, n12472, n152_adj_2062, 
        n12471, n155_adj_2063, n12470, n158_adj_2064, n12469, n161_adj_2065, 
        n12468, n12467, n12466, n12465, n12464, n12463, n12462, 
        n12461, n12460, n12459, n12458, n12457, n12456, n12455, 
        n12454, n12453, n12452, n12451, n12450, n12449, n12448, 
        n12447, n12446, n12445, n12444, n12443, n12442, n12440, 
        n12439, n12438, n12437, n12436, n12435, n12434, n12433, 
        n12432, n12431, n12430, n12429, n12428, n12427, n12426, 
        n12425, n12421, n12420, n12419, n12418, n12417, n12416, 
        n12415, n12414, n12413, n12412, n12411, n12410, n12409, 
        n12408, n12407, n12406, n12405, n12404, n12403, n12402, 
        n68_adj_2066, n12401, n71_adj_2067, n12400, n74_adj_2068, 
        n12399, n77_adj_2069, n12398, n80_adj_2070, n12397, n83_adj_2071, 
        n12396, n86_adj_2072, n12395, n89_adj_2073, n12394, n92_adj_2074, 
        n12393, n95_adj_2075, n12392, n98_adj_2076, n12391, n101_adj_2077, 
        n104_adj_2078, n107_adj_2079, n110_adj_2080, n113_adj_2081, 
        n116_adj_2082, n119_adj_2083, n122_adj_2084, n125_adj_2085, 
        n128_adj_2086, n131_adj_2087, n134_adj_2088, n137_adj_2089, 
        n140_adj_2090, n143_adj_2091, n146_adj_2092, n149_adj_2093, 
        n152_adj_2094, n155_adj_2095, n158_adj_2096, n161_adj_2097, 
        n68_adj_2098, n71_adj_2099, n74_adj_2100, n77_adj_2101, n80_adj_2102, 
        n83_adj_2103, n86_adj_2104, n89_adj_2105, n92_adj_2106, n95_adj_2107, 
        n98_adj_2108, n101_adj_2109, n104_adj_2110, n107_adj_2111, n110_adj_2112, 
        n113_adj_2113, n116_adj_2114, n119_adj_2115, n122_adj_2116, 
        n125_adj_2117, n128_adj_2118, n131_adj_2119, n134_adj_2120, 
        n137_adj_2121, n140_adj_2122, n143_adj_2123, n146_adj_2124, 
        n149_adj_2125, n152_adj_2126, n155_adj_2127, n158_adj_2128, 
        n161_adj_2129, n68_adj_2130, n71_adj_2131, n74_adj_2132, n77_adj_2133, 
        n80_adj_2134, n83_adj_2135, n86_adj_2136, n89_adj_2137, n92_adj_2138, 
        n95_adj_2139, n98_adj_2140, n101_adj_2141, n104_adj_2142, n107_adj_2143, 
        n110_adj_2144, n113_adj_2145, n116_adj_2146, n119_adj_2147, 
        n122_adj_2148, n125_adj_2149, n128_adj_2150, n131_adj_2151, 
        n134_adj_2152, n137_adj_2153, n140_adj_2154, n143_adj_2155, 
        n146_adj_2156, n149_adj_2157, n152_adj_2158, n155_adj_2159, 
        n158_adj_2160, n161_adj_2161, n68_adj_2162, n71_adj_2163, n74_adj_2164, 
        n77_adj_2165, n80_adj_2166, n83_adj_2167, n86_adj_2168, n89_adj_2169, 
        n92_adj_2170, n95_adj_2171, n98_adj_2172, n101_adj_2173, n104_adj_2174, 
        n107_adj_2175, n110_adj_2176, n113_adj_2177, n116_adj_2178, 
        n119_adj_2179, n122_adj_2180, n125_adj_2181, n128_adj_2182, 
        n131_adj_2183, n134_adj_2184, n137_adj_2185, n140_adj_2186, 
        n143_adj_2187, n146_adj_2188, n149_adj_2189, n152_adj_2190, 
        n155_adj_2191, n158_adj_2192, n161_adj_2193, n62_adj_2194, n13836, 
        n60_adj_2195, n13835, n11713, n57_adj_2196, n55_adj_2197, 
        n54_adj_2198, n13834, n52_adj_2199, n51_adj_2200, n50_adj_2201, 
        n48_adj_2202, n13833, n42_adj_2203, n41_adj_2204, n34_adj_2205, 
        n13832, n13840, n13839, n13838, n13831, n13830, n13829, 
        n13828, n13827, n13826, n13825, n13824, n13823, n13822, 
        n13821, n13820, n13819, n13818;
    
    VHI i2 (.Z(VCC_net));
    LUT4 i1495_2_lut_4_lut (.A(n68_adj_474), .B(n68_adj_442), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n61)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1495_2_lut_4_lut.init = 16'h0035;
    FD1S3AX b1_reg_i0 (.D(b_c_0), .CK(clk_c), .Q(b1_reg[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i0.GSR = "ENABLED";
    FD1S3AX c1_reg_i0 (.D(c_c_0), .CK(clk_c), .Q(c1_reg[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i0.GSR = "ENABLED";
    FD1S3AX d1_reg_i0 (.D(d_c_0), .CK(clk_c), .Q(d1_reg[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i0.GSR = "ENABLED";
    FD1S3AX b2_reg_i0 (.D(b1_reg[0]), .CK(clk_c), .Q(b2_reg[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i0.GSR = "ENABLED";
    FD1S3AX det_q4_28_i4 (.D(det_q4_28_31__N_65[4]), .CK(clk_c), .Q(det_q4_28[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i4.GSR = "ENABLED";
    FD1S3AX c2_reg_i0 (.D(c1_reg[0]), .CK(clk_c), .Q(c2_reg[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i0.GSR = "ENABLED";
    FD1S3AX det_q4_28_i3 (.D(det_q4_28_31__N_65[3]), .CK(clk_c), .Q(det_q4_28[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i3.GSR = "ENABLED";
    CCU2C _add_1_532_add_4_25 (.A0(n95_adj_707), .B0(n13822), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_706), .B1(n13822), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12621), .COUT(n12622), .S0(n92_adj_642), 
          .S1(n89_adj_641));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_25.INJECT1_1 = "NO";
    FD1S3AY det_zero_stage2_49 (.D(det_zero_reg), .CK(clk_c), .Q(det_zero_stage2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam det_zero_stage2_49.GSR = "ENABLED";
    FD1S3AX det_q4_28_i2 (.D(det_q4_28_31__N_65[2]), .CK(clk_c), .Q(det_q4_28[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i2.GSR = "ENABLED";
    FD1S3AX det_q4_28_i1 (.D(det_q4_28_31__N_65[1]), .CK(clk_c), .Q(det_q4_28[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i1.GSR = "ENABLED";
    FD1S3AX c2_reg_i15 (.D(c1_reg[15]), .CK(clk_c), .Q(c2_reg[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i15.GSR = "ENABLED";
    FD1S3AX det_q4_28_i0 (.D(det_q4_28_31__N_65[0]), .CK(clk_c), .Q(det_q4_28[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i0.GSR = "ENABLED";
    FD1S3AX c2_reg_i14 (.D(c1_reg[14]), .CK(clk_c), .Q(c2_reg[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i14.GSR = "ENABLED";
    FD1S3AX c2_reg_i13 (.D(c1_reg[13]), .CK(clk_c), .Q(c2_reg[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i13.GSR = "ENABLED";
    FD1S3JX error_reg_54 (.D(error_recip), .CK(clk_c), .PD(det_zero_stage2), 
            .Q(error_c));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam error_reg_54.GSR = "ENABLED";
    FD1S3AY det_zero_reg_40 (.D(det_zero_reg_N_162), .CK(clk_c), .Q(det_zero_reg));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_zero_reg_40.GSR = "ENABLED";
    FD1S3AX c2_reg_i12 (.D(c1_reg[12]), .CK(clk_c), .Q(c2_reg[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i12.GSR = "ENABLED";
    FD1S3AX c2_reg_i11 (.D(c1_reg[11]), .CK(clk_c), .Q(c2_reg[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i11.GSR = "ENABLED";
    FD1S3AX c2_reg_i10 (.D(c1_reg[10]), .CK(clk_c), .Q(c2_reg[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i10.GSR = "ENABLED";
    FD1S3AX c2_reg_i9 (.D(c1_reg[9]), .CK(clk_c), .Q(c2_reg[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i9.GSR = "ENABLED";
    FD1S3AX c2_reg_i8 (.D(c1_reg[8]), .CK(clk_c), .Q(c2_reg[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i8.GSR = "ENABLED";
    OB c_inv_pad_9 (.I(c_inv_c_9), .O(c_inv[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    FD1S3AX c2_reg_i7 (.D(c1_reg[7]), .CK(clk_c), .Q(c2_reg[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i7.GSR = "ENABLED";
    FD1S3AX c2_reg_i6 (.D(c1_reg[6]), .CK(clk_c), .Q(c2_reg[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i6.GSR = "ENABLED";
    FD1S3AX c2_reg_i5 (.D(c1_reg[5]), .CK(clk_c), .Q(c2_reg[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i5.GSR = "ENABLED";
    FD1S3AX c2_reg_i4 (.D(c1_reg[4]), .CK(clk_c), .Q(c2_reg[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i4.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i1 (.D(a_inv_15__N_1[32]), .CK(clk_c), .Q(a_inv_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i1.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i1 (.D(d_inv_15__N_49[32]), .CK(clk_c), .Q(d_inv_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i1.GSR = "ENABLED";
    FD1S3AX c2_reg_i3 (.D(c1_reg[3]), .CK(clk_c), .Q(c2_reg[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i3.GSR = "ENABLED";
    FD1S3AX c2_reg_i2 (.D(c1_reg[2]), .CK(clk_c), .Q(c2_reg[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i2.GSR = "ENABLED";
    FD1S3AX c2_reg_i1 (.D(c1_reg[1]), .CK(clk_c), .Q(c2_reg[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam c2_reg_i1.GSR = "ENABLED";
    FD1S3AX b2_reg_i15 (.D(b1_reg[15]), .CK(clk_c), .Q(b2_reg[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i15.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i1 (.D(b_inv_15__N_17[32]), .CK(clk_c), .Q(b_inv_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i1.GSR = "ENABLED";
    FD1S3AX b2_reg_i14 (.D(b1_reg[14]), .CK(clk_c), .Q(b2_reg[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i14.GSR = "ENABLED";
    CCU2C _add_1_532_add_4_23 (.A0(n101_adj_709), .B0(n13822), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_708), .B1(n13822), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12620), .COUT(n12621), .S0(n98_adj_644), 
          .S1(n95_adj_643));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_23.INJECT1_1 = "NO";
    FD1S3AX b2_reg_i13 (.D(b1_reg[13]), .CK(clk_c), .Q(b2_reg[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i13.GSR = "ENABLED";
    FD1S3AX b2_reg_i12 (.D(b1_reg[12]), .CK(clk_c), .Q(b2_reg[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i12.GSR = "ENABLED";
    FD1S3AX b2_reg_i11 (.D(b1_reg[11]), .CK(clk_c), .Q(b2_reg[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i11.GSR = "ENABLED";
    FD1S3AX b2_reg_i10 (.D(b1_reg[10]), .CK(clk_c), .Q(b2_reg[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i10.GSR = "ENABLED";
    FD1S3AX b2_reg_i9 (.D(b1_reg[9]), .CK(clk_c), .Q(b2_reg[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i9.GSR = "ENABLED";
    FD1S3AX b2_reg_i8 (.D(b1_reg[8]), .CK(clk_c), .Q(b2_reg[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i8.GSR = "ENABLED";
    FD1S3AX b2_reg_i7 (.D(b1_reg[7]), .CK(clk_c), .Q(b2_reg[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i7.GSR = "ENABLED";
    FD1S3AX b2_reg_i6 (.D(b1_reg[6]), .CK(clk_c), .Q(b2_reg[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i6.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i1 (.D(c_inv_15__N_33[32]), .CK(clk_c), .Q(c_inv_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i1.GSR = "ENABLED";
    CCU2C _add_1_532_add_4_21 (.A0(n107_adj_711), .B0(n13822), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_710), .B1(n13822), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12619), .COUT(n12620), .S0(n104_adj_646), 
          .S1(n101_adj_645));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_19 (.A0(n113_adj_713), .B0(n13822), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_712), .B1(n13822), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12618), .COUT(n12619), .S0(n110_adj_648), 
          .S1(n107_adj_647));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_17 (.A0(n119_adj_715), .B0(n13822), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_714), .B1(n13822), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12617), .COUT(n12618), .S0(n116_adj_650), 
          .S1(n113_adj_649));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_15 (.A0(n125_adj_717), .B0(n13822), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_716), .B1(n13822), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12616), .COUT(n12617), .S0(n122_adj_652), 
          .S1(n119_adj_651));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_13 (.A0(n131_adj_719), .B0(n13822), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_718), .B1(n13822), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12615), .COUT(n12616), .S0(n128_adj_654), 
          .S1(n125_adj_653));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_11 (.A0(n137_adj_721), .B0(n13822), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_720), .B1(n13822), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12614), .COUT(n12615), .S0(n134_adj_656), 
          .S1(n131_adj_655));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_9 (.A0(n143_adj_723), .B0(n13822), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_722), .B1(n13822), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12613), .COUT(n12614), .S0(n140_adj_658), 
          .S1(n137_adj_657));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_7 (.A0(n149_adj_725), .B0(n13822), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_724), .B1(n13822), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12612), .COUT(n12613), .S0(n146_adj_660), 
          .S1(n143_adj_659));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_5 (.A0(n155_adj_727), .B0(n13822), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_726), .B1(n13822), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12611), .COUT(n12612), .S0(n152_adj_662), 
          .S1(n149_adj_661));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_3 (.A0(n161_adj_729), .B0(n13822), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_728), .B1(n13822), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12610), .COUT(n12611), .S0(n158_adj_664), 
          .S1(n155_adj_663));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13822), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12610), .S1(n161_adj_665));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_532_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_33 (.A0(n1444), .B0(n2583), .C0(n71_adj_1495), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12609), .S0(n68_adj_347));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_31 (.A0(n77_adj_1497), .B0(n2583), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1496), .B1(n2583), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12608), .COUT(n12609), .S0(n74_adj_349), 
          .S1(n71_adj_348));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_29 (.A0(n83_adj_1499), .B0(n2583), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1498), .B1(n2583), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12607), .COUT(n12608), .S0(n80_adj_351), 
          .S1(n77_adj_350));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_27 (.A0(n89_adj_1501), .B0(n2583), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1500), .B1(n2583), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12606), .COUT(n12607), .S0(n86_adj_353), 
          .S1(n83_adj_352));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_25 (.A0(n95_adj_1503), .B0(n2583), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1502), .B1(n2583), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12605), .COUT(n12606), .S0(n92_adj_355), 
          .S1(n89_adj_354));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_23 (.A0(n101_adj_1505), .B0(n2583), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1504), .B1(n2583), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12604), .COUT(n12605), .S0(n98_adj_357), 
          .S1(n95_adj_356));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_21 (.A0(n107_adj_1507), .B0(n2583), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1506), .B1(n2583), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12603), .COUT(n12604), .S0(n104_adj_359), 
          .S1(n101_adj_358));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_add_4_21.INJECT1_1 = "NO";
    FD1S3AX d2_reg_15__I_0_e2__i1 (.D(d1_reg[0]), .CK(clk_c), .Q(n130_adj_231));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i1.GSR = "ENABLED";
    CCU2C _add_1_add_4_19 (.A0(n113_adj_1509), .B0(n2583), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1508), .B1(n2583), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12602), .COUT(n12603), .S0(n110_adj_361), 
          .S1(n107_adj_360));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_17 (.A0(n119_adj_1511), .B0(n2583), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1510), .B1(n2583), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12601), .COUT(n12602), .S0(n116_adj_363), 
          .S1(n113_adj_362));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_15 (.A0(n125_adj_1513), .B0(n2583), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1512), .B1(n2583), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12600), .COUT(n12601), .S0(n122_adj_365), 
          .S1(n119_adj_364));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_13 (.A0(n131_adj_1515), .B0(n2583), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1514), .B1(n2583), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12599), .COUT(n12600), .S0(n128_adj_367), 
          .S1(n125_adj_366));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_11 (.A0(n137_adj_1517), .B0(n2583), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1516), .B1(n2583), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12598), .COUT(n12599), .S0(n134_adj_369), 
          .S1(n131_adj_368));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_add_4_11.INJECT1_1 = "NO";
    FD1S3AX b2_reg_i5 (.D(b1_reg[5]), .CK(clk_c), .Q(b2_reg[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i5.GSR = "ENABLED";
    FD1S3AX b2_reg_i4 (.D(b1_reg[4]), .CK(clk_c), .Q(b2_reg[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i4.GSR = "ENABLED";
    FD1S3AX b2_reg_i3 (.D(b1_reg[3]), .CK(clk_c), .Q(b2_reg[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i3.GSR = "ENABLED";
    FD1S3AX b2_reg_i2 (.D(b1_reg[2]), .CK(clk_c), .Q(b2_reg[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i2.GSR = "ENABLED";
    FD1S3AX b2_reg_i1 (.D(b1_reg[1]), .CK(clk_c), .Q(b2_reg[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(76[18] 82[12])
    defparam b2_reg_i1.GSR = "ENABLED";
    FD1S3AX d1_reg_i15 (.D(d_c_15), .CK(clk_c), .Q(d1_reg[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i15.GSR = "ENABLED";
    FD1S3AX d1_reg_i14 (.D(d_c_14), .CK(clk_c), .Q(d1_reg[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i14.GSR = "ENABLED";
    FD1S3AX d1_reg_i13 (.D(d_c_13), .CK(clk_c), .Q(d1_reg[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i13.GSR = "ENABLED";
    FD1S3AX d1_reg_i12 (.D(d_c_12), .CK(clk_c), .Q(d1_reg[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i12.GSR = "ENABLED";
    FD1S3AX d1_reg_i11 (.D(d_c_11), .CK(clk_c), .Q(d1_reg[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i11.GSR = "ENABLED";
    FD1S3AX d1_reg_i10 (.D(d_c_10), .CK(clk_c), .Q(d1_reg[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i10.GSR = "ENABLED";
    FD1S3AX d1_reg_i9 (.D(d_c_9), .CK(clk_c), .Q(d1_reg[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i9.GSR = "ENABLED";
    FD1S3AX d1_reg_i8 (.D(d_c_8), .CK(clk_c), .Q(d1_reg[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i8.GSR = "ENABLED";
    FD1S3AX d1_reg_i7 (.D(d_c_7), .CK(clk_c), .Q(d1_reg[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i7.GSR = "ENABLED";
    FD1S3AX d1_reg_i6 (.D(d_c_6), .CK(clk_c), .Q(d1_reg[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i6.GSR = "ENABLED";
    FD1S3AX d1_reg_i5 (.D(d_c_5), .CK(clk_c), .Q(d1_reg[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i5.GSR = "ENABLED";
    FD1S3AX d1_reg_i4 (.D(d_c_4), .CK(clk_c), .Q(d1_reg[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i4.GSR = "ENABLED";
    FD1S3AX d1_reg_i3 (.D(d_c_3), .CK(clk_c), .Q(d1_reg[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i3.GSR = "ENABLED";
    FD1S3AX d1_reg_i2 (.D(d_c_2), .CK(clk_c), .Q(d1_reg[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i2.GSR = "ENABLED";
    FD1S3AX d1_reg_i1 (.D(d_c_1), .CK(clk_c), .Q(d1_reg[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam d1_reg_i1.GSR = "ENABLED";
    MULT18X18D mult_3 (.A17(d_c_15), .A16(d_c_15), .A15(d_c_15), .A14(d_c_14), 
            .A13(d_c_13), .A12(d_c_12), .A11(d_c_11), .A10(d_c_10), 
            .A9(d_c_9), .A8(d_c_8), .A7(d_c_7), .A6(d_c_6), .A5(d_c_5), 
            .A4(d_c_4), .A3(d_c_3), .A2(d_c_2), .A1(d_c_1), .A0(d_c_0), 
            .B17(a_c_15), .B16(a_c_15), .B15(a_c_15), .B14(a_c_14), 
            .B13(a_c_13), .B12(a_c_12), .B11(a_c_11), .B10(a_c_10), 
            .B9(a_c_9), .B8(a_c_8), .B7(a_c_7), .B6(a_c_6), .B5(a_c_5), 
            .B4(a_c_4), .B3(a_c_3), .B2(a_c_2), .B1(a_c_1), .B0(a_c_0), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P31(det_q4_28_31__N_97[31]), 
            .P30(det_q4_28_31__N_97[30]), .P29(det_q4_28_31__N_97[29]), 
            .P28(det_q4_28_31__N_97[28]), .P27(det_q4_28_31__N_97[27]), 
            .P26(det_q4_28_31__N_97[26]), .P25(det_q4_28_31__N_97[25]), 
            .P24(det_q4_28_31__N_97[24]), .P23(det_q4_28_31__N_97[23]), 
            .P22(det_q4_28_31__N_97[22]), .P21(det_q4_28_31__N_97[21]), 
            .P20(det_q4_28_31__N_97[20]), .P19(det_q4_28_31__N_97[19]), 
            .P18(det_q4_28_31__N_97[18]), .P17(det_q4_28_31__N_97[17]), 
            .P16(det_q4_28_31__N_97[16]), .P15(det_q4_28_31__N_97[15]), 
            .P14(det_q4_28_31__N_97[14]), .P13(det_q4_28_31__N_97[13]), 
            .P12(det_q4_28_31__N_97[12]), .P11(det_q4_28_31__N_97[11]), 
            .P10(det_q4_28_31__N_97[10]), .P9(det_q4_28_31__N_97[9]), .P8(det_q4_28_31__N_97[8]), 
            .P7(det_q4_28_31__N_97[7]), .P6(det_q4_28_31__N_97[6]), .P5(det_q4_28_31__N_97[5]), 
            .P4(det_q4_28_31__N_97[4]), .P3(det_q4_28_31__N_97[3]), .P2(det_q4_28_31__N_97[2]), 
            .P1(det_q4_28_31__N_97[1]), .P0(det_q4_28_31__N_97[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:33])
    defparam mult_3.REG_INPUTA_CLK = "NONE";
    defparam mult_3.REG_INPUTA_CE = "CE0";
    defparam mult_3.REG_INPUTA_RST = "RST0";
    defparam mult_3.REG_INPUTB_CLK = "NONE";
    defparam mult_3.REG_INPUTB_CE = "CE0";
    defparam mult_3.REG_INPUTB_RST = "RST0";
    defparam mult_3.REG_INPUTC_CLK = "NONE";
    defparam mult_3.REG_INPUTC_CE = "CE0";
    defparam mult_3.REG_INPUTC_RST = "RST0";
    defparam mult_3.REG_PIPELINE_CLK = "NONE";
    defparam mult_3.REG_PIPELINE_CE = "CE0";
    defparam mult_3.REG_PIPELINE_RST = "RST0";
    defparam mult_3.REG_OUTPUT_CLK = "NONE";
    defparam mult_3.REG_OUTPUT_CE = "CE0";
    defparam mult_3.REG_OUTPUT_RST = "RST0";
    defparam mult_3.CLK0_DIV = "ENABLED";
    defparam mult_3.CLK1_DIV = "ENABLED";
    defparam mult_3.CLK2_DIV = "ENABLED";
    defparam mult_3.CLK3_DIV = "ENABLED";
    defparam mult_3.HIGHSPEED_CLK = "NONE";
    defparam mult_3.GSR = "DISABLED";
    defparam mult_3.CAS_MATCH_REG = "FALSE";
    defparam mult_3.SOURCEB_MODE = "B_SHIFT";
    defparam mult_3.MULT_BYPASS = "DISABLED";
    defparam mult_3.RESETMODE = "SYNC";
    FD1S3AX c1_reg_i15 (.D(c_c_15), .CK(clk_c), .Q(c1_reg[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i15.GSR = "ENABLED";
    MULT18X18D mult_4 (.A17(c_c_15), .A16(c_c_15), .A15(c_c_15), .A14(c_c_14), 
            .A13(c_c_13), .A12(c_c_12), .A11(c_c_11), .A10(c_c_10), 
            .A9(c_c_9), .A8(c_c_8), .A7(c_c_7), .A6(c_c_6), .A5(c_c_5), 
            .A4(c_c_4), .A3(c_c_3), .A2(c_c_2), .A1(c_c_1), .A0(c_c_0), 
            .B17(b_c_15), .B16(b_c_15), .B15(b_c_15), .B14(b_c_14), 
            .B13(b_c_13), .B12(b_c_12), .B11(b_c_11), .B10(b_c_10), 
            .B9(b_c_9), .B8(b_c_8), .B7(b_c_7), .B6(b_c_6), .B5(b_c_5), 
            .B4(b_c_4), .B3(b_c_3), .B2(b_c_2), .B1(b_c_1), .B0(b_c_0), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P31(det_q4_28_31__N_129[31]), 
            .P30(det_q4_28_31__N_129[30]), .P29(det_q4_28_31__N_129[29]), 
            .P28(det_q4_28_31__N_129[28]), .P27(det_q4_28_31__N_129[27]), 
            .P26(det_q4_28_31__N_129[26]), .P25(det_q4_28_31__N_129[25]), 
            .P24(det_q4_28_31__N_129[24]), .P23(det_q4_28_31__N_129[23]), 
            .P22(det_q4_28_31__N_129[22]), .P21(det_q4_28_31__N_129[21]), 
            .P20(det_q4_28_31__N_129[20]), .P19(det_q4_28_31__N_129[19]), 
            .P18(det_q4_28_31__N_129[18]), .P17(det_q4_28_31__N_129[17]), 
            .P16(det_q4_28_31__N_129[16]), .P15(det_q4_28_31__N_129[15]), 
            .P14(det_q4_28_31__N_129[14]), .P13(det_q4_28_31__N_129[13]), 
            .P12(det_q4_28_31__N_129[12]), .P11(det_q4_28_31__N_129[11]), 
            .P10(det_q4_28_31__N_129[10]), .P9(det_q4_28_31__N_129[9]), 
            .P8(det_q4_28_31__N_129[8]), .P7(det_q4_28_31__N_129[7]), .P6(det_q4_28_31__N_129[6]), 
            .P5(det_q4_28_31__N_129[5]), .P4(det_q4_28_31__N_129[4]), .P3(det_q4_28_31__N_129[3]), 
            .P2(det_q4_28_31__N_129[2]), .P1(det_q4_28_31__N_129[1]), .P0(det_q4_28_31__N_129[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[36:43])
    defparam mult_4.REG_INPUTA_CLK = "NONE";
    defparam mult_4.REG_INPUTA_CE = "CE0";
    defparam mult_4.REG_INPUTA_RST = "RST0";
    defparam mult_4.REG_INPUTB_CLK = "NONE";
    defparam mult_4.REG_INPUTB_CE = "CE0";
    defparam mult_4.REG_INPUTB_RST = "RST0";
    defparam mult_4.REG_INPUTC_CLK = "NONE";
    defparam mult_4.REG_INPUTC_CE = "CE0";
    defparam mult_4.REG_INPUTC_RST = "RST0";
    defparam mult_4.REG_PIPELINE_CLK = "NONE";
    defparam mult_4.REG_PIPELINE_CE = "CE0";
    defparam mult_4.REG_PIPELINE_RST = "RST0";
    defparam mult_4.REG_OUTPUT_CLK = "NONE";
    defparam mult_4.REG_OUTPUT_CE = "CE0";
    defparam mult_4.REG_OUTPUT_RST = "RST0";
    defparam mult_4.CLK0_DIV = "ENABLED";
    defparam mult_4.CLK1_DIV = "ENABLED";
    defparam mult_4.CLK2_DIV = "ENABLED";
    defparam mult_4.CLK3_DIV = "ENABLED";
    defparam mult_4.HIGHSPEED_CLK = "NONE";
    defparam mult_4.GSR = "DISABLED";
    defparam mult_4.CAS_MATCH_REG = "FALSE";
    defparam mult_4.SOURCEB_MODE = "B_SHIFT";
    defparam mult_4.MULT_BYPASS = "DISABLED";
    defparam mult_4.RESETMODE = "SYNC";
    FD1S3AX c1_reg_i14 (.D(c_c_14), .CK(clk_c), .Q(c1_reg[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i14.GSR = "ENABLED";
    ALU54B lat_alu_19 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n11483), .SIGNEDIB(n11556), .SIGNEDCIN(n11629), .A35(n11482), 
           .A34(n11481), .A33(n11480), .A32(n11479), .A31(n11478), .A30(n11477), 
           .A29(n11476), .A28(n11475), .A27(n11474), .A26(n11473), .A25(n11472), 
           .A24(n11471), .A23(n11470), .A22(n11469), .A21(n11468), .A20(n11467), 
           .A19(n11466), .A18(n11465), .A17(n11464), .A16(n11463), .A15(n11462), 
           .A14(n11461), .A13(n11460), .A12(n11459), .A11(n11458), .A10(n11457), 
           .A9(n11456), .A8(n11455), .A7(n11454), .A6(n11453), .A5(n11452), 
           .A4(n11451), .A3(n11450), .A2(n11449), .A1(n11448), .A0(n11447), 
           .B35(n11555), .B34(n11554), .B33(n11553), .B32(n11552), .B31(n11551), 
           .B30(n11550), .B29(n11549), .B28(n11548), .B27(n11547), .B26(n11546), 
           .B25(n11545), .B24(n11544), .B23(n11543), .B22(n11542), .B21(n11541), 
           .B20(n11540), .B19(n11539), .B18(n11538), .B17(n11537), .B16(n11536), 
           .B15(n11535), .B14(n11534), .B13(n11533), .B12(n11532), .B11(n11531), 
           .B10(n11530), .B9(n11529), .B8(n11528), .B7(n11527), .B6(n11526), 
           .B5(n11525), .B4(n11524), .B3(n11523), .B2(n11522), .B1(n11521), 
           .B0(n11520), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n11519), .MA34(n11518), .MA33(n11517), .MA32(n11516), 
           .MA31(n11515), .MA30(n11514), .MA29(n11513), .MA28(n11512), 
           .MA27(n11511), .MA26(n11510), .MA25(n11509), .MA24(n11508), 
           .MA23(n11507), .MA22(n11506), .MA21(n11505), .MA20(n11504), 
           .MA19(n11503), .MA18(n11502), .MA17(n11501), .MA16(n11500), 
           .MA15(n11499), .MA14(n11498), .MA13(n11497), .MA12(n11496), 
           .MA11(n11495), .MA10(n11494), .MA9(n11493), .MA8(n11492), 
           .MA7(n11491), .MA6(n11490), .MA5(n11489), .MA4(n11488), .MA3(n11487), 
           .MA2(n11486), .MA1(n11485), .MA0(n11484), .MB35(n11592), 
           .MB34(n11591), .MB33(n11590), .MB32(n11589), .MB31(n11588), 
           .MB30(n11587), .MB29(n11586), .MB28(n11585), .MB27(n11584), 
           .MB26(n11583), .MB25(n11582), .MB24(n11581), .MB23(n11580), 
           .MB22(n11579), .MB21(n11578), .MB20(n11577), .MB19(n11576), 
           .MB18(n11575), .MB17(n11574), .MB16(n11573), .MB15(n11572), 
           .MB14(n11571), .MB13(n11570), .MB12(n11569), .MB11(n11568), 
           .MB10(n11567), .MB9(n11566), .MB8(n11565), .MB7(n11564), 
           .MB6(n11563), .MB5(n11562), .MB4(n11561), .MB3(n11560), .MB2(n11559), 
           .MB1(n11558), .MB0(n11557), .CIN53(n11628), .CIN52(n11627), 
           .CIN51(n11626), .CIN50(n11625), .CIN49(n11624), .CIN48(n11623), 
           .CIN47(n11622), .CIN46(n11621), .CIN45(n11620), .CIN44(n11619), 
           .CIN43(n11618), .CIN42(n11617), .CIN41(n11616), .CIN40(n11615), 
           .CIN39(n11614), .CIN38(n11613), .CIN37(n11612), .CIN36(n11611), 
           .CIN35(n11610), .CIN34(n11609), .CIN33(n11608), .CIN32(n11607), 
           .CIN31(n11606), .CIN30(n11605), .CIN29(n11604), .CIN28(n11603), 
           .CIN27(n11602), .CIN26(n11601), .CIN25(n11600), .CIN24(n11599), 
           .CIN23(n11598), .CIN22(n11597), .CIN21(n11596), .CIN20(n11595), 
           .CIN19(n11594), .CIN18(n11593), .CIN17(prod_d[17]), .CIN16(prod_d[16]), 
           .CIN15(prod_d[15]), .CIN14(n11286), .CIN13(n11287), .CIN12(n11288), 
           .CIN11(n11289), .CIN10(n11290), .CIN9(n11291), .CIN8(n11292), 
           .CIN7(n11293), .CIN6(n11294), .CIN5(n11295), .CIN4(n11296), 
           .CIN3(n11297), .CIN2(n11298), .CIN1(n11299), .CIN0(n11300), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R29(prod_d[47]), 
           .R28(prod_d[46]), .R27(prod_d[45]), .R26(prod_d[44]), .R25(prod_d[43]), 
           .R24(prod_d[42]), .R23(prod_d[41]), .R22(prod_d[40]), .R21(prod_d[39]), 
           .R20(prod_d[38]), .R19(prod_d[37]), .R18(prod_d[36]), .R17(prod_d[35]), 
           .R16(prod_d[34]), .R15(prod_d[33]), .R14(prod_d[32]), .R13(prod_d[31]), 
           .R12(prod_d[30]), .R11(prod_d[29]), .R10(prod_d[28]), .R9(prod_d[27]), 
           .R8(prod_d[26]), .R7(prod_d[25]), .R6(prod_d[24]), .R5(prod_d[23]), 
           .R4(prod_d[22]), .R3(prod_d[21]), .R2(prod_d[20]), .R1(prod_d[19]), 
           .R0(prod_d[18]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam lat_alu_19.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_19.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_19.REG_FLAG_CLK = "NONE";
    defparam lat_alu_19.REG_FLAG_CE = "CE0";
    defparam lat_alu_19.REG_FLAG_RST = "RST0";
    defparam lat_alu_19.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASK01 = "0x00000000000000";
    defparam lat_alu_19.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_19.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_19.CLK0_DIV = "ENABLED";
    defparam lat_alu_19.CLK1_DIV = "ENABLED";
    defparam lat_alu_19.CLK2_DIV = "ENABLED";
    defparam lat_alu_19.CLK3_DIV = "ENABLED";
    defparam lat_alu_19.MCPAT = "0x00000000000000";
    defparam lat_alu_19.MASKPAT = "0x00000000000000";
    defparam lat_alu_19.RNDPAT = "0x00000000000000";
    defparam lat_alu_19.GSR = "DISABLED";
    defparam lat_alu_19.RESETMODE = "SYNC";
    defparam lat_alu_19.MULT9_MODE = "DISABLED";
    defparam lat_alu_19.LEGACY = "DISABLED";
    FD1S3AX a2_reg_15__I_0_e2__i1 (.D(a1_reg[0]), .CK(clk_c), .Q(n130));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i1.GSR = "ENABLED";
    ALU54B lat_alu_18 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n11337), .SIGNEDIB(n11410), .SIGNEDCIN(GND_net), 
           .A35(n11336), .A34(n11335), .A33(n11334), .A32(n11333), .A31(n11332), 
           .A30(n11331), .A29(n11330), .A28(n11329), .A27(n11328), .A26(n11327), 
           .A25(n11326), .A24(n11325), .A23(n11324), .A22(n11323), .A21(n11322), 
           .A20(n11321), .A19(n11320), .A18(n11319), .A17(n11318), .A16(n11317), 
           .A15(n11316), .A14(n11315), .A13(n11314), .A12(n11313), .A11(n11312), 
           .A10(n11311), .A9(n11310), .A8(n11309), .A7(n11308), .A6(n11307), 
           .A5(n11306), .A4(n11305), .A3(n11304), .A2(n11303), .A1(n11302), 
           .A0(n11301), .B35(n11409), .B34(n11408), .B33(n11407), .B32(n11406), 
           .B31(n11405), .B30(n11404), .B29(n11403), .B28(n11402), .B27(n11401), 
           .B26(n11400), .B25(n11399), .B24(n11398), .B23(n11397), .B22(n11396), 
           .B21(n11395), .B20(n11394), .B19(n11393), .B18(n11392), .B17(n11391), 
           .B16(n11390), .B15(n11389), .B14(n11388), .B13(n11387), .B12(n11386), 
           .B11(n11385), .B10(n11384), .B9(n11383), .B8(n11382), .B7(n11381), 
           .B6(n11380), .B5(n11379), .B4(n11378), .B3(n11377), .B2(n11376), 
           .B1(n11375), .B0(n11374), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n11373), .MA34(n11372), .MA33(n11371), .MA32(n11370), 
           .MA31(n11369), .MA30(n11368), .MA29(n11367), .MA28(n11366), 
           .MA27(n11365), .MA26(n11364), .MA25(n11363), .MA24(n11362), 
           .MA23(n11361), .MA22(n11360), .MA21(n11359), .MA20(n11358), 
           .MA19(n11357), .MA18(n11356), .MA17(n11355), .MA16(n11354), 
           .MA15(n11353), .MA14(n11352), .MA13(n11351), .MA12(n11350), 
           .MA11(n11349), .MA10(n11348), .MA9(n11347), .MA8(n11346), 
           .MA7(n11345), .MA6(n11344), .MA5(n11343), .MA4(n11342), .MA3(n11341), 
           .MA2(n11340), .MA1(n11339), .MA0(n11338), .MB35(n11446), 
           .MB34(n11445), .MB33(n11444), .MB32(n11443), .MB31(n11442), 
           .MB30(n11441), .MB29(n11440), .MB28(n11439), .MB27(n11438), 
           .MB26(n11437), .MB25(n11436), .MB24(n11435), .MB23(n11434), 
           .MB22(n11433), .MB21(n11432), .MB20(n11431), .MB19(n11430), 
           .MB18(n11429), .MB17(n11428), .MB16(n11427), .MB15(n11426), 
           .MB14(n11425), .MB13(n11424), .MB12(n11423), .MB11(n11422), 
           .MB10(n11421), .MB9(n11420), .MB8(n11419), .MB7(n11418), 
           .MB6(n11417), .MB5(n11416), .MB4(n11415), .MB3(n11414), .MB2(n11413), 
           .MB1(n11412), .MB0(n11411), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n11628), 
           .R52(n11627), .R51(n11626), .R50(n11625), .R49(n11624), .R48(n11623), 
           .R47(n11622), .R46(n11621), .R45(n11620), .R44(n11619), .R43(n11618), 
           .R42(n11617), .R41(n11616), .R40(n11615), .R39(n11614), .R38(n11613), 
           .R37(n11612), .R36(n11611), .R35(n11610), .R34(n11609), .R33(n11608), 
           .R32(n11607), .R31(n11606), .R30(n11605), .R29(n11604), .R28(n11603), 
           .R27(n11602), .R26(n11601), .R25(n11600), .R24(n11599), .R23(n11598), 
           .R22(n11597), .R21(n11596), .R20(n11595), .R19(n11594), .R18(n11593), 
           .R17(prod_d[17]), .R16(prod_d[16]), .R15(prod_d[15]), .R14(n11286), 
           .R13(n11287), .R12(n11288), .R11(n11289), .R10(n11290), .R9(n11291), 
           .R8(n11292), .R7(n11293), .R6(n11294), .R5(n11295), .R4(n11296), 
           .R3(n11297), .R2(n11298), .R1(n11299), .R0(n11300), .SIGNEDR(n11629));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam lat_alu_18.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_18.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_18.REG_FLAG_CLK = "NONE";
    defparam lat_alu_18.REG_FLAG_CE = "CE0";
    defparam lat_alu_18.REG_FLAG_RST = "RST0";
    defparam lat_alu_18.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASK01 = "0x00000000000000";
    defparam lat_alu_18.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_18.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_18.CLK0_DIV = "ENABLED";
    defparam lat_alu_18.CLK1_DIV = "ENABLED";
    defparam lat_alu_18.CLK2_DIV = "ENABLED";
    defparam lat_alu_18.CLK3_DIV = "ENABLED";
    defparam lat_alu_18.MCPAT = "0x00000000000000";
    defparam lat_alu_18.MASKPAT = "0x00000000000000";
    defparam lat_alu_18.RNDPAT = "0x00000000000000";
    defparam lat_alu_18.GSR = "DISABLED";
    defparam lat_alu_18.RESETMODE = "SYNC";
    defparam lat_alu_18.MULT9_MODE = "DISABLED";
    defparam lat_alu_18.LEGACY = "DISABLED";
    FD1S3AX c1_reg_i13 (.D(c_c_13), .CK(clk_c), .Q(c1_reg[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i13.GSR = "ENABLED";
    MULT18X18D lat_mult_17 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68), .B16(n68), .B15(n68), 
            .B14(n68), .B13(n68), .B12(n68), .B11(n68), .B10(n68), 
            .B9(n68), .B8(n68), .B7(n68), .B6(n68), .B5(n68), .B4(n68), 
            .B3(n68), .B2(n68), .B1(n68), .B0(n68), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n11537), .ROA16(n11536), .ROA15(n11535), 
            .ROA14(n11534), .ROA13(n11533), .ROA12(n11532), .ROA11(n11531), 
            .ROA10(n11530), .ROA9(n11529), .ROA8(n11528), .ROA7(n11527), 
            .ROA6(n11526), .ROA5(n11525), .ROA4(n11524), .ROA3(n11523), 
            .ROA2(n11522), .ROA1(n11521), .ROA0(n11520), .ROB17(n11555), 
            .ROB16(n11554), .ROB15(n11553), .ROB14(n11552), .ROB13(n11551), 
            .ROB12(n11550), .ROB11(n11549), .ROB10(n11548), .ROB9(n11547), 
            .ROB8(n11546), .ROB7(n11545), .ROB6(n11544), .ROB5(n11543), 
            .ROB4(n11542), .ROB3(n11541), .ROB2(n11540), .ROB1(n11539), 
            .ROB0(n11538), .P35(n11592), .P34(n11591), .P33(n11590), 
            .P32(n11589), .P31(n11588), .P30(n11587), .P29(n11586), 
            .P28(n11585), .P27(n11584), .P26(n11583), .P25(n11582), 
            .P24(n11581), .P23(n11580), .P22(n11579), .P21(n11578), 
            .P20(n11577), .P19(n11576), .P18(n11575), .P17(n11574), 
            .P16(n11573), .P15(n11572), .P14(n11571), .P13(n11570), 
            .P12(n11569), .P11(n11568), .P10(n11567), .P9(n11566), .P8(n11565), 
            .P7(n11564), .P6(n11563), .P5(n11562), .P4(n11561), .P3(n11560), 
            .P2(n11559), .P1(n11558), .P0(n11557), .SIGNEDP(n11556));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam lat_mult_17.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_17.REG_INPUTA_CE = "CE3";
    defparam lat_mult_17.REG_INPUTA_RST = "RST3";
    defparam lat_mult_17.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTB_CE = "CE0";
    defparam lat_mult_17.REG_INPUTB_RST = "RST0";
    defparam lat_mult_17.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTC_CE = "CE0";
    defparam lat_mult_17.REG_INPUTC_RST = "RST0";
    defparam lat_mult_17.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_17.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_17.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_17.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_17.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_17.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_17.CLK0_DIV = "ENABLED";
    defparam lat_mult_17.CLK1_DIV = "ENABLED";
    defparam lat_mult_17.CLK2_DIV = "ENABLED";
    defparam lat_mult_17.CLK3_DIV = "ENABLED";
    defparam lat_mult_17.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_17.GSR = "DISABLED";
    defparam lat_mult_17.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_17.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_17.MULT_BYPASS = "DISABLED";
    defparam lat_mult_17.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i12 (.D(c_c_12), .CK(clk_c), .Q(c1_reg[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i12.GSR = "ENABLED";
    MULT18X18D lat_mult_16 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(n68), .B16(n68), .B15(n68), 
            .B14(n68), .B13(n68), .B12(n68), .B11(n68), .B10(n68), 
            .B9(n68), .B8(n68), .B7(n68), .B6(n68), .B5(n68), .B4(n68), 
            .B3(n68), .B2(n68), .B1(n68), .B0(n68), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n11464), .ROA16(n11463), .ROA15(n11462), 
            .ROA14(n11461), .ROA13(n11460), .ROA12(n11459), .ROA11(n11458), 
            .ROA10(n11457), .ROA9(n11456), .ROA8(n11455), .ROA7(n11454), 
            .ROA6(n11453), .ROA5(n11452), .ROA4(n11451), .ROA3(n11450), 
            .ROA2(n11449), .ROA1(n11448), .ROA0(n11447), .ROB17(n11482), 
            .ROB16(n11481), .ROB15(n11480), .ROB14(n11479), .ROB13(n11478), 
            .ROB12(n11477), .ROB11(n11476), .ROB10(n11475), .ROB9(n11474), 
            .ROB8(n11473), .ROB7(n11472), .ROB6(n11471), .ROB5(n11470), 
            .ROB4(n11469), .ROB3(n11468), .ROB2(n11467), .ROB1(n11466), 
            .ROB0(n11465), .P35(n11519), .P34(n11518), .P33(n11517), 
            .P32(n11516), .P31(n11515), .P30(n11514), .P29(n11513), 
            .P28(n11512), .P27(n11511), .P26(n11510), .P25(n11509), 
            .P24(n11508), .P23(n11507), .P22(n11506), .P21(n11505), 
            .P20(n11504), .P19(n11503), .P18(n11502), .P17(n11501), 
            .P16(n11500), .P15(n11499), .P14(n11498), .P13(n11497), 
            .P12(n11496), .P11(n11495), .P10(n11494), .P9(n11493), .P8(n11492), 
            .P7(n11491), .P6(n11490), .P5(n11489), .P4(n11488), .P3(n11487), 
            .P2(n11486), .P1(n11485), .P0(n11484), .SIGNEDP(n11483));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam lat_mult_16.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_16.REG_INPUTA_CE = "CE3";
    defparam lat_mult_16.REG_INPUTA_RST = "RST3";
    defparam lat_mult_16.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTB_CE = "CE0";
    defparam lat_mult_16.REG_INPUTB_RST = "RST0";
    defparam lat_mult_16.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTC_CE = "CE0";
    defparam lat_mult_16.REG_INPUTC_RST = "RST0";
    defparam lat_mult_16.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_16.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_16.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_16.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_16.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_16.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_16.CLK0_DIV = "ENABLED";
    defparam lat_mult_16.CLK1_DIV = "ENABLED";
    defparam lat_mult_16.CLK2_DIV = "ENABLED";
    defparam lat_mult_16.CLK3_DIV = "ENABLED";
    defparam lat_mult_16.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_16.GSR = "DISABLED";
    defparam lat_mult_16.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_16.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_16.MULT_BYPASS = "DISABLED";
    defparam lat_mult_16.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i11 (.D(c_c_11), .CK(clk_c), .Q(c1_reg[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i11.GSR = "ENABLED";
    MULT18X18D lat_mult_15 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68), .B16(n68), .B15(n68), 
            .B14(n102), .B13(n104), .B12(n106), .B11(n108), .B10(n110), 
            .B9(n112), .B8(n114), .B7(n116), .B6(n118), .B5(n120), 
            .B4(n122), .B3(n124), .B2(n126), .B1(n128), .B0(n130), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n11391), .ROA16(n11390), 
            .ROA15(n11389), .ROA14(n11388), .ROA13(n11387), .ROA12(n11386), 
            .ROA11(n11385), .ROA10(n11384), .ROA9(n11383), .ROA8(n11382), 
            .ROA7(n11381), .ROA6(n11380), .ROA5(n11379), .ROA4(n11378), 
            .ROA3(n11377), .ROA2(n11376), .ROA1(n11375), .ROA0(n11374), 
            .ROB17(n11409), .ROB16(n11408), .ROB15(n11407), .ROB14(n11406), 
            .ROB13(n11405), .ROB12(n11404), .ROB11(n11403), .ROB10(n11402), 
            .ROB9(n11401), .ROB8(n11400), .ROB7(n11399), .ROB6(n11398), 
            .ROB5(n11397), .ROB4(n11396), .ROB3(n11395), .ROB2(n11394), 
            .ROB1(n11393), .ROB0(n11392), .P35(n11446), .P34(n11445), 
            .P33(n11444), .P32(n11443), .P31(n11442), .P30(n11441), 
            .P29(n11440), .P28(n11439), .P27(n11438), .P26(n11437), 
            .P25(n11436), .P24(n11435), .P23(n11434), .P22(n11433), 
            .P21(n11432), .P20(n11431), .P19(n11430), .P18(n11429), 
            .P17(n11428), .P16(n11427), .P15(n11426), .P14(n11425), 
            .P13(n11424), .P12(n11423), .P11(n11422), .P10(n11421), 
            .P9(n11420), .P8(n11419), .P7(n11418), .P6(n11417), .P5(n11416), 
            .P4(n11415), .P3(n11414), .P2(n11413), .P1(n11412), .P0(n11411), 
            .SIGNEDP(n11410));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam lat_mult_15.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_15.REG_INPUTA_CE = "CE3";
    defparam lat_mult_15.REG_INPUTA_RST = "RST3";
    defparam lat_mult_15.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTB_CE = "CE0";
    defparam lat_mult_15.REG_INPUTB_RST = "RST0";
    defparam lat_mult_15.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTC_CE = "CE0";
    defparam lat_mult_15.REG_INPUTC_RST = "RST0";
    defparam lat_mult_15.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_15.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_15.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_15.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_15.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_15.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_15.CLK0_DIV = "ENABLED";
    defparam lat_mult_15.CLK1_DIV = "ENABLED";
    defparam lat_mult_15.CLK2_DIV = "ENABLED";
    defparam lat_mult_15.CLK3_DIV = "ENABLED";
    defparam lat_mult_15.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_15.GSR = "DISABLED";
    defparam lat_mult_15.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_15.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_15.MULT_BYPASS = "DISABLED";
    defparam lat_mult_15.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i10 (.D(c_c_10), .CK(clk_c), .Q(c1_reg[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i10.GSR = "ENABLED";
    MULT18X18D a2_reg_15__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), 
            .A14(n50), .A13(n51), .A12(n52), .A11(n53), .A10(n54), 
            .A9(n55), .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), 
            .A3(n61), .A2(n62), .A1(n63), .A0(n64), .B17(n68), .B16(n68), 
            .B15(n68), .B14(n102), .B13(n104), .B12(n106), .B11(n108), 
            .B10(n110), .B9(n112), .B8(n114), .B7(n116), .B6(n118), 
            .B5(n120), .B4(n122), .B3(n124), .B2(n126), .B1(n128), 
            .B0(n130), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n11318), 
            .ROA16(n11317), .ROA15(n11316), .ROA14(n11315), .ROA13(n11314), 
            .ROA12(n11313), .ROA11(n11312), .ROA10(n11311), .ROA9(n11310), 
            .ROA8(n11309), .ROA7(n11308), .ROA6(n11307), .ROA5(n11306), 
            .ROA4(n11305), .ROA3(n11304), .ROA2(n11303), .ROA1(n11302), 
            .ROA0(n11301), .ROB17(n11336), .ROB16(n11335), .ROB15(n11334), 
            .ROB14(n11333), .ROB13(n11332), .ROB12(n11331), .ROB11(n11330), 
            .ROB10(n11329), .ROB9(n11328), .ROB8(n11327), .ROB7(n11326), 
            .ROB6(n11325), .ROB5(n11324), .ROB4(n11323), .ROB3(n11322), 
            .ROB2(n11321), .ROB1(n11320), .ROB0(n11319), .P35(n11373), 
            .P34(n11372), .P33(n11371), .P32(n11370), .P31(n11369), 
            .P30(n11368), .P29(n11367), .P28(n11366), .P27(n11365), 
            .P26(n11364), .P25(n11363), .P24(n11362), .P23(n11361), 
            .P22(n11360), .P21(n11359), .P20(n11358), .P19(n11357), 
            .P18(n11356), .P17(n11355), .P16(n11354), .P15(n11353), 
            .P14(n11352), .P13(n11351), .P12(n11350), .P11(n11349), 
            .P10(n11348), .P9(n11347), .P8(n11346), .P7(n11345), .P6(n11344), 
            .P5(n11343), .P4(n11342), .P3(n11341), .P2(n11340), .P1(n11339), 
            .P0(n11338), .SIGNEDP(n11337));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam a2_reg_15__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam a2_reg_15__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam a2_reg_15__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam a2_reg_15__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam a2_reg_15__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam a2_reg_15__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam a2_reg_15__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam a2_reg_15__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam a2_reg_15__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam a2_reg_15__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam a2_reg_15__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam a2_reg_15__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam a2_reg_15__I_0_mult_2.GSR = "DISABLED";
    defparam a2_reg_15__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam a2_reg_15__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam a2_reg_15__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam a2_reg_15__I_0_mult_2.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i9 (.D(c_c_9), .CK(clk_c), .Q(c1_reg[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i9.GSR = "ENABLED";
    ALU54B lat_alu_14 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n11123), .SIGNEDIB(n11196), .SIGNEDCIN(n11269), .A35(n11122), 
           .A34(n11121), .A33(n11120), .A32(n11119), .A31(n11118), .A30(n11117), 
           .A29(n11116), .A28(n11115), .A27(n11114), .A26(n11113), .A25(n11112), 
           .A24(n11111), .A23(n11110), .A22(n11109), .A21(n11108), .A20(n11107), 
           .A19(n11106), .A18(n11105), .A17(n11104), .A16(n11103), .A15(n11102), 
           .A14(n11101), .A13(n11100), .A12(n11099), .A11(n11098), .A10(n11097), 
           .A9(n11096), .A8(n11095), .A7(n11094), .A6(n11093), .A5(n11092), 
           .A4(n11091), .A3(n11090), .A2(n11089), .A1(n11088), .A0(n11087), 
           .B35(n11195), .B34(n11194), .B33(n11193), .B32(n11192), .B31(n11191), 
           .B30(n11190), .B29(n11189), .B28(n11188), .B27(n11187), .B26(n11186), 
           .B25(n11185), .B24(n11184), .B23(n11183), .B22(n11182), .B21(n11181), 
           .B20(n11180), .B19(n11179), .B18(n11178), .B17(n11177), .B16(n11176), 
           .B15(n11175), .B14(n11174), .B13(n11173), .B12(n11172), .B11(n11171), 
           .B10(n11170), .B9(n11169), .B8(n11168), .B7(n11167), .B6(n11166), 
           .B5(n11165), .B4(n11164), .B3(n11163), .B2(n11162), .B1(n11161), 
           .B0(n11160), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n11159), .MA34(n11158), .MA33(n11157), .MA32(n11156), 
           .MA31(n11155), .MA30(n11154), .MA29(n11153), .MA28(n11152), 
           .MA27(n11151), .MA26(n11150), .MA25(n11149), .MA24(n11148), 
           .MA23(n11147), .MA22(n11146), .MA21(n11145), .MA20(n11144), 
           .MA19(n11143), .MA18(n11142), .MA17(n11141), .MA16(n11140), 
           .MA15(n11139), .MA14(n11138), .MA13(n11137), .MA12(n11136), 
           .MA11(n11135), .MA10(n11134), .MA9(n11133), .MA8(n11132), 
           .MA7(n11131), .MA6(n11130), .MA5(n11129), .MA4(n11128), .MA3(n11127), 
           .MA2(n11126), .MA1(n11125), .MA0(n11124), .MB35(n11232), 
           .MB34(n11231), .MB33(n11230), .MB32(n11229), .MB31(n11228), 
           .MB30(n11227), .MB29(n11226), .MB28(n11225), .MB27(n11224), 
           .MB26(n11223), .MB25(n11222), .MB24(n11221), .MB23(n11220), 
           .MB22(n11219), .MB21(n11218), .MB20(n11217), .MB19(n11216), 
           .MB18(n11215), .MB17(n11214), .MB16(n11213), .MB15(n11212), 
           .MB14(n11211), .MB13(n11210), .MB12(n11209), .MB11(n11208), 
           .MB10(n11207), .MB9(n11206), .MB8(n11205), .MB7(n11204), 
           .MB6(n11203), .MB5(n11202), .MB4(n11201), .MB3(n11200), .MB2(n11199), 
           .MB1(n11198), .MB0(n11197), .CIN53(n11268), .CIN52(n11267), 
           .CIN51(n11266), .CIN50(n11265), .CIN49(n11264), .CIN48(n11263), 
           .CIN47(n11262), .CIN46(n11261), .CIN45(n11260), .CIN44(n11259), 
           .CIN43(n11258), .CIN42(n11257), .CIN41(n11256), .CIN40(n11255), 
           .CIN39(n11254), .CIN38(n11253), .CIN37(n11252), .CIN36(n11251), 
           .CIN35(n11250), .CIN34(n11249), .CIN33(n11248), .CIN32(n11247), 
           .CIN31(n11246), .CIN30(n11245), .CIN29(n11244), .CIN28(n11243), 
           .CIN27(n11242), .CIN26(n11241), .CIN25(n11240), .CIN24(n11239), 
           .CIN23(n11238), .CIN22(n11237), .CIN21(n11236), .CIN20(n11235), 
           .CIN19(n11234), .CIN18(n11233), .CIN17(prod_c[17]), .CIN16(prod_c[16]), 
           .CIN15(prod_c[15]), .CIN14(n10926), .CIN13(n10927), .CIN12(n10928), 
           .CIN11(n10929), .CIN10(n10930), .CIN9(n10931), .CIN8(n10932), 
           .CIN7(n10933), .CIN6(n10934), .CIN5(n10935), .CIN4(n10936), 
           .CIN3(n10937), .CIN2(n10938), .CIN1(n10939), .CIN0(n10940), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R29(prod_c[47]), 
           .R28(prod_c[46]), .R27(prod_c[45]), .R26(prod_c[44]), .R25(prod_c[43]), 
           .R24(prod_c[42]), .R23(prod_c[41]), .R22(prod_c[40]), .R21(prod_c[39]), 
           .R20(prod_c[38]), .R19(prod_c[37]), .R18(prod_c[36]), .R17(prod_c[35]), 
           .R16(prod_c[34]), .R15(prod_c[33]), .R14(prod_c[32]), .R13(prod_c[31]), 
           .R12(prod_c[30]), .R11(prod_c[29]), .R10(prod_c[28]), .R9(prod_c[27]), 
           .R8(prod_c[26]), .R7(prod_c[25]), .R6(prod_c[24]), .R5(prod_c[23]), 
           .R4(prod_c[22]), .R3(prod_c[21]), .R2(prod_c[20]), .R1(prod_c[19]), 
           .R0(prod_c[18]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[44:57])
    defparam lat_alu_14.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_14.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_14.REG_FLAG_CLK = "NONE";
    defparam lat_alu_14.REG_FLAG_CE = "CE0";
    defparam lat_alu_14.REG_FLAG_RST = "RST0";
    defparam lat_alu_14.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASK01 = "0x00000000000000";
    defparam lat_alu_14.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_14.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_14.CLK0_DIV = "ENABLED";
    defparam lat_alu_14.CLK1_DIV = "ENABLED";
    defparam lat_alu_14.CLK2_DIV = "ENABLED";
    defparam lat_alu_14.CLK3_DIV = "ENABLED";
    defparam lat_alu_14.MCPAT = "0x00000000000000";
    defparam lat_alu_14.MASKPAT = "0x00000000000000";
    defparam lat_alu_14.RNDPAT = "0x00000000000000";
    defparam lat_alu_14.GSR = "DISABLED";
    defparam lat_alu_14.RESETMODE = "SYNC";
    defparam lat_alu_14.MULT9_MODE = "DISABLED";
    defparam lat_alu_14.LEGACY = "DISABLED";
    FD1S3AX c1_reg_i8 (.D(c_c_8), .CK(clk_c), .Q(c1_reg[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i8.GSR = "ENABLED";
    ALU54B lat_alu_13 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10977), .SIGNEDIB(n11050), .SIGNEDCIN(GND_net), 
           .A35(n10976), .A34(n10975), .A33(n10974), .A32(n10973), .A31(n10972), 
           .A30(n10971), .A29(n10970), .A28(n10969), .A27(n10968), .A26(n10967), 
           .A25(n10966), .A24(n10965), .A23(n10964), .A22(n10963), .A21(n10962), 
           .A20(n10961), .A19(n10960), .A18(n10959), .A17(n10958), .A16(n10957), 
           .A15(n10956), .A14(n10955), .A13(n10954), .A12(n10953), .A11(n10952), 
           .A10(n10951), .A9(n10950), .A8(n10949), .A7(n10948), .A6(n10947), 
           .A5(n10946), .A4(n10945), .A3(n10944), .A2(n10943), .A1(n10942), 
           .A0(n10941), .B35(n11049), .B34(n11048), .B33(n11047), .B32(n11046), 
           .B31(n11045), .B30(n11044), .B29(n11043), .B28(n11042), .B27(n11041), 
           .B26(n11040), .B25(n11039), .B24(n11038), .B23(n11037), .B22(n11036), 
           .B21(n11035), .B20(n11034), .B19(n11033), .B18(n11032), .B17(n11031), 
           .B16(n11030), .B15(n11029), .B14(n11028), .B13(n11027), .B12(n11026), 
           .B11(n11025), .B10(n11024), .B9(n11023), .B8(n11022), .B7(n11021), 
           .B6(n11020), .B5(n11019), .B4(n11018), .B3(n11017), .B2(n11016), 
           .B1(n11015), .B0(n11014), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n11013), .MA34(n11012), .MA33(n11011), .MA32(n11010), 
           .MA31(n11009), .MA30(n11008), .MA29(n11007), .MA28(n11006), 
           .MA27(n11005), .MA26(n11004), .MA25(n11003), .MA24(n11002), 
           .MA23(n11001), .MA22(n11000), .MA21(n10999), .MA20(n10998), 
           .MA19(n10997), .MA18(n10996), .MA17(n10995), .MA16(n10994), 
           .MA15(n10993), .MA14(n10992), .MA13(n10991), .MA12(n10990), 
           .MA11(n10989), .MA10(n10988), .MA9(n10987), .MA8(n10986), 
           .MA7(n10985), .MA6(n10984), .MA5(n10983), .MA4(n10982), .MA3(n10981), 
           .MA2(n10980), .MA1(n10979), .MA0(n10978), .MB35(n11086), 
           .MB34(n11085), .MB33(n11084), .MB32(n11083), .MB31(n11082), 
           .MB30(n11081), .MB29(n11080), .MB28(n11079), .MB27(n11078), 
           .MB26(n11077), .MB25(n11076), .MB24(n11075), .MB23(n11074), 
           .MB22(n11073), .MB21(n11072), .MB20(n11071), .MB19(n11070), 
           .MB18(n11069), .MB17(n11068), .MB16(n11067), .MB15(n11066), 
           .MB14(n11065), .MB13(n11064), .MB12(n11063), .MB11(n11062), 
           .MB10(n11061), .MB9(n11060), .MB8(n11059), .MB7(n11058), 
           .MB6(n11057), .MB5(n11056), .MB4(n11055), .MB3(n11054), .MB2(n11053), 
           .MB1(n11052), .MB0(n11051), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n11268), 
           .R52(n11267), .R51(n11266), .R50(n11265), .R49(n11264), .R48(n11263), 
           .R47(n11262), .R46(n11261), .R45(n11260), .R44(n11259), .R43(n11258), 
           .R42(n11257), .R41(n11256), .R40(n11255), .R39(n11254), .R38(n11253), 
           .R37(n11252), .R36(n11251), .R35(n11250), .R34(n11249), .R33(n11248), 
           .R32(n11247), .R31(n11246), .R30(n11245), .R29(n11244), .R28(n11243), 
           .R27(n11242), .R26(n11241), .R25(n11240), .R24(n11239), .R23(n11238), 
           .R22(n11237), .R21(n11236), .R20(n11235), .R19(n11234), .R18(n11233), 
           .R17(prod_c[17]), .R16(prod_c[16]), .R15(prod_c[15]), .R14(n10926), 
           .R13(n10927), .R12(n10928), .R11(n10929), .R10(n10930), .R9(n10931), 
           .R8(n10932), .R7(n10933), .R6(n10934), .R5(n10935), .R4(n10936), 
           .R3(n10937), .R2(n10938), .R1(n10939), .R0(n10940), .SIGNEDR(n11269));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[44:57])
    defparam lat_alu_13.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_13.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_13.REG_FLAG_CLK = "NONE";
    defparam lat_alu_13.REG_FLAG_CE = "CE0";
    defparam lat_alu_13.REG_FLAG_RST = "RST0";
    defparam lat_alu_13.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASK01 = "0x00000000000000";
    defparam lat_alu_13.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_13.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_13.CLK0_DIV = "ENABLED";
    defparam lat_alu_13.CLK1_DIV = "ENABLED";
    defparam lat_alu_13.CLK2_DIV = "ENABLED";
    defparam lat_alu_13.CLK3_DIV = "ENABLED";
    defparam lat_alu_13.MCPAT = "0x00000000000000";
    defparam lat_alu_13.MASKPAT = "0x00000000000000";
    defparam lat_alu_13.RNDPAT = "0x00000000000000";
    defparam lat_alu_13.GSR = "DISABLED";
    defparam lat_alu_13.RESETMODE = "SYNC";
    defparam lat_alu_13.MULT9_MODE = "DISABLED";
    defparam lat_alu_13.LEGACY = "DISABLED";
    FD1S3AX c1_reg_i7 (.D(c_c_7), .CK(clk_c), .Q(c1_reg[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i7.GSR = "ENABLED";
    MULT18X18D lat_mult_12 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[16]), .B14(c_s[16]), .B13(c_s[16]), .B12(c_s[16]), 
            .B11(c_s[16]), .B10(c_s[16]), .B9(c_s[16]), .B8(c_s[16]), 
            .B7(c_s[16]), .B6(c_s[16]), .B5(c_s[16]), .B4(c_s[16]), 
            .B3(c_s[16]), .B2(c_s[16]), .B1(c_s[16]), .B0(c_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n11177), .ROA16(n11176), 
            .ROA15(n11175), .ROA14(n11174), .ROA13(n11173), .ROA12(n11172), 
            .ROA11(n11171), .ROA10(n11170), .ROA9(n11169), .ROA8(n11168), 
            .ROA7(n11167), .ROA6(n11166), .ROA5(n11165), .ROA4(n11164), 
            .ROA3(n11163), .ROA2(n11162), .ROA1(n11161), .ROA0(n11160), 
            .ROB17(n11195), .ROB16(n11194), .ROB15(n11193), .ROB14(n11192), 
            .ROB13(n11191), .ROB12(n11190), .ROB11(n11189), .ROB10(n11188), 
            .ROB9(n11187), .ROB8(n11186), .ROB7(n11185), .ROB6(n11184), 
            .ROB5(n11183), .ROB4(n11182), .ROB3(n11181), .ROB2(n11180), 
            .ROB1(n11179), .ROB0(n11178), .P35(n11232), .P34(n11231), 
            .P33(n11230), .P32(n11229), .P31(n11228), .P30(n11227), 
            .P29(n11226), .P28(n11225), .P27(n11224), .P26(n11223), 
            .P25(n11222), .P24(n11221), .P23(n11220), .P22(n11219), 
            .P21(n11218), .P20(n11217), .P19(n11216), .P18(n11215), 
            .P17(n11214), .P16(n11213), .P15(n11212), .P14(n11211), 
            .P13(n11210), .P12(n11209), .P11(n11208), .P10(n11207), 
            .P9(n11206), .P8(n11205), .P7(n11204), .P6(n11203), .P5(n11202), 
            .P4(n11201), .P3(n11200), .P2(n11199), .P1(n11198), .P0(n11197), 
            .SIGNEDP(n11196));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[44:57])
    defparam lat_mult_12.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_12.REG_INPUTA_CE = "CE3";
    defparam lat_mult_12.REG_INPUTA_RST = "RST3";
    defparam lat_mult_12.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTB_CE = "CE0";
    defparam lat_mult_12.REG_INPUTB_RST = "RST0";
    defparam lat_mult_12.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTC_CE = "CE0";
    defparam lat_mult_12.REG_INPUTC_RST = "RST0";
    defparam lat_mult_12.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_12.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_12.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_12.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_12.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_12.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_12.CLK0_DIV = "ENABLED";
    defparam lat_mult_12.CLK1_DIV = "ENABLED";
    defparam lat_mult_12.CLK2_DIV = "ENABLED";
    defparam lat_mult_12.CLK3_DIV = "ENABLED";
    defparam lat_mult_12.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_12.GSR = "DISABLED";
    defparam lat_mult_12.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_12.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_12.MULT_BYPASS = "DISABLED";
    defparam lat_mult_12.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i6 (.D(c_c_6), .CK(clk_c), .Q(c1_reg[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i6.GSR = "ENABLED";
    MULT18X18D lat_mult_11 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[16]), .B14(c_s[16]), .B13(c_s[16]), .B12(c_s[16]), 
            .B11(c_s[16]), .B10(c_s[16]), .B9(c_s[16]), .B8(c_s[16]), 
            .B7(c_s[16]), .B6(c_s[16]), .B5(c_s[16]), .B4(c_s[16]), 
            .B3(c_s[16]), .B2(c_s[16]), .B1(c_s[16]), .B0(c_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n11104), .ROA16(n11103), 
            .ROA15(n11102), .ROA14(n11101), .ROA13(n11100), .ROA12(n11099), 
            .ROA11(n11098), .ROA10(n11097), .ROA9(n11096), .ROA8(n11095), 
            .ROA7(n11094), .ROA6(n11093), .ROA5(n11092), .ROA4(n11091), 
            .ROA3(n11090), .ROA2(n11089), .ROA1(n11088), .ROA0(n11087), 
            .ROB17(n11122), .ROB16(n11121), .ROB15(n11120), .ROB14(n11119), 
            .ROB13(n11118), .ROB12(n11117), .ROB11(n11116), .ROB10(n11115), 
            .ROB9(n11114), .ROB8(n11113), .ROB7(n11112), .ROB6(n11111), 
            .ROB5(n11110), .ROB4(n11109), .ROB3(n11108), .ROB2(n11107), 
            .ROB1(n11106), .ROB0(n11105), .P35(n11159), .P34(n11158), 
            .P33(n11157), .P32(n11156), .P31(n11155), .P30(n11154), 
            .P29(n11153), .P28(n11152), .P27(n11151), .P26(n11150), 
            .P25(n11149), .P24(n11148), .P23(n11147), .P22(n11146), 
            .P21(n11145), .P20(n11144), .P19(n11143), .P18(n11142), 
            .P17(n11141), .P16(n11140), .P15(n11139), .P14(n11138), 
            .P13(n11137), .P12(n11136), .P11(n11135), .P10(n11134), 
            .P9(n11133), .P8(n11132), .P7(n11131), .P6(n11130), .P5(n11129), 
            .P4(n11128), .P3(n11127), .P2(n11126), .P1(n11125), .P0(n11124), 
            .SIGNEDP(n11123));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[44:57])
    defparam lat_mult_11.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_11.REG_INPUTA_CE = "CE3";
    defparam lat_mult_11.REG_INPUTA_RST = "RST3";
    defparam lat_mult_11.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTB_CE = "CE0";
    defparam lat_mult_11.REG_INPUTB_RST = "RST0";
    defparam lat_mult_11.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTC_CE = "CE0";
    defparam lat_mult_11.REG_INPUTC_RST = "RST0";
    defparam lat_mult_11.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_11.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_11.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_11.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_11.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_11.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_11.CLK0_DIV = "ENABLED";
    defparam lat_mult_11.CLK1_DIV = "ENABLED";
    defparam lat_mult_11.CLK2_DIV = "ENABLED";
    defparam lat_mult_11.CLK3_DIV = "ENABLED";
    defparam lat_mult_11.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_11.GSR = "DISABLED";
    defparam lat_mult_11.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_11.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_11.MULT_BYPASS = "DISABLED";
    defparam lat_mult_11.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i5 (.D(c_c_5), .CK(clk_c), .Q(c1_reg[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i5.GSR = "ENABLED";
    MULT18X18D lat_mult_10 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[15]), .B14(c_s[14]), .B13(c_s[13]), .B12(c_s[12]), 
            .B11(c_s[11]), .B10(c_s[10]), .B9(c_s[9]), .B8(c_s[8]), 
            .B7(c_s[7]), .B6(c_s[6]), .B5(c_s[5]), .B4(c_s[4]), .B3(c_s[3]), 
            .B2(c_s[2]), .B1(c_s[1]), .B0(c_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n11031), .ROA16(n11030), .ROA15(n11029), .ROA14(n11028), 
            .ROA13(n11027), .ROA12(n11026), .ROA11(n11025), .ROA10(n11024), 
            .ROA9(n11023), .ROA8(n11022), .ROA7(n11021), .ROA6(n11020), 
            .ROA5(n11019), .ROA4(n11018), .ROA3(n11017), .ROA2(n11016), 
            .ROA1(n11015), .ROA0(n11014), .ROB17(n11049), .ROB16(n11048), 
            .ROB15(n11047), .ROB14(n11046), .ROB13(n11045), .ROB12(n11044), 
            .ROB11(n11043), .ROB10(n11042), .ROB9(n11041), .ROB8(n11040), 
            .ROB7(n11039), .ROB6(n11038), .ROB5(n11037), .ROB4(n11036), 
            .ROB3(n11035), .ROB2(n11034), .ROB1(n11033), .ROB0(n11032), 
            .P35(n11086), .P34(n11085), .P33(n11084), .P32(n11083), 
            .P31(n11082), .P30(n11081), .P29(n11080), .P28(n11079), 
            .P27(n11078), .P26(n11077), .P25(n11076), .P24(n11075), 
            .P23(n11074), .P22(n11073), .P21(n11072), .P20(n11071), 
            .P19(n11070), .P18(n11069), .P17(n11068), .P16(n11067), 
            .P15(n11066), .P14(n11065), .P13(n11064), .P12(n11063), 
            .P11(n11062), .P10(n11061), .P9(n11060), .P8(n11059), .P7(n11058), 
            .P6(n11057), .P5(n11056), .P4(n11055), .P3(n11054), .P2(n11053), 
            .P1(n11052), .P0(n11051), .SIGNEDP(n11050));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[44:57])
    defparam lat_mult_10.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_10.REG_INPUTA_CE = "CE3";
    defparam lat_mult_10.REG_INPUTA_RST = "RST3";
    defparam lat_mult_10.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTB_CE = "CE0";
    defparam lat_mult_10.REG_INPUTB_RST = "RST0";
    defparam lat_mult_10.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTC_CE = "CE0";
    defparam lat_mult_10.REG_INPUTC_RST = "RST0";
    defparam lat_mult_10.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_10.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_10.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_10.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_10.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_10.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_10.CLK0_DIV = "ENABLED";
    defparam lat_mult_10.CLK1_DIV = "ENABLED";
    defparam lat_mult_10.CLK2_DIV = "ENABLED";
    defparam lat_mult_10.CLK3_DIV = "ENABLED";
    defparam lat_mult_10.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_10.GSR = "DISABLED";
    defparam lat_mult_10.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_10.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_10.MULT_BYPASS = "DISABLED";
    defparam lat_mult_10.RESETMODE = "ASYNC";
    MULT18X18D c_s_31__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[15]), .B14(c_s[14]), .B13(c_s[13]), .B12(c_s[12]), 
            .B11(c_s[11]), .B10(c_s[10]), .B9(c_s[9]), .B8(c_s[8]), 
            .B7(c_s[7]), .B6(c_s[6]), .B5(c_s[5]), .B4(c_s[4]), .B3(c_s[3]), 
            .B2(c_s[2]), .B1(c_s[1]), .B0(c_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10958), .ROA16(n10957), .ROA15(n10956), .ROA14(n10955), 
            .ROA13(n10954), .ROA12(n10953), .ROA11(n10952), .ROA10(n10951), 
            .ROA9(n10950), .ROA8(n10949), .ROA7(n10948), .ROA6(n10947), 
            .ROA5(n10946), .ROA4(n10945), .ROA3(n10944), .ROA2(n10943), 
            .ROA1(n10942), .ROA0(n10941), .ROB17(n10976), .ROB16(n10975), 
            .ROB15(n10974), .ROB14(n10973), .ROB13(n10972), .ROB12(n10971), 
            .ROB11(n10970), .ROB10(n10969), .ROB9(n10968), .ROB8(n10967), 
            .ROB7(n10966), .ROB6(n10965), .ROB5(n10964), .ROB4(n10963), 
            .ROB3(n10962), .ROB2(n10961), .ROB1(n10960), .ROB0(n10959), 
            .P35(n11013), .P34(n11012), .P33(n11011), .P32(n11010), 
            .P31(n11009), .P30(n11008), .P29(n11007), .P28(n11006), 
            .P27(n11005), .P26(n11004), .P25(n11003), .P24(n11002), 
            .P23(n11001), .P22(n11000), .P21(n10999), .P20(n10998), 
            .P19(n10997), .P18(n10996), .P17(n10995), .P16(n10994), 
            .P15(n10993), .P14(n10992), .P13(n10991), .P12(n10990), 
            .P11(n10989), .P10(n10988), .P9(n10987), .P8(n10986), .P7(n10985), 
            .P6(n10984), .P5(n10983), .P4(n10982), .P3(n10981), .P2(n10980), 
            .P1(n10979), .P0(n10978), .SIGNEDP(n10977));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(103[44:57])
    defparam c_s_31__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam c_s_31__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam c_s_31__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam c_s_31__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam c_s_31__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam c_s_31__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam c_s_31__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam c_s_31__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.GSR = "DISABLED";
    defparam c_s_31__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam c_s_31__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam c_s_31__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam c_s_31__I_0_mult_2.RESETMODE = "ASYNC";
    FD1S3AX c1_reg_i4 (.D(c_c_4), .CK(clk_c), .Q(c1_reg[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i4.GSR = "ENABLED";
    ALU54B lat_alu_9 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10763), .SIGNEDIB(n10836), .SIGNEDCIN(n10909), .A35(n10762), 
           .A34(n10761), .A33(n10760), .A32(n10759), .A31(n10758), .A30(n10757), 
           .A29(n10756), .A28(n10755), .A27(n10754), .A26(n10753), .A25(n10752), 
           .A24(n10751), .A23(n10750), .A22(n10749), .A21(n10748), .A20(n10747), 
           .A19(n10746), .A18(n10745), .A17(n10744), .A16(n10743), .A15(n10742), 
           .A14(n10741), .A13(n10740), .A12(n10739), .A11(n10738), .A10(n10737), 
           .A9(n10736), .A8(n10735), .A7(n10734), .A6(n10733), .A5(n10732), 
           .A4(n10731), .A3(n10730), .A2(n10729), .A1(n10728), .A0(n10727), 
           .B35(n10835), .B34(n10834), .B33(n10833), .B32(n10832), .B31(n10831), 
           .B30(n10830), .B29(n10829), .B28(n10828), .B27(n10827), .B26(n10826), 
           .B25(n10825), .B24(n10824), .B23(n10823), .B22(n10822), .B21(n10821), 
           .B20(n10820), .B19(n10819), .B18(n10818), .B17(n10817), .B16(n10816), 
           .B15(n10815), .B14(n10814), .B13(n10813), .B12(n10812), .B11(n10811), 
           .B10(n10810), .B9(n10809), .B8(n10808), .B7(n10807), .B6(n10806), 
           .B5(n10805), .B4(n10804), .B3(n10803), .B2(n10802), .B1(n10801), 
           .B0(n10800), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10799), .MA34(n10798), .MA33(n10797), .MA32(n10796), 
           .MA31(n10795), .MA30(n10794), .MA29(n10793), .MA28(n10792), 
           .MA27(n10791), .MA26(n10790), .MA25(n10789), .MA24(n10788), 
           .MA23(n10787), .MA22(n10786), .MA21(n10785), .MA20(n10784), 
           .MA19(n10783), .MA18(n10782), .MA17(n10781), .MA16(n10780), 
           .MA15(n10779), .MA14(n10778), .MA13(n10777), .MA12(n10776), 
           .MA11(n10775), .MA10(n10774), .MA9(n10773), .MA8(n10772), 
           .MA7(n10771), .MA6(n10770), .MA5(n10769), .MA4(n10768), .MA3(n10767), 
           .MA2(n10766), .MA1(n10765), .MA0(n10764), .MB35(n10872), 
           .MB34(n10871), .MB33(n10870), .MB32(n10869), .MB31(n10868), 
           .MB30(n10867), .MB29(n10866), .MB28(n10865), .MB27(n10864), 
           .MB26(n10863), .MB25(n10862), .MB24(n10861), .MB23(n10860), 
           .MB22(n10859), .MB21(n10858), .MB20(n10857), .MB19(n10856), 
           .MB18(n10855), .MB17(n10854), .MB16(n10853), .MB15(n10852), 
           .MB14(n10851), .MB13(n10850), .MB12(n10849), .MB11(n10848), 
           .MB10(n10847), .MB9(n10846), .MB8(n10845), .MB7(n10844), 
           .MB6(n10843), .MB5(n10842), .MB4(n10841), .MB3(n10840), .MB2(n10839), 
           .MB1(n10838), .MB0(n10837), .CIN53(n10908), .CIN52(n10907), 
           .CIN51(n10906), .CIN50(n10905), .CIN49(n10904), .CIN48(n10903), 
           .CIN47(n10902), .CIN46(n10901), .CIN45(n10900), .CIN44(n10899), 
           .CIN43(n10898), .CIN42(n10897), .CIN41(n10896), .CIN40(n10895), 
           .CIN39(n10894), .CIN38(n10893), .CIN37(n10892), .CIN36(n10891), 
           .CIN35(n10890), .CIN34(n10889), .CIN33(n10888), .CIN32(n10887), 
           .CIN31(n10886), .CIN30(n10885), .CIN29(n10884), .CIN28(n10883), 
           .CIN27(n10882), .CIN26(n10881), .CIN25(n10880), .CIN24(n10879), 
           .CIN23(n10878), .CIN22(n10877), .CIN21(n10876), .CIN20(n10875), 
           .CIN19(n10874), .CIN18(n10873), .CIN17(prod_b[17]), .CIN16(prod_b[16]), 
           .CIN15(prod_b[15]), .CIN14(n10566), .CIN13(n10567), .CIN12(n10568), 
           .CIN11(n10569), .CIN10(n10570), .CIN9(n10571), .CIN8(n10572), 
           .CIN7(n10573), .CIN6(n10574), .CIN5(n10575), .CIN4(n10576), 
           .CIN3(n10577), .CIN2(n10578), .CIN1(n10579), .CIN0(n10580), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R29(prod_b[47]), 
           .R28(prod_b[46]), .R27(prod_b[45]), .R26(prod_b[44]), .R25(prod_b[43]), 
           .R24(prod_b[42]), .R23(prod_b[41]), .R22(prod_b[40]), .R21(prod_b[39]), 
           .R20(prod_b[38]), .R19(prod_b[37]), .R18(prod_b[36]), .R17(prod_b[35]), 
           .R16(prod_b[34]), .R15(prod_b[33]), .R14(prod_b[32]), .R13(prod_b[31]), 
           .R12(prod_b[30]), .R11(prod_b[29]), .R10(prod_b[28]), .R9(prod_b[27]), 
           .R8(prod_b[26]), .R7(prod_b[25]), .R6(prod_b[24]), .R5(prod_b[23]), 
           .R4(prod_b[22]), .R3(prod_b[21]), .R2(prod_b[20]), .R1(prod_b[19]), 
           .R0(prod_b[18]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[44:57])
    defparam lat_alu_9.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_9.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_9.REG_FLAG_CLK = "NONE";
    defparam lat_alu_9.REG_FLAG_CE = "CE0";
    defparam lat_alu_9.REG_FLAG_RST = "RST0";
    defparam lat_alu_9.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASK01 = "0x00000000000000";
    defparam lat_alu_9.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_9.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_9.CLK0_DIV = "ENABLED";
    defparam lat_alu_9.CLK1_DIV = "ENABLED";
    defparam lat_alu_9.CLK2_DIV = "ENABLED";
    defparam lat_alu_9.CLK3_DIV = "ENABLED";
    defparam lat_alu_9.MCPAT = "0x00000000000000";
    defparam lat_alu_9.MASKPAT = "0x00000000000000";
    defparam lat_alu_9.RNDPAT = "0x00000000000000";
    defparam lat_alu_9.GSR = "DISABLED";
    defparam lat_alu_9.RESETMODE = "SYNC";
    defparam lat_alu_9.MULT9_MODE = "DISABLED";
    defparam lat_alu_9.LEGACY = "DISABLED";
    ALU54B lat_alu_8 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10617), .SIGNEDIB(n10690), .SIGNEDCIN(GND_net), 
           .A35(n10616), .A34(n10615), .A33(n10614), .A32(n10613), .A31(n10612), 
           .A30(n10611), .A29(n10610), .A28(n10609), .A27(n10608), .A26(n10607), 
           .A25(n10606), .A24(n10605), .A23(n10604), .A22(n10603), .A21(n10602), 
           .A20(n10601), .A19(n10600), .A18(n10599), .A17(n10598), .A16(n10597), 
           .A15(n10596), .A14(n10595), .A13(n10594), .A12(n10593), .A11(n10592), 
           .A10(n10591), .A9(n10590), .A8(n10589), .A7(n10588), .A6(n10587), 
           .A5(n10586), .A4(n10585), .A3(n10584), .A2(n10583), .A1(n10582), 
           .A0(n10581), .B35(n10689), .B34(n10688), .B33(n10687), .B32(n10686), 
           .B31(n10685), .B30(n10684), .B29(n10683), .B28(n10682), .B27(n10681), 
           .B26(n10680), .B25(n10679), .B24(n10678), .B23(n10677), .B22(n10676), 
           .B21(n10675), .B20(n10674), .B19(n10673), .B18(n10672), .B17(n10671), 
           .B16(n10670), .B15(n10669), .B14(n10668), .B13(n10667), .B12(n10666), 
           .B11(n10665), .B10(n10664), .B9(n10663), .B8(n10662), .B7(n10661), 
           .B6(n10660), .B5(n10659), .B4(n10658), .B3(n10657), .B2(n10656), 
           .B1(n10655), .B0(n10654), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10653), .MA34(n10652), .MA33(n10651), .MA32(n10650), 
           .MA31(n10649), .MA30(n10648), .MA29(n10647), .MA28(n10646), 
           .MA27(n10645), .MA26(n10644), .MA25(n10643), .MA24(n10642), 
           .MA23(n10641), .MA22(n10640), .MA21(n10639), .MA20(n10638), 
           .MA19(n10637), .MA18(n10636), .MA17(n10635), .MA16(n10634), 
           .MA15(n10633), .MA14(n10632), .MA13(n10631), .MA12(n10630), 
           .MA11(n10629), .MA10(n10628), .MA9(n10627), .MA8(n10626), 
           .MA7(n10625), .MA6(n10624), .MA5(n10623), .MA4(n10622), .MA3(n10621), 
           .MA2(n10620), .MA1(n10619), .MA0(n10618), .MB35(n10726), 
           .MB34(n10725), .MB33(n10724), .MB32(n10723), .MB31(n10722), 
           .MB30(n10721), .MB29(n10720), .MB28(n10719), .MB27(n10718), 
           .MB26(n10717), .MB25(n10716), .MB24(n10715), .MB23(n10714), 
           .MB22(n10713), .MB21(n10712), .MB20(n10711), .MB19(n10710), 
           .MB18(n10709), .MB17(n10708), .MB16(n10707), .MB15(n10706), 
           .MB14(n10705), .MB13(n10704), .MB12(n10703), .MB11(n10702), 
           .MB10(n10701), .MB9(n10700), .MB8(n10699), .MB7(n10698), 
           .MB6(n10697), .MB5(n10696), .MB4(n10695), .MB3(n10694), .MB2(n10693), 
           .MB1(n10692), .MB0(n10691), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n10908), 
           .R52(n10907), .R51(n10906), .R50(n10905), .R49(n10904), .R48(n10903), 
           .R47(n10902), .R46(n10901), .R45(n10900), .R44(n10899), .R43(n10898), 
           .R42(n10897), .R41(n10896), .R40(n10895), .R39(n10894), .R38(n10893), 
           .R37(n10892), .R36(n10891), .R35(n10890), .R34(n10889), .R33(n10888), 
           .R32(n10887), .R31(n10886), .R30(n10885), .R29(n10884), .R28(n10883), 
           .R27(n10882), .R26(n10881), .R25(n10880), .R24(n10879), .R23(n10878), 
           .R22(n10877), .R21(n10876), .R20(n10875), .R19(n10874), .R18(n10873), 
           .R17(prod_b[17]), .R16(prod_b[16]), .R15(prod_b[15]), .R14(n10566), 
           .R13(n10567), .R12(n10568), .R11(n10569), .R10(n10570), .R9(n10571), 
           .R8(n10572), .R7(n10573), .R6(n10574), .R5(n10575), .R4(n10576), 
           .R3(n10577), .R2(n10578), .R1(n10579), .R0(n10580), .SIGNEDR(n10909));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[44:57])
    defparam lat_alu_8.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_8.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_8.REG_FLAG_CLK = "NONE";
    defparam lat_alu_8.REG_FLAG_CE = "CE0";
    defparam lat_alu_8.REG_FLAG_RST = "RST0";
    defparam lat_alu_8.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASK01 = "0x00000000000000";
    defparam lat_alu_8.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_8.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_8.CLK0_DIV = "ENABLED";
    defparam lat_alu_8.CLK1_DIV = "ENABLED";
    defparam lat_alu_8.CLK2_DIV = "ENABLED";
    defparam lat_alu_8.CLK3_DIV = "ENABLED";
    defparam lat_alu_8.MCPAT = "0x00000000000000";
    defparam lat_alu_8.MASKPAT = "0x00000000000000";
    defparam lat_alu_8.RNDPAT = "0x00000000000000";
    defparam lat_alu_8.GSR = "DISABLED";
    defparam lat_alu_8.RESETMODE = "SYNC";
    defparam lat_alu_8.MULT9_MODE = "DISABLED";
    defparam lat_alu_8.LEGACY = "DISABLED";
    MULT18X18D lat_mult_7 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[16]), .B14(b_s[16]), .B13(b_s[16]), .B12(b_s[16]), 
            .B11(b_s[16]), .B10(b_s[16]), .B9(b_s[16]), .B8(b_s[16]), 
            .B7(b_s[16]), .B6(b_s[16]), .B5(b_s[16]), .B4(b_s[16]), 
            .B3(b_s[16]), .B2(b_s[16]), .B1(b_s[16]), .B0(b_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10817), .ROA16(n10816), 
            .ROA15(n10815), .ROA14(n10814), .ROA13(n10813), .ROA12(n10812), 
            .ROA11(n10811), .ROA10(n10810), .ROA9(n10809), .ROA8(n10808), 
            .ROA7(n10807), .ROA6(n10806), .ROA5(n10805), .ROA4(n10804), 
            .ROA3(n10803), .ROA2(n10802), .ROA1(n10801), .ROA0(n10800), 
            .ROB17(n10835), .ROB16(n10834), .ROB15(n10833), .ROB14(n10832), 
            .ROB13(n10831), .ROB12(n10830), .ROB11(n10829), .ROB10(n10828), 
            .ROB9(n10827), .ROB8(n10826), .ROB7(n10825), .ROB6(n10824), 
            .ROB5(n10823), .ROB4(n10822), .ROB3(n10821), .ROB2(n10820), 
            .ROB1(n10819), .ROB0(n10818), .P35(n10872), .P34(n10871), 
            .P33(n10870), .P32(n10869), .P31(n10868), .P30(n10867), 
            .P29(n10866), .P28(n10865), .P27(n10864), .P26(n10863), 
            .P25(n10862), .P24(n10861), .P23(n10860), .P22(n10859), 
            .P21(n10858), .P20(n10857), .P19(n10856), .P18(n10855), 
            .P17(n10854), .P16(n10853), .P15(n10852), .P14(n10851), 
            .P13(n10850), .P12(n10849), .P11(n10848), .P10(n10847), 
            .P9(n10846), .P8(n10845), .P7(n10844), .P6(n10843), .P5(n10842), 
            .P4(n10841), .P3(n10840), .P2(n10839), .P1(n10838), .P0(n10837), 
            .SIGNEDP(n10836));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[44:57])
    defparam lat_mult_7.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_7.REG_INPUTA_CE = "CE3";
    defparam lat_mult_7.REG_INPUTA_RST = "RST3";
    defparam lat_mult_7.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTB_CE = "CE0";
    defparam lat_mult_7.REG_INPUTB_RST = "RST0";
    defparam lat_mult_7.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTC_CE = "CE0";
    defparam lat_mult_7.REG_INPUTC_RST = "RST0";
    defparam lat_mult_7.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_7.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_7.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_7.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_7.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_7.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_7.CLK0_DIV = "ENABLED";
    defparam lat_mult_7.CLK1_DIV = "ENABLED";
    defparam lat_mult_7.CLK2_DIV = "ENABLED";
    defparam lat_mult_7.CLK3_DIV = "ENABLED";
    defparam lat_mult_7.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_7.GSR = "DISABLED";
    defparam lat_mult_7.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_7.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_7.MULT_BYPASS = "DISABLED";
    defparam lat_mult_7.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_6 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[16]), .B14(b_s[16]), .B13(b_s[16]), .B12(b_s[16]), 
            .B11(b_s[16]), .B10(b_s[16]), .B9(b_s[16]), .B8(b_s[16]), 
            .B7(b_s[16]), .B6(b_s[16]), .B5(b_s[16]), .B4(b_s[16]), 
            .B3(b_s[16]), .B2(b_s[16]), .B1(b_s[16]), .B0(b_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10744), .ROA16(n10743), 
            .ROA15(n10742), .ROA14(n10741), .ROA13(n10740), .ROA12(n10739), 
            .ROA11(n10738), .ROA10(n10737), .ROA9(n10736), .ROA8(n10735), 
            .ROA7(n10734), .ROA6(n10733), .ROA5(n10732), .ROA4(n10731), 
            .ROA3(n10730), .ROA2(n10729), .ROA1(n10728), .ROA0(n10727), 
            .ROB17(n10762), .ROB16(n10761), .ROB15(n10760), .ROB14(n10759), 
            .ROB13(n10758), .ROB12(n10757), .ROB11(n10756), .ROB10(n10755), 
            .ROB9(n10754), .ROB8(n10753), .ROB7(n10752), .ROB6(n10751), 
            .ROB5(n10750), .ROB4(n10749), .ROB3(n10748), .ROB2(n10747), 
            .ROB1(n10746), .ROB0(n10745), .P35(n10799), .P34(n10798), 
            .P33(n10797), .P32(n10796), .P31(n10795), .P30(n10794), 
            .P29(n10793), .P28(n10792), .P27(n10791), .P26(n10790), 
            .P25(n10789), .P24(n10788), .P23(n10787), .P22(n10786), 
            .P21(n10785), .P20(n10784), .P19(n10783), .P18(n10782), 
            .P17(n10781), .P16(n10780), .P15(n10779), .P14(n10778), 
            .P13(n10777), .P12(n10776), .P11(n10775), .P10(n10774), 
            .P9(n10773), .P8(n10772), .P7(n10771), .P6(n10770), .P5(n10769), 
            .P4(n10768), .P3(n10767), .P2(n10766), .P1(n10765), .P0(n10764), 
            .SIGNEDP(n10763));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[44:57])
    defparam lat_mult_6.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_6.REG_INPUTA_CE = "CE3";
    defparam lat_mult_6.REG_INPUTA_RST = "RST3";
    defparam lat_mult_6.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTB_CE = "CE0";
    defparam lat_mult_6.REG_INPUTB_RST = "RST0";
    defparam lat_mult_6.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTC_CE = "CE0";
    defparam lat_mult_6.REG_INPUTC_RST = "RST0";
    defparam lat_mult_6.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_6.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_6.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_6.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_6.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_6.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_6.CLK0_DIV = "ENABLED";
    defparam lat_mult_6.CLK1_DIV = "ENABLED";
    defparam lat_mult_6.CLK2_DIV = "ENABLED";
    defparam lat_mult_6.CLK3_DIV = "ENABLED";
    defparam lat_mult_6.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_6.GSR = "DISABLED";
    defparam lat_mult_6.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_6.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_6.MULT_BYPASS = "DISABLED";
    defparam lat_mult_6.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_5 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[15]), .B14(b_s[14]), .B13(b_s[13]), .B12(b_s[12]), 
            .B11(b_s[11]), .B10(b_s[10]), .B9(b_s[9]), .B8(b_s[8]), 
            .B7(b_s[7]), .B6(b_s[6]), .B5(b_s[5]), .B4(b_s[4]), .B3(b_s[3]), 
            .B2(b_s[2]), .B1(b_s[1]), .B0(b_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10671), .ROA16(n10670), .ROA15(n10669), .ROA14(n10668), 
            .ROA13(n10667), .ROA12(n10666), .ROA11(n10665), .ROA10(n10664), 
            .ROA9(n10663), .ROA8(n10662), .ROA7(n10661), .ROA6(n10660), 
            .ROA5(n10659), .ROA4(n10658), .ROA3(n10657), .ROA2(n10656), 
            .ROA1(n10655), .ROA0(n10654), .ROB17(n10689), .ROB16(n10688), 
            .ROB15(n10687), .ROB14(n10686), .ROB13(n10685), .ROB12(n10684), 
            .ROB11(n10683), .ROB10(n10682), .ROB9(n10681), .ROB8(n10680), 
            .ROB7(n10679), .ROB6(n10678), .ROB5(n10677), .ROB4(n10676), 
            .ROB3(n10675), .ROB2(n10674), .ROB1(n10673), .ROB0(n10672), 
            .P35(n10726), .P34(n10725), .P33(n10724), .P32(n10723), 
            .P31(n10722), .P30(n10721), .P29(n10720), .P28(n10719), 
            .P27(n10718), .P26(n10717), .P25(n10716), .P24(n10715), 
            .P23(n10714), .P22(n10713), .P21(n10712), .P20(n10711), 
            .P19(n10710), .P18(n10709), .P17(n10708), .P16(n10707), 
            .P15(n10706), .P14(n10705), .P13(n10704), .P12(n10703), 
            .P11(n10702), .P10(n10701), .P9(n10700), .P8(n10699), .P7(n10698), 
            .P6(n10697), .P5(n10696), .P4(n10695), .P3(n10694), .P2(n10693), 
            .P1(n10692), .P0(n10691), .SIGNEDP(n10690));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[44:57])
    defparam lat_mult_5.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_5.REG_INPUTA_CE = "CE3";
    defparam lat_mult_5.REG_INPUTA_RST = "RST3";
    defparam lat_mult_5.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTB_CE = "CE0";
    defparam lat_mult_5.REG_INPUTB_RST = "RST0";
    defparam lat_mult_5.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTC_CE = "CE0";
    defparam lat_mult_5.REG_INPUTC_RST = "RST0";
    defparam lat_mult_5.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_5.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_5.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_5.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_5.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_5.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_5.CLK0_DIV = "ENABLED";
    defparam lat_mult_5.CLK1_DIV = "ENABLED";
    defparam lat_mult_5.CLK2_DIV = "ENABLED";
    defparam lat_mult_5.CLK3_DIV = "ENABLED";
    defparam lat_mult_5.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_5.GSR = "DISABLED";
    defparam lat_mult_5.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_5.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_5.MULT_BYPASS = "DISABLED";
    defparam lat_mult_5.RESETMODE = "ASYNC";
    MULT18X18D b_s_31__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[15]), .B14(b_s[14]), .B13(b_s[13]), .B12(b_s[12]), 
            .B11(b_s[11]), .B10(b_s[10]), .B9(b_s[9]), .B8(b_s[8]), 
            .B7(b_s[7]), .B6(b_s[6]), .B5(b_s[5]), .B4(b_s[4]), .B3(b_s[3]), 
            .B2(b_s[2]), .B1(b_s[1]), .B0(b_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10598), .ROA16(n10597), .ROA15(n10596), .ROA14(n10595), 
            .ROA13(n10594), .ROA12(n10593), .ROA11(n10592), .ROA10(n10591), 
            .ROA9(n10590), .ROA8(n10589), .ROA7(n10588), .ROA6(n10587), 
            .ROA5(n10586), .ROA4(n10585), .ROA3(n10584), .ROA2(n10583), 
            .ROA1(n10582), .ROA0(n10581), .ROB17(n10616), .ROB16(n10615), 
            .ROB15(n10614), .ROB14(n10613), .ROB13(n10612), .ROB12(n10611), 
            .ROB11(n10610), .ROB10(n10609), .ROB9(n10608), .ROB8(n10607), 
            .ROB7(n10606), .ROB6(n10605), .ROB5(n10604), .ROB4(n10603), 
            .ROB3(n10602), .ROB2(n10601), .ROB1(n10600), .ROB0(n10599), 
            .P35(n10653), .P34(n10652), .P33(n10651), .P32(n10650), 
            .P31(n10649), .P30(n10648), .P29(n10647), .P28(n10646), 
            .P27(n10645), .P26(n10644), .P25(n10643), .P24(n10642), 
            .P23(n10641), .P22(n10640), .P21(n10639), .P20(n10638), 
            .P19(n10637), .P18(n10636), .P17(n10635), .P16(n10634), 
            .P15(n10633), .P14(n10632), .P13(n10631), .P12(n10630), 
            .P11(n10629), .P10(n10628), .P9(n10627), .P8(n10626), .P7(n10625), 
            .P6(n10624), .P5(n10623), .P4(n10622), .P3(n10621), .P2(n10620), 
            .P1(n10619), .P0(n10618), .SIGNEDP(n10617));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(102[44:57])
    defparam b_s_31__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam b_s_31__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam b_s_31__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam b_s_31__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam b_s_31__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam b_s_31__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam b_s_31__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam b_s_31__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.GSR = "DISABLED";
    defparam b_s_31__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam b_s_31__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam b_s_31__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam b_s_31__I_0_mult_2.RESETMODE = "ASYNC";
    ALU54B lat_alu_4 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10403), .SIGNEDIB(n10476), .SIGNEDCIN(n10549), .A35(n10402), 
           .A34(n10401), .A33(n10400), .A32(n10399), .A31(n10398), .A30(n10397), 
           .A29(n10396), .A28(n10395), .A27(n10394), .A26(n10393), .A25(n10392), 
           .A24(n10391), .A23(n10390), .A22(n10389), .A21(n10388), .A20(n10387), 
           .A19(n10386), .A18(n10385), .A17(n10384), .A16(n10383), .A15(n10382), 
           .A14(n10381), .A13(n10380), .A12(n10379), .A11(n10378), .A10(n10377), 
           .A9(n10376), .A8(n10375), .A7(n10374), .A6(n10373), .A5(n10372), 
           .A4(n10371), .A3(n10370), .A2(n10369), .A1(n10368), .A0(n10367), 
           .B35(n10475), .B34(n10474), .B33(n10473), .B32(n10472), .B31(n10471), 
           .B30(n10470), .B29(n10469), .B28(n10468), .B27(n10467), .B26(n10466), 
           .B25(n10465), .B24(n10464), .B23(n10463), .B22(n10462), .B21(n10461), 
           .B20(n10460), .B19(n10459), .B18(n10458), .B17(n10457), .B16(n10456), 
           .B15(n10455), .B14(n10454), .B13(n10453), .B12(n10452), .B11(n10451), 
           .B10(n10450), .B9(n10449), .B8(n10448), .B7(n10447), .B6(n10446), 
           .B5(n10445), .B4(n10444), .B3(n10443), .B2(n10442), .B1(n10441), 
           .B0(n10440), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10439), .MA34(n10438), .MA33(n10437), .MA32(n10436), 
           .MA31(n10435), .MA30(n10434), .MA29(n10433), .MA28(n10432), 
           .MA27(n10431), .MA26(n10430), .MA25(n10429), .MA24(n10428), 
           .MA23(n10427), .MA22(n10426), .MA21(n10425), .MA20(n10424), 
           .MA19(n10423), .MA18(n10422), .MA17(n10421), .MA16(n10420), 
           .MA15(n10419), .MA14(n10418), .MA13(n10417), .MA12(n10416), 
           .MA11(n10415), .MA10(n10414), .MA9(n10413), .MA8(n10412), 
           .MA7(n10411), .MA6(n10410), .MA5(n10409), .MA4(n10408), .MA3(n10407), 
           .MA2(n10406), .MA1(n10405), .MA0(n10404), .MB35(n10512), 
           .MB34(n10511), .MB33(n10510), .MB32(n10509), .MB31(n10508), 
           .MB30(n10507), .MB29(n10506), .MB28(n10505), .MB27(n10504), 
           .MB26(n10503), .MB25(n10502), .MB24(n10501), .MB23(n10500), 
           .MB22(n10499), .MB21(n10498), .MB20(n10497), .MB19(n10496), 
           .MB18(n10495), .MB17(n10494), .MB16(n10493), .MB15(n10492), 
           .MB14(n10491), .MB13(n10490), .MB12(n10489), .MB11(n10488), 
           .MB10(n10487), .MB9(n10486), .MB8(n10485), .MB7(n10484), 
           .MB6(n10483), .MB5(n10482), .MB4(n10481), .MB3(n10480), .MB2(n10479), 
           .MB1(n10478), .MB0(n10477), .CIN53(n10548), .CIN52(n10547), 
           .CIN51(n10546), .CIN50(n10545), .CIN49(n10544), .CIN48(n10543), 
           .CIN47(n10542), .CIN46(n10541), .CIN45(n10540), .CIN44(n10539), 
           .CIN43(n10538), .CIN42(n10537), .CIN41(n10536), .CIN40(n10535), 
           .CIN39(n10534), .CIN38(n10533), .CIN37(n10532), .CIN36(n10531), 
           .CIN35(n10530), .CIN34(n10529), .CIN33(n10528), .CIN32(n10527), 
           .CIN31(n10526), .CIN30(n10525), .CIN29(n10524), .CIN28(n10523), 
           .CIN27(n10522), .CIN26(n10521), .CIN25(n10520), .CIN24(n10519), 
           .CIN23(n10518), .CIN22(n10517), .CIN21(n10516), .CIN20(n10515), 
           .CIN19(n10514), .CIN18(n10513), .CIN17(prod_a[17]), .CIN16(prod_a[16]), 
           .CIN15(prod_a[15]), .CIN14(n10206), .CIN13(n10207), .CIN12(n10208), 
           .CIN11(n10209), .CIN10(n10210), .CIN9(n10211), .CIN8(n10212), 
           .CIN7(n10213), .CIN6(n10214), .CIN5(n10215), .CIN4(n10216), 
           .CIN3(n10217), .CIN2(n10218), .CIN1(n10219), .CIN0(n10220), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R29(prod_a[47]), 
           .R28(prod_a[46]), .R27(prod_a[45]), .R26(prod_a[44]), .R25(prod_a[43]), 
           .R24(prod_a[42]), .R23(prod_a[41]), .R22(prod_a[40]), .R21(prod_a[39]), 
           .R20(prod_a[38]), .R19(prod_a[37]), .R18(prod_a[36]), .R17(prod_a[35]), 
           .R16(prod_a[34]), .R15(prod_a[33]), .R14(prod_a[32]), .R13(prod_a[31]), 
           .R12(prod_a[30]), .R11(prod_a[29]), .R10(prod_a[28]), .R9(prod_a[27]), 
           .R8(prod_a[26]), .R7(prod_a[25]), .R6(prod_a[24]), .R5(prod_a[23]), 
           .R4(prod_a[22]), .R3(prod_a[21]), .R2(prod_a[20]), .R1(prod_a[19]), 
           .R0(prod_a[18]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam lat_alu_4.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_4.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_4.REG_FLAG_CLK = "NONE";
    defparam lat_alu_4.REG_FLAG_CE = "CE0";
    defparam lat_alu_4.REG_FLAG_RST = "RST0";
    defparam lat_alu_4.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASK01 = "0x00000000000000";
    defparam lat_alu_4.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_4.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_4.CLK0_DIV = "ENABLED";
    defparam lat_alu_4.CLK1_DIV = "ENABLED";
    defparam lat_alu_4.CLK2_DIV = "ENABLED";
    defparam lat_alu_4.CLK3_DIV = "ENABLED";
    defparam lat_alu_4.MCPAT = "0x00000000000000";
    defparam lat_alu_4.MASKPAT = "0x00000000000000";
    defparam lat_alu_4.RNDPAT = "0x00000000000000";
    defparam lat_alu_4.GSR = "DISABLED";
    defparam lat_alu_4.RESETMODE = "SYNC";
    defparam lat_alu_4.MULT9_MODE = "DISABLED";
    defparam lat_alu_4.LEGACY = "DISABLED";
    ALU54B lat_alu_3 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10257), .SIGNEDIB(n10330), .SIGNEDCIN(GND_net), 
           .A35(n10256), .A34(n10255), .A33(n10254), .A32(n10253), .A31(n10252), 
           .A30(n10251), .A29(n10250), .A28(n10249), .A27(n10248), .A26(n10247), 
           .A25(n10246), .A24(n10245), .A23(n10244), .A22(n10243), .A21(n10242), 
           .A20(n10241), .A19(n10240), .A18(n10239), .A17(n10238), .A16(n10237), 
           .A15(n10236), .A14(n10235), .A13(n10234), .A12(n10233), .A11(n10232), 
           .A10(n10231), .A9(n10230), .A8(n10229), .A7(n10228), .A6(n10227), 
           .A5(n10226), .A4(n10225), .A3(n10224), .A2(n10223), .A1(n10222), 
           .A0(n10221), .B35(n10329), .B34(n10328), .B33(n10327), .B32(n10326), 
           .B31(n10325), .B30(n10324), .B29(n10323), .B28(n10322), .B27(n10321), 
           .B26(n10320), .B25(n10319), .B24(n10318), .B23(n10317), .B22(n10316), 
           .B21(n10315), .B20(n10314), .B19(n10313), .B18(n10312), .B17(n10311), 
           .B16(n10310), .B15(n10309), .B14(n10308), .B13(n10307), .B12(n10306), 
           .B11(n10305), .B10(n10304), .B9(n10303), .B8(n10302), .B7(n10301), 
           .B6(n10300), .B5(n10299), .B4(n10298), .B3(n10297), .B2(n10296), 
           .B1(n10295), .B0(n10294), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10293), .MA34(n10292), .MA33(n10291), .MA32(n10290), 
           .MA31(n10289), .MA30(n10288), .MA29(n10287), .MA28(n10286), 
           .MA27(n10285), .MA26(n10284), .MA25(n10283), .MA24(n10282), 
           .MA23(n10281), .MA22(n10280), .MA21(n10279), .MA20(n10278), 
           .MA19(n10277), .MA18(n10276), .MA17(n10275), .MA16(n10274), 
           .MA15(n10273), .MA14(n10272), .MA13(n10271), .MA12(n10270), 
           .MA11(n10269), .MA10(n10268), .MA9(n10267), .MA8(n10266), 
           .MA7(n10265), .MA6(n10264), .MA5(n10263), .MA4(n10262), .MA3(n10261), 
           .MA2(n10260), .MA1(n10259), .MA0(n10258), .MB35(n10366), 
           .MB34(n10365), .MB33(n10364), .MB32(n10363), .MB31(n10362), 
           .MB30(n10361), .MB29(n10360), .MB28(n10359), .MB27(n10358), 
           .MB26(n10357), .MB25(n10356), .MB24(n10355), .MB23(n10354), 
           .MB22(n10353), .MB21(n10352), .MB20(n10351), .MB19(n10350), 
           .MB18(n10349), .MB17(n10348), .MB16(n10347), .MB15(n10346), 
           .MB14(n10345), .MB13(n10344), .MB12(n10343), .MB11(n10342), 
           .MB10(n10341), .MB9(n10340), .MB8(n10339), .MB7(n10338), 
           .MB6(n10337), .MB5(n10336), .MB4(n10335), .MB3(n10334), .MB2(n10333), 
           .MB1(n10332), .MB0(n10331), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n10548), 
           .R52(n10547), .R51(n10546), .R50(n10545), .R49(n10544), .R48(n10543), 
           .R47(n10542), .R46(n10541), .R45(n10540), .R44(n10539), .R43(n10538), 
           .R42(n10537), .R41(n10536), .R40(n10535), .R39(n10534), .R38(n10533), 
           .R37(n10532), .R36(n10531), .R35(n10530), .R34(n10529), .R33(n10528), 
           .R32(n10527), .R31(n10526), .R30(n10525), .R29(n10524), .R28(n10523), 
           .R27(n10522), .R26(n10521), .R25(n10520), .R24(n10519), .R23(n10518), 
           .R22(n10517), .R21(n10516), .R20(n10515), .R19(n10514), .R18(n10513), 
           .R17(prod_a[17]), .R16(prod_a[16]), .R15(prod_a[15]), .R14(n10206), 
           .R13(n10207), .R12(n10208), .R11(n10209), .R10(n10210), .R9(n10211), 
           .R8(n10212), .R7(n10213), .R6(n10214), .R5(n10215), .R4(n10216), 
           .R3(n10217), .R2(n10218), .R1(n10219), .R0(n10220), .SIGNEDR(n10549));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam lat_alu_3.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_3.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_3.REG_FLAG_CLK = "NONE";
    defparam lat_alu_3.REG_FLAG_CE = "CE0";
    defparam lat_alu_3.REG_FLAG_RST = "RST0";
    defparam lat_alu_3.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASK01 = "0x00000000000000";
    defparam lat_alu_3.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_3.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_3.CLK0_DIV = "ENABLED";
    defparam lat_alu_3.CLK1_DIV = "ENABLED";
    defparam lat_alu_3.CLK2_DIV = "ENABLED";
    defparam lat_alu_3.CLK3_DIV = "ENABLED";
    defparam lat_alu_3.MCPAT = "0x00000000000000";
    defparam lat_alu_3.MASKPAT = "0x00000000000000";
    defparam lat_alu_3.RNDPAT = "0x00000000000000";
    defparam lat_alu_3.GSR = "DISABLED";
    defparam lat_alu_3.RESETMODE = "SYNC";
    defparam lat_alu_3.MULT9_MODE = "DISABLED";
    defparam lat_alu_3.LEGACY = "DISABLED";
    FD1S3AX d_inv_reg_res4_i16 (.D(d_inv_15__N_49[47]), .CK(clk_c), .Q(d_inv_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i16.GSR = "ENABLED";
    MULT18X18D lat_mult_2 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68_adj_245), .B16(n68_adj_245), 
            .B15(n68_adj_245), .B14(n68_adj_245), .B13(n68_adj_245), .B12(n68_adj_245), 
            .B11(n68_adj_245), .B10(n68_adj_245), .B9(n68_adj_245), .B8(n68_adj_245), 
            .B7(n68_adj_245), .B6(n68_adj_245), .B5(n68_adj_245), .B4(n68_adj_245), 
            .B3(n68_adj_245), .B2(n68_adj_245), .B1(n68_adj_245), .B0(n68_adj_245), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10457), .ROA16(n10456), 
            .ROA15(n10455), .ROA14(n10454), .ROA13(n10453), .ROA12(n10452), 
            .ROA11(n10451), .ROA10(n10450), .ROA9(n10449), .ROA8(n10448), 
            .ROA7(n10447), .ROA6(n10446), .ROA5(n10445), .ROA4(n10444), 
            .ROA3(n10443), .ROA2(n10442), .ROA1(n10441), .ROA0(n10440), 
            .ROB17(n10475), .ROB16(n10474), .ROB15(n10473), .ROB14(n10472), 
            .ROB13(n10471), .ROB12(n10470), .ROB11(n10469), .ROB10(n10468), 
            .ROB9(n10467), .ROB8(n10466), .ROB7(n10465), .ROB6(n10464), 
            .ROB5(n10463), .ROB4(n10462), .ROB3(n10461), .ROB2(n10460), 
            .ROB1(n10459), .ROB0(n10458), .P35(n10512), .P34(n10511), 
            .P33(n10510), .P32(n10509), .P31(n10508), .P30(n10507), 
            .P29(n10506), .P28(n10505), .P27(n10504), .P26(n10503), 
            .P25(n10502), .P24(n10501), .P23(n10500), .P22(n10499), 
            .P21(n10498), .P20(n10497), .P19(n10496), .P18(n10495), 
            .P17(n10494), .P16(n10493), .P15(n10492), .P14(n10491), 
            .P13(n10490), .P12(n10489), .P11(n10488), .P10(n10487), 
            .P9(n10486), .P8(n10485), .P7(n10484), .P6(n10483), .P5(n10482), 
            .P4(n10481), .P3(n10480), .P2(n10479), .P1(n10478), .P0(n10477), 
            .SIGNEDP(n10476));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam lat_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_2.REG_INPUTA_CE = "CE3";
    defparam lat_mult_2.REG_INPUTA_RST = "RST3";
    defparam lat_mult_2.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTB_CE = "CE0";
    defparam lat_mult_2.REG_INPUTB_RST = "RST0";
    defparam lat_mult_2.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTC_CE = "CE0";
    defparam lat_mult_2.REG_INPUTC_RST = "RST0";
    defparam lat_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_2.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_2.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_2.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_2.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_2.CLK0_DIV = "ENABLED";
    defparam lat_mult_2.CLK1_DIV = "ENABLED";
    defparam lat_mult_2.CLK2_DIV = "ENABLED";
    defparam lat_mult_2.CLK3_DIV = "ENABLED";
    defparam lat_mult_2.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_2.GSR = "DISABLED";
    defparam lat_mult_2.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_2.MULT_BYPASS = "DISABLED";
    defparam lat_mult_2.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_1 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(n68_adj_245), .B16(n68_adj_245), 
            .B15(n68_adj_245), .B14(n68_adj_245), .B13(n68_adj_245), .B12(n68_adj_245), 
            .B11(n68_adj_245), .B10(n68_adj_245), .B9(n68_adj_245), .B8(n68_adj_245), 
            .B7(n68_adj_245), .B6(n68_adj_245), .B5(n68_adj_245), .B4(n68_adj_245), 
            .B3(n68_adj_245), .B2(n68_adj_245), .B1(n68_adj_245), .B0(n68_adj_245), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10384), .ROA16(n10383), 
            .ROA15(n10382), .ROA14(n10381), .ROA13(n10380), .ROA12(n10379), 
            .ROA11(n10378), .ROA10(n10377), .ROA9(n10376), .ROA8(n10375), 
            .ROA7(n10374), .ROA6(n10373), .ROA5(n10372), .ROA4(n10371), 
            .ROA3(n10370), .ROA2(n10369), .ROA1(n10368), .ROA0(n10367), 
            .ROB17(n10402), .ROB16(n10401), .ROB15(n10400), .ROB14(n10399), 
            .ROB13(n10398), .ROB12(n10397), .ROB11(n10396), .ROB10(n10395), 
            .ROB9(n10394), .ROB8(n10393), .ROB7(n10392), .ROB6(n10391), 
            .ROB5(n10390), .ROB4(n10389), .ROB3(n10388), .ROB2(n10387), 
            .ROB1(n10386), .ROB0(n10385), .P35(n10439), .P34(n10438), 
            .P33(n10437), .P32(n10436), .P31(n10435), .P30(n10434), 
            .P29(n10433), .P28(n10432), .P27(n10431), .P26(n10430), 
            .P25(n10429), .P24(n10428), .P23(n10427), .P22(n10426), 
            .P21(n10425), .P20(n10424), .P19(n10423), .P18(n10422), 
            .P17(n10421), .P16(n10420), .P15(n10419), .P14(n10418), 
            .P13(n10417), .P12(n10416), .P11(n10415), .P10(n10414), 
            .P9(n10413), .P8(n10412), .P7(n10411), .P6(n10410), .P5(n10409), 
            .P4(n10408), .P3(n10407), .P2(n10406), .P1(n10405), .P0(n10404), 
            .SIGNEDP(n10403));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam lat_mult_1.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_1.REG_INPUTA_CE = "CE3";
    defparam lat_mult_1.REG_INPUTA_RST = "RST3";
    defparam lat_mult_1.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTB_CE = "CE0";
    defparam lat_mult_1.REG_INPUTB_RST = "RST0";
    defparam lat_mult_1.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTC_CE = "CE0";
    defparam lat_mult_1.REG_INPUTC_RST = "RST0";
    defparam lat_mult_1.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_1.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_1.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_1.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_1.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_1.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_1.CLK0_DIV = "ENABLED";
    defparam lat_mult_1.CLK1_DIV = "ENABLED";
    defparam lat_mult_1.CLK2_DIV = "ENABLED";
    defparam lat_mult_1.CLK3_DIV = "ENABLED";
    defparam lat_mult_1.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_1.GSR = "DISABLED";
    defparam lat_mult_1.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_1.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_1.MULT_BYPASS = "DISABLED";
    defparam lat_mult_1.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_0 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68_adj_245), .B16(n68_adj_245), 
            .B15(n68_adj_245), .B14(n102_adj_244), .B13(n104_adj_243), 
            .B12(n106_adj_230), .B11(n108_adj_242), .B10(n110_adj_241), 
            .B9(n112_adj_240), .B8(n114_adj_239), .B7(n116_adj_238), .B6(n118_adj_237), 
            .B5(n120_adj_236), .B4(n122_adj_235), .B3(n124_adj_234), .B2(n126_adj_233), 
            .B1(n128_adj_232), .B0(n130_adj_231), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10311), .ROA16(n10310), .ROA15(n10309), .ROA14(n10308), 
            .ROA13(n10307), .ROA12(n10306), .ROA11(n10305), .ROA10(n10304), 
            .ROA9(n10303), .ROA8(n10302), .ROA7(n10301), .ROA6(n10300), 
            .ROA5(n10299), .ROA4(n10298), .ROA3(n10297), .ROA2(n10296), 
            .ROA1(n10295), .ROA0(n10294), .ROB17(n10329), .ROB16(n10328), 
            .ROB15(n10327), .ROB14(n10326), .ROB13(n10325), .ROB12(n10324), 
            .ROB11(n10323), .ROB10(n10322), .ROB9(n10321), .ROB8(n10320), 
            .ROB7(n10319), .ROB6(n10318), .ROB5(n10317), .ROB4(n10316), 
            .ROB3(n10315), .ROB2(n10314), .ROB1(n10313), .ROB0(n10312), 
            .P35(n10366), .P34(n10365), .P33(n10364), .P32(n10363), 
            .P31(n10362), .P30(n10361), .P29(n10360), .P28(n10359), 
            .P27(n10358), .P26(n10357), .P25(n10356), .P24(n10355), 
            .P23(n10354), .P22(n10353), .P21(n10352), .P20(n10351), 
            .P19(n10350), .P18(n10349), .P17(n10348), .P16(n10347), 
            .P15(n10346), .P14(n10345), .P13(n10344), .P12(n10343), 
            .P11(n10342), .P10(n10341), .P9(n10340), .P8(n10339), .P7(n10338), 
            .P6(n10337), .P5(n10336), .P4(n10335), .P3(n10334), .P2(n10333), 
            .P1(n10332), .P0(n10331), .SIGNEDP(n10330));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam lat_mult_0.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_0.REG_INPUTA_CE = "CE3";
    defparam lat_mult_0.REG_INPUTA_RST = "RST3";
    defparam lat_mult_0.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTB_CE = "CE0";
    defparam lat_mult_0.REG_INPUTB_RST = "RST0";
    defparam lat_mult_0.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTC_CE = "CE0";
    defparam lat_mult_0.REG_INPUTC_RST = "RST0";
    defparam lat_mult_0.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_0.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_0.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_0.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_0.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_0.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_0.CLK0_DIV = "ENABLED";
    defparam lat_mult_0.CLK1_DIV = "ENABLED";
    defparam lat_mult_0.CLK2_DIV = "ENABLED";
    defparam lat_mult_0.CLK3_DIV = "ENABLED";
    defparam lat_mult_0.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_0.GSR = "DISABLED";
    defparam lat_mult_0.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_0.MULT_BYPASS = "DISABLED";
    defparam lat_mult_0.RESETMODE = "ASYNC";
    MULT18X18D d2_reg_15__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), 
            .A14(n50), .A13(n51), .A12(n52), .A11(n53), .A10(n54), 
            .A9(n55), .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), 
            .A3(n61), .A2(n62), .A1(n63), .A0(n64), .B17(n68_adj_245), 
            .B16(n68_adj_245), .B15(n68_adj_245), .B14(n102_adj_244), 
            .B13(n104_adj_243), .B12(n106_adj_230), .B11(n108_adj_242), 
            .B10(n110_adj_241), .B9(n112_adj_240), .B8(n114_adj_239), 
            .B7(n116_adj_238), .B6(n118_adj_237), .B5(n120_adj_236), .B4(n122_adj_235), 
            .B3(n124_adj_234), .B2(n126_adj_233), .B1(n128_adj_232), .B0(n130_adj_231), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10238), .ROA16(n10237), 
            .ROA15(n10236), .ROA14(n10235), .ROA13(n10234), .ROA12(n10233), 
            .ROA11(n10232), .ROA10(n10231), .ROA9(n10230), .ROA8(n10229), 
            .ROA7(n10228), .ROA6(n10227), .ROA5(n10226), .ROA4(n10225), 
            .ROA3(n10224), .ROA2(n10223), .ROA1(n10222), .ROA0(n10221), 
            .ROB17(n10256), .ROB16(n10255), .ROB15(n10254), .ROB14(n10253), 
            .ROB13(n10252), .ROB12(n10251), .ROB11(n10250), .ROB10(n10249), 
            .ROB9(n10248), .ROB8(n10247), .ROB7(n10246), .ROB6(n10245), 
            .ROB5(n10244), .ROB4(n10243), .ROB3(n10242), .ROB2(n10241), 
            .ROB1(n10240), .ROB0(n10239), .P35(n10293), .P34(n10292), 
            .P33(n10291), .P32(n10290), .P31(n10289), .P30(n10288), 
            .P29(n10287), .P28(n10286), .P27(n10285), .P26(n10284), 
            .P25(n10283), .P24(n10282), .P23(n10281), .P22(n10280), 
            .P21(n10279), .P20(n10278), .P19(n10277), .P18(n10276), 
            .P17(n10275), .P16(n10274), .P15(n10273), .P14(n10272), 
            .P13(n10271), .P12(n10270), .P11(n10269), .P10(n10268), 
            .P9(n10267), .P8(n10266), .P7(n10265), .P6(n10264), .P5(n10263), 
            .P4(n10262), .P3(n10261), .P2(n10260), .P1(n10259), .P0(n10258), 
            .SIGNEDP(n10257));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam d2_reg_15__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam d2_reg_15__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam d2_reg_15__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam d2_reg_15__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam d2_reg_15__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam d2_reg_15__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam d2_reg_15__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam d2_reg_15__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam d2_reg_15__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam d2_reg_15__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam d2_reg_15__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam d2_reg_15__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam d2_reg_15__I_0_mult_2.GSR = "DISABLED";
    defparam d2_reg_15__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam d2_reg_15__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam d2_reg_15__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam d2_reg_15__I_0_mult_2.RESETMODE = "ASYNC";
    FD1S3AX d_inv_reg_res4_i9 (.D(d_inv_15__N_49[40]), .CK(clk_c), .Q(d_inv_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i9.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i10 (.D(d_inv_15__N_49[41]), .CK(clk_c), .Q(d_inv_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i10.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i13 (.D(d_inv_15__N_49[44]), .CK(clk_c), .Q(d_inv_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i13.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i14 (.D(d_inv_15__N_49[45]), .CK(clk_c), .Q(d_inv_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i14.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i15 (.D(d_inv_15__N_49[46]), .CK(clk_c), .Q(d_inv_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i15.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i2 (.D(d_inv_15__N_49[33]), .CK(clk_c), .Q(d_inv_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i2.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i3 (.D(d_inv_15__N_49[34]), .CK(clk_c), .Q(d_inv_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i3.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i12 (.D(d_inv_15__N_49[43]), .CK(clk_c), .Q(d_inv_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i12.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i11 (.D(d_inv_15__N_49[42]), .CK(clk_c), .Q(d_inv_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i11.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i6 (.D(d_inv_15__N_49[37]), .CK(clk_c), .Q(d_inv_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i6.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i7 (.D(d_inv_15__N_49[38]), .CK(clk_c), .Q(d_inv_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i7.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i8 (.D(d_inv_15__N_49[39]), .CK(clk_c), .Q(d_inv_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i8.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i10 (.D(a_inv_15__N_1[41]), .CK(clk_c), .Q(a_inv_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i10.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i11 (.D(a_inv_15__N_1[42]), .CK(clk_c), .Q(a_inv_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i11.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i5 (.D(d_inv_15__N_49[36]), .CK(clk_c), .Q(d_inv_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i5.GSR = "ENABLED";
    FD1S3AX d_inv_reg_res4_i4 (.D(d_inv_15__N_49[35]), .CK(clk_c), .Q(d_inv_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam d_inv_reg_res4_i4.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i14 (.D(a_inv_15__N_1[45]), .CK(clk_c), .Q(a_inv_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i14.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i15 (.D(a_inv_15__N_1[46]), .CK(clk_c), .Q(a_inv_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i15.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i16 (.D(a_inv_15__N_1[47]), .CK(clk_c), .Q(a_inv_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i16.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i3 (.D(a_inv_15__N_1[34]), .CK(clk_c), .Q(a_inv_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i3.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i4 (.D(a_inv_15__N_1[35]), .CK(clk_c), .Q(a_inv_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i4.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i13 (.D(a_inv_15__N_1[44]), .CK(clk_c), .Q(a_inv_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i13.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i12 (.D(a_inv_15__N_1[43]), .CK(clk_c), .Q(a_inv_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i12.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i7 (.D(a_inv_15__N_1[38]), .CK(clk_c), .Q(a_inv_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i7.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i8 (.D(a_inv_15__N_1[39]), .CK(clk_c), .Q(a_inv_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i8.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i9 (.D(a_inv_15__N_1[40]), .CK(clk_c), .Q(a_inv_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i9.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i6 (.D(a_inv_15__N_1[37]), .CK(clk_c), .Q(a_inv_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i6.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i5 (.D(a_inv_15__N_1[36]), .CK(clk_c), .Q(a_inv_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i5.GSR = "ENABLED";
    FD1S3AX a_inv_reg_res3_i2 (.D(a_inv_15__N_1[33]), .CK(clk_c), .Q(a_inv_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam a_inv_reg_res3_i2.GSR = "ENABLED";
    FD1S3AX c1_reg_i3 (.D(c_c_3), .CK(clk_c), .Q(c1_reg[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i3.GSR = "ENABLED";
    OB b_inv_pad_3 (.I(b_inv_c_3), .O(b_inv[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_4 (.I(b_inv_c_4), .O(b_inv[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_5 (.I(b_inv_c_5), .O(b_inv[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_6 (.I(b_inv_c_6), .O(b_inv[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB a_inv_pad_6 (.I(a_inv_c_6), .O(a_inv[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB b_inv_pad_7 (.I(b_inv_c_7), .O(b_inv[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB a_inv_pad_5 (.I(a_inv_c_5), .O(a_inv[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_4 (.I(a_inv_c_4), .O(a_inv[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_0 (.I(a_inv_c_0), .O(a_inv[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    LUT4 i1344_2_lut (.A(n1475), .B(det_q4_28[0]), .Z(n161_adj_1366)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1344_2_lut.init = 16'h6666;
    IB b_pad_7 (.I(b[7]), .O(b_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_8 (.I(b[8]), .O(b_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    FD1S3AX c1_reg_i2 (.D(c_c_2), .CK(clk_c), .Q(c1_reg[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i2.GSR = "ENABLED";
    FD1S3AX det_q4_28_i28 (.D(det_q4_28_31__N_65[28]), .CK(clk_c), .Q(det_q4_28[28]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i28.GSR = "ENABLED";
    CCU2C _add_1_add_4_9 (.A0(n143_adj_1519), .B0(n2583), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1518), .B1(n2583), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12597), .COUT(n12598), .S0(n140_adj_371), 
          .S1(n137_adj_370));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_add_4_9.INJECT1_1 = "NO";
    OB a_inv_pad_2 (.I(a_inv_c_2), .O(a_inv[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_14 (.I(a_inv_c_14), .O(a_inv[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_13 (.I(a_inv_c_13), .O(a_inv[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_3 (.I(a_inv_c_3), .O(a_inv[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB c_inv_pad_8 (.I(c_inv_c_8), .O(c_inv[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB a_inv_pad_12 (.I(a_inv_c_12), .O(a_inv[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_11 (.I(a_inv_c_11), .O(a_inv[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB a_inv_pad_8 (.I(a_inv_c_8), .O(a_inv[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    LUT4 mux_343_i1_3_lut_rep_68 (.A(n68_adj_474), .B(n68_adj_442), .C(n2650), 
         .Z(n13818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_343_i1_3_lut_rep_68.init = 16'hcaca;
    LUT4 mux_341_i1_3_lut_rep_70 (.A(n68_adj_602), .B(n68_adj_570), .C(n2650), 
         .Z(n13820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_341_i1_3_lut_rep_70.init = 16'hcaca;
    OB b_inv_pad_8 (.I(b_inv_c_8), .O(b_inv[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_9 (.I(b_inv_c_9), .O(b_inv[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    LUT4 mux_340_i1_3_lut_rep_71 (.A(n68_adj_666), .B(n68_adj_634), .C(n2650), 
         .Z(n13821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_340_i1_3_lut_rep_71.init = 16'hcaca;
    LUT4 i1504_2_lut_4_lut (.A(n68_adj_666), .B(n68_adj_634), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n58)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1504_2_lut_4_lut.init = 16'h0035;
    OB b_inv_pad_10 (.I(b_inv_c_10), .O(b_inv[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_11 (.I(b_inv_c_11), .O(b_inv[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_2 (.I(b_inv_c_2), .O(b_inv[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    LUT4 mux_339_i1_3_lut_rep_72 (.A(n68_adj_730), .B(n68_adj_698), .C(n2650), 
         .Z(n13822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_339_i1_3_lut_rep_72.init = 16'hcaca;
    LUT4 i1507_2_lut_4_lut (.A(n68_adj_730), .B(n68_adj_698), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n57)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1507_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_338_i1_3_lut_rep_73 (.A(n68_adj_826), .B(n68_adj_762), .C(n2650), 
         .Z(n13823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_338_i1_3_lut_rep_73.init = 16'hcaca;
    LUT4 i1510_2_lut_4_lut (.A(n68_adj_826), .B(n68_adj_762), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n56)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1510_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_337_i1_3_lut_rep_74 (.A(n68_adj_1717), .B(n68_adj_1685), .C(n2650), 
         .Z(n13824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_337_i1_3_lut_rep_74.init = 16'hcaca;
    LUT4 i1513_2_lut_4_lut (.A(n68_adj_1717), .B(n68_adj_1685), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n55)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1513_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_336_i1_3_lut_rep_75 (.A(n68_adj_1908), .B(n68_adj_1844), .C(n2650), 
         .Z(n13825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_336_i1_3_lut_rep_75.init = 16'hcaca;
    FD1S3AX det_q4_28_i29 (.D(det_q4_28_31__N_65[29]), .CK(clk_c), .Q(det_q4_28[29]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i29.GSR = "ENABLED";
    FD1S3AX det_q4_28_i21 (.D(det_q4_28_31__N_65[21]), .CK(clk_c), .Q(det_q4_28[21]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i21.GSR = "ENABLED";
    LUT4 i1516_2_lut_4_lut (.A(n68_adj_1908), .B(n68_adj_1844), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n54)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1516_2_lut_4_lut.init = 16'h0035;
    LUT4 i1501_2_lut_4_lut (.A(n68_adj_602), .B(n68_adj_570), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n59)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1501_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_335_i1_3_lut_rep_76 (.A(n68_adj_2003), .B(n68_adj_1971), .C(n2650), 
         .Z(n13826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_335_i1_3_lut_rep_76.init = 16'hcaca;
    LUT4 i767_2_lut_4_lut (.A(n68_adj_474), .B(n68_adj_442), .C(n2650), 
         .D(n1444), .Z(n3421)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i767_2_lut_4_lut.init = 16'h3500;
    LUT4 i1519_2_lut_4_lut (.A(n68_adj_2003), .B(n68_adj_1971), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n53)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1519_2_lut_4_lut.init = 16'h0035;
    FD1S3AX det_q4_28_i22 (.D(det_q4_28_31__N_65[22]), .CK(clk_c), .Q(det_q4_28[22]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i22.GSR = "ENABLED";
    FD1S3AX det_q4_28_i31 (.D(det_q4_28_31__N_65[31]), .CK(clk_c), .Q(det_q4_28[31]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i31.GSR = "ENABLED";
    FD1S3AX c1_reg_i1 (.D(c_c_1), .CK(clk_c), .Q(c1_reg[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam c1_reg_i1.GSR = "ENABLED";
    FD1S3AX det_q4_28_i30 (.D(det_q4_28_31__N_65[30]), .CK(clk_c), .Q(det_q4_28[30]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i30.GSR = "ENABLED";
    FD1S3AX det_q4_28_i25 (.D(det_q4_28_31__N_65[25]), .CK(clk_c), .Q(det_q4_28[25]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i25.GSR = "ENABLED";
    FD1S3AX det_q4_28_i26 (.D(det_q4_28_31__N_65[26]), .CK(clk_c), .Q(det_q4_28[26]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i26.GSR = "ENABLED";
    FD1S3AX b1_reg_i15 (.D(b_c_15), .CK(clk_c), .Q(b1_reg[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i15.GSR = "ENABLED";
    FD1S3AX det_q4_28_i27 (.D(det_q4_28_31__N_65[27]), .CK(clk_c), .Q(det_q4_28[27]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i27.GSR = "ENABLED";
    FD1S3AX det_q4_28_i14 (.D(det_q4_28_31__N_65[14]), .CK(clk_c), .Q(det_q4_28[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i14.GSR = "ENABLED";
    FD1S3AX det_q4_28_i15 (.D(det_q4_28_31__N_65[15]), .CK(clk_c), .Q(det_q4_28[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i15.GSR = "ENABLED";
    FD1S3AX det_q4_28_i24 (.D(det_q4_28_31__N_65[24]), .CK(clk_c), .Q(det_q4_28[24]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i24.GSR = "ENABLED";
    FD1S3AX b1_reg_i14 (.D(b_c_14), .CK(clk_c), .Q(b1_reg[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i14.GSR = "ENABLED";
    FD1S3AX det_q4_28_i23 (.D(det_q4_28_31__N_65[23]), .CK(clk_c), .Q(det_q4_28[23]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i23.GSR = "ENABLED";
    FD1S3AX det_q4_28_i18 (.D(det_q4_28_31__N_65[18]), .CK(clk_c), .Q(det_q4_28[18]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i18.GSR = "ENABLED";
    FD1S3AX det_q4_28_i19 (.D(det_q4_28_31__N_65[19]), .CK(clk_c), .Q(det_q4_28[19]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i19.GSR = "ENABLED";
    FD1S3AX b1_reg_i13 (.D(b_c_13), .CK(clk_c), .Q(b1_reg[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i13.GSR = "ENABLED";
    FD1S3AX det_q4_28_i20 (.D(det_q4_28_31__N_65[20]), .CK(clk_c), .Q(det_q4_28[20]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i20.GSR = "ENABLED";
    FD1S3AX det_q4_28_i7 (.D(det_q4_28_31__N_65[7]), .CK(clk_c), .Q(det_q4_28[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i7.GSR = "ENABLED";
    FD1S3AX det_q4_28_i8 (.D(det_q4_28_31__N_65[8]), .CK(clk_c), .Q(det_q4_28[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i8.GSR = "ENABLED";
    FD1S3AX det_q4_28_i17 (.D(det_q4_28_31__N_65[17]), .CK(clk_c), .Q(det_q4_28[17]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i17.GSR = "ENABLED";
    FD1S3AX b1_reg_i12 (.D(b_c_12), .CK(clk_c), .Q(b1_reg[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i12.GSR = "ENABLED";
    FD1S3AX det_q4_28_i16 (.D(det_q4_28_31__N_65[16]), .CK(clk_c), .Q(det_q4_28[16]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i16.GSR = "ENABLED";
    FD1S3AX det_q4_28_i11 (.D(det_q4_28_31__N_65[11]), .CK(clk_c), .Q(det_q4_28[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i11.GSR = "ENABLED";
    FD1S3AX det_q4_28_i12 (.D(det_q4_28_31__N_65[12]), .CK(clk_c), .Q(det_q4_28[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i12.GSR = "ENABLED";
    FD1S3AX b1_reg_i11 (.D(b_c_11), .CK(clk_c), .Q(b1_reg[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i11.GSR = "ENABLED";
    FD1S3AX det_q4_28_i13 (.D(det_q4_28_31__N_65[13]), .CK(clk_c), .Q(det_q4_28[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i13.GSR = "ENABLED";
    FD1S3AX det_q4_28_i10 (.D(det_q4_28_31__N_65[10]), .CK(clk_c), .Q(det_q4_28[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i10.GSR = "ENABLED";
    IB d_pad_5 (.I(d[5]), .O(d_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_4 (.I(d[4]), .O(d_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    FD1S3AX b1_reg_i10 (.D(b_c_10), .CK(clk_c), .Q(b1_reg[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i10.GSR = "ENABLED";
    FD1S3AX det_q4_28_i9 (.D(det_q4_28_31__N_65[9]), .CK(clk_c), .Q(det_q4_28[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i9.GSR = "ENABLED";
    FD1S3AX b1_reg_i9 (.D(b_c_9), .CK(clk_c), .Q(b1_reg[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i9.GSR = "ENABLED";
    IB d_pad_1 (.I(d[1]), .O(d_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_0 (.I(d[0]), .O(d_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    FD1S3AX det_q4_28_i6 (.D(det_q4_28_31__N_65[6]), .CK(clk_c), .Q(det_q4_28[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i6.GSR = "ENABLED";
    FD1S3AX b1_reg_i8 (.D(b_c_8), .CK(clk_c), .Q(b1_reg[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i8.GSR = "ENABLED";
    IB d_pad_12 (.I(d[12]), .O(d_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_11 (.I(d[11]), .O(d_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_2 (.I(d[2]), .O(d_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    FD1S3AX b1_reg_i7 (.D(b_c_7), .CK(clk_c), .Q(b1_reg[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i7.GSR = "ENABLED";
    IB d_pad_3 (.I(d[3]), .O(d_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_8 (.I(d[8]), .O(d_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_7 (.I(d[7]), .O(d_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    FD1S3AX b1_reg_i6 (.D(b_c_6), .CK(clk_c), .Q(b1_reg[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i6.GSR = "ENABLED";
    IB d_pad_6 (.I(d[6]), .O(d_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB c_pad_3 (.I(c[3]), .O(c_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_2 (.I(c[2]), .O(c_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB d_pad_9 (.I(d[9]), .O(d_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    FD1S3AX b1_reg_i5 (.D(b_c_5), .CK(clk_c), .Q(b1_reg[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i5.GSR = "ENABLED";
    IB d_pad_10 (.I(d[10]), .O(d_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_15 (.I(d[15]), .O(d_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB d_pad_14 (.I(d[14]), .O(d_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    FD1S3AX b1_reg_i4 (.D(b_c_4), .CK(clk_c), .Q(b1_reg[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i4.GSR = "ENABLED";
    IB d_pad_13 (.I(d[13]), .O(d_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[35:36])
    IB c_pad_10 (.I(c[10]), .O(c_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_9 (.I(c[9]), .O(c_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_0 (.I(c[0]), .O(c_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    FD1S3AX b1_reg_i3 (.D(b_c_3), .CK(clk_c), .Q(b1_reg[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i3.GSR = "ENABLED";
    IB c_pad_1 (.I(c[1]), .O(c_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_6 (.I(c[6]), .O(c_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_5 (.I(c[5]), .O(c_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    FD1S3AX b1_reg_i2 (.D(b_c_2), .CK(clk_c), .Q(b1_reg[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i2.GSR = "ENABLED";
    IB c_pad_4 (.I(c[4]), .O(c_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_15 (.I(c[15]), .O(c_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_14 (.I(c[14]), .O(c_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_7 (.I(c[7]), .O(c_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    FD1S3AX b1_reg_i1 (.D(b_c_1), .CK(clk_c), .Q(b1_reg[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam b1_reg_i1.GSR = "ENABLED";
    IB c_pad_8 (.I(c[8]), .O(c_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_13 (.I(c[13]), .O(c_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    IB c_pad_12 (.I(c[12]), .O(c_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    FD1S3AX a1_reg_i15 (.D(a_c_15), .CK(clk_c), .Q(a1_reg[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i15.GSR = "ENABLED";
    IB c_pad_11 (.I(c[11]), .O(c_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[32:33])
    OB b_inv_pad_12 (.I(b_inv_c_12), .O(b_inv[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_13 (.I(b_inv_c_13), .O(b_inv[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB a_inv_pad_10 (.I(a_inv_c_10), .O(a_inv[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    FD1S3AX a1_reg_i14 (.D(a_c_14), .CK(clk_c), .Q(a1_reg[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i14.GSR = "ENABLED";
    OB a_inv_pad_9 (.I(a_inv_c_9), .O(a_inv[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB b_inv_pad_14 (.I(b_inv_c_14), .O(b_inv[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB b_inv_pad_15 (.I(b_inv_c_15), .O(b_inv[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    FD1S3AX a1_reg_i13 (.D(a_c_13), .CK(clk_c), .Q(a1_reg[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i13.GSR = "ENABLED";
    OB a_inv_pad_1 (.I(a_inv_c_1), .O(a_inv[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    IB b_pad_15 (.I(b[15]), .O(b_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_14 (.I(b[14]), .O(b_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_5 (.I(b[5]), .O(b_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    FD1S3AX a1_reg_i12 (.D(a_c_12), .CK(clk_c), .Q(a1_reg[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i12.GSR = "ENABLED";
    IB b_pad_6 (.I(b[6]), .O(b_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_11 (.I(b[11]), .O(b_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_10 (.I(b[10]), .O(b_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    FD1S3AX a1_reg_i11 (.D(a_c_11), .CK(clk_c), .Q(a1_reg[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i11.GSR = "ENABLED";
    IB b_pad_9 (.I(b[9]), .O(b_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB a_pad_6 (.I(a[6]), .O(a_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_5 (.I(a[5]), .O(a_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB b_pad_12 (.I(b[12]), .O(b_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    FD1S3AX a1_reg_i10 (.D(a_c_10), .CK(clk_c), .Q(a1_reg[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i10.GSR = "ENABLED";
    IB b_pad_13 (.I(b[13]), .O(b_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB a_pad_2 (.I(a[2]), .O(a_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_1 (.I(a[1]), .O(a_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    FD1S3AX a1_reg_i9 (.D(a_c_9), .CK(clk_c), .Q(a1_reg[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i9.GSR = "ENABLED";
    IB a_pad_0 (.I(a[0]), .O(a_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_13 (.I(a[13]), .O(a_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_12 (.I(a[12]), .O(a_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_3 (.I(a[3]), .O(a_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    FD1S3AX a1_reg_i8 (.D(a_c_8), .CK(clk_c), .Q(a1_reg[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i8.GSR = "ENABLED";
    IB a_pad_4 (.I(a[4]), .O(a_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_9 (.I(a[9]), .O(a_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB a_pad_8 (.I(a[8]), .O(a_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    FD1S3AX a1_reg_i7 (.D(a_c_7), .CK(clk_c), .Q(a1_reg[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i7.GSR = "ENABLED";
    IB a_pad_7 (.I(a[7]), .O(a_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    OB d_inv_pad_1 (.I(d_inv_c_1), .O(d_inv[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_0 (.I(d_inv_c_0), .O(d_inv[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    IB a_pad_10 (.I(a[10]), .O(a_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    FD1S3AX a1_reg_i6 (.D(a_c_6), .CK(clk_c), .Q(a1_reg[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i6.GSR = "ENABLED";
    IB a_pad_11 (.I(a[11]), .O(a_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    IB reset_pad (.I(reset), .O(reset_c));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[25:30])
    IB a_pad_15 (.I(a[15]), .O(a_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    FD1S3AX a1_reg_i5 (.D(a_c_5), .CK(clk_c), .Q(a1_reg[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i5.GSR = "ENABLED";
    IB a_pad_14 (.I(a[14]), .O(a_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[26:27])
    OB d_inv_pad_8 (.I(d_inv_c_8), .O(d_inv[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_7 (.I(d_inv_c_7), .O(d_inv[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[20:23])
    FD1S3AX a1_reg_i4 (.D(a_c_4), .CK(clk_c), .Q(a1_reg[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i4.GSR = "ENABLED";
    OB error_pad (.I(error_c), .O(error));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(19[26:31])
    OB d_inv_pad_4 (.I(d_inv_c_4), .O(d_inv[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_3 (.I(d_inv_c_3), .O(d_inv[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    FD1S3AX a1_reg_i3 (.D(a_c_3), .CK(clk_c), .Q(a1_reg[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i3.GSR = "ENABLED";
    OB d_inv_pad_2 (.I(d_inv_c_2), .O(d_inv[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_15 (.I(d_inv_c_15), .O(d_inv[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_14 (.I(d_inv_c_14), .O(d_inv[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_5 (.I(d_inv_c_5), .O(d_inv[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    FD1S3AX a1_reg_i2 (.D(a_c_2), .CK(clk_c), .Q(a1_reg[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i2.GSR = "ENABLED";
    OB d_inv_pad_6 (.I(d_inv_c_6), .O(d_inv[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_11 (.I(d_inv_c_11), .O(d_inv[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB d_inv_pad_10 (.I(d_inv_c_10), .O(d_inv[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    FD1S3AX a1_reg_i1 (.D(a_c_1), .CK(clk_c), .Q(a1_reg[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i1.GSR = "ENABLED";
    OB d_inv_pad_9 (.I(d_inv_c_9), .O(d_inv[9]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB c_inv_pad_6 (.I(c_inv_c_6), .O(c_inv[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_5 (.I(c_inv_c_5), .O(c_inv[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB d_inv_pad_12 (.I(d_inv_c_12), .O(d_inv[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    FD1S3AX a1_reg_i0 (.D(a_c_0), .CK(clk_c), .Q(a1_reg[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam a1_reg_i0.GSR = "ENABLED";
    OB d_inv_pad_13 (.I(d_inv_c_13), .O(d_inv[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[47:52])
    OB c_inv_pad_4 (.I(c_inv_c_4), .O(c_inv[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_1 (.I(c_inv_c_1), .O(c_inv[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    FD1S3AX b_inv_reg_res2_i2 (.D(b_inv_15__N_17[33]), .CK(clk_c), .Q(b_inv_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i2.GSR = "ENABLED";
    OB c_inv_pad_0 (.I(c_inv_c_0), .O(c_inv[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_15 (.I(c_inv_c_15), .O(c_inv[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_14 (.I(c_inv_c_14), .O(c_inv[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_2 (.I(c_inv_c_2), .O(c_inv[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB a_inv_pad_15 (.I(a_inv_c_15), .O(a_inv[15]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    OB c_inv_pad_3 (.I(c_inv_c_3), .O(c_inv[3]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_13 (.I(c_inv_c_13), .O(c_inv[13]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_12 (.I(c_inv_c_12), .O(c_inv[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    GSR GSR_INST (.GSR(n11713));
    OB b_inv_pad_0 (.I(b_inv_c_0), .O(b_inv[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB c_inv_pad_11 (.I(c_inv_c_11), .O(c_inv[11]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB c_inv_pad_10 (.I(c_inv_c_10), .O(c_inv[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB b_inv_pad_1 (.I(b_inv_c_1), .O(b_inv[1]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[33:38])
    OB c_inv_pad_7 (.I(c_inv_c_7), .O(c_inv[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[40:45])
    OB a_inv_pad_7 (.I(a_inv_c_7), .O(a_inv[7]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(18[26:31])
    LUT4 i1498_2_lut_4_lut (.A(n68_adj_538), .B(n68_adj_506), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n60)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1498_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_334_i1_3_lut_rep_77 (.A(n68_adj_1620), .B(n68_adj_2098), .C(n2650), 
         .Z(n13827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_334_i1_3_lut_rep_77.init = 16'hcaca;
    LUT4 mux_342_i1_3_lut_rep_69 (.A(n68_adj_538), .B(n68_adj_506), .C(n2650), 
         .Z(n13819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_342_i1_3_lut_rep_69.init = 16'hcaca;
    LUT4 i1486_4_lut (.A(n57_adj_2196), .B(n62_adj_2194), .C(n51_adj_2200), 
         .D(n52_adj_2199), .Z(det_zero_reg_N_162)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i1486_4_lut.init = 16'h0001;
    IB b_pad_0 (.I(b[0]), .O(b_c_0));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_1 (.I(b[1]), .O(b_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_2 (.I(b[2]), .O(b_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_3 (.I(b[3]), .O(b_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    IB b_pad_4 (.I(b[4]), .O(b_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(17[29:30])
    LUT4 i25_4_lut (.A(det_q4_28_31__N_65[0]), .B(n50_adj_2201), .C(n34_adj_2205), 
         .D(det_q4_28_31__N_65[27]), .Z(n57_adj_2196)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41_adj_2204), .B(n60_adj_2195), .C(n54_adj_2198), 
         .D(n42_adj_2203), .Z(n62_adj_2194)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(det_q4_28_31__N_65[3]), .B(det_q4_28_31__N_65[5]), 
         .C(det_q4_28_31__N_65[15]), .D(det_q4_28_31__N_65[7]), .Z(n51_adj_2200)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i20_4_lut (.A(det_q4_28_31__N_65[1]), .B(det_q4_28_31__N_65[21]), 
         .C(det_q4_28_31__N_65[11]), .D(det_q4_28_31__N_65[16]), .Z(n52_adj_2199)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(det_q4_28_31__N_65[29]), .B(det_q4_28_31__N_65[17]), 
         .C(det_q4_28_31__N_65[19]), .D(det_q4_28_31__N_65[8]), .Z(n50_adj_2201)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(det_q4_28_31__N_65[10]), .B(det_q4_28_31__N_65[25]), 
         .Z(n34_adj_2205)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i9_2_lut (.A(det_q4_28_31__N_65[9]), .B(det_q4_28_31__N_65[26]), 
         .Z(n41_adj_2204)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(n55_adj_2197), .B(det_q4_28_31__N_65[30]), .C(n48_adj_2202), 
         .D(det_q4_28_31__N_65[4]), .Z(n60_adj_2195)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(det_q4_28_31__N_65[28]), .B(det_q4_28_31__N_65[13]), 
         .C(det_q4_28_31__N_65[31]), .D(det_q4_28_31__N_65[23]), .Z(n54_adj_2198)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(det_q4_28_31__N_65[18]), .B(det_q4_28_31__N_65[2]), 
         .Z(n42_adj_2203)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(det_q4_28_31__N_65[20]), .B(det_q4_28_31__N_65[22]), 
         .C(det_q4_28_31__N_65[6]), .D(det_q4_28_31__N_65[14]), .Z(n55_adj_2197)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i16_2_lut (.A(det_q4_28_31__N_65[24]), .B(det_q4_28_31__N_65[12]), 
         .Z(n48_adj_2202)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(60[29:53])
    defparam i16_2_lut.init = 16'heeee;
    LUT4 i1522_2_lut_4_lut (.A(n68_adj_1620), .B(n68_adj_2098), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n52)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1522_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_333_i1_3_lut_rep_78 (.A(n68_adj_1940), .B(n68_adj_1749), .C(n2650), 
         .Z(n13828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_333_i1_3_lut_rep_78.init = 16'hcaca;
    LUT4 i1525_2_lut_4_lut (.A(n68_adj_1940), .B(n68_adj_1749), .C(n2650), 
         .D(inv_det_31__N_227), .Z(n51)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1525_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_320_i1_3_lut_rep_79 (.A(n68_adj_1588), .B(n68_adj_1556), .C(n1846), 
         .Z(n13829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_320_i1_3_lut_rep_79.init = 16'hcaca;
    LUT4 i1543_2_lut_4_lut (.A(n68_adj_1588), .B(n68_adj_1556), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n45)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1543_2_lut_4_lut.init = 16'h0035;
    LUT4 i696_2_lut_4_lut (.A(n68_adj_1588), .B(n68_adj_1556), .C(n1846), 
         .D(n1444), .Z(n2349)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i696_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_321_i1_3_lut_rep_80 (.A(n68_adj_1780), .B(n68_adj_794), .C(n1846), 
         .Z(n13830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_321_i1_3_lut_rep_80.init = 16'hcaca;
    LUT4 i1546_2_lut_4_lut (.A(n68_adj_1780), .B(n68_adj_794), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n44)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1546_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_322_i1_3_lut_rep_81 (.A(n68_adj_251), .B(n68_adj_1876), .C(n1846), 
         .Z(n13831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_322_i1_3_lut_rep_81.init = 16'hcaca;
    LUT4 i1549_2_lut_4_lut (.A(n68_adj_251), .B(n68_adj_1876), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n43)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1549_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_323_i1_3_lut_rep_82 (.A(n68_adj_1812), .B(n68_adj_1653), .C(n1846), 
         .Z(n13832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_323_i1_3_lut_rep_82.init = 16'hcaca;
    LUT4 i686_1_lut (.A(reset_c), .Z(n11713)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[25:30])
    defparam i686_1_lut.init = 16'h5555;
    LUT4 i1340_2_lut (.A(det_q4_28[1]), .B(det_q4_28[0]), .Z(n161_adj_1272)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1340_2_lut.init = 16'h6666;
    FD1S3AX b_inv_reg_res2_i3 (.D(b_inv_15__N_17[34]), .CK(clk_c), .Q(b_inv_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i3.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i4 (.D(b_inv_15__N_17[35]), .CK(clk_c), .Q(b_inv_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i4.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i5 (.D(b_inv_15__N_17[36]), .CK(clk_c), .Q(b_inv_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i5.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i6 (.D(b_inv_15__N_17[37]), .CK(clk_c), .Q(b_inv_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i6.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i7 (.D(b_inv_15__N_17[38]), .CK(clk_c), .Q(b_inv_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i7.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i8 (.D(b_inv_15__N_17[39]), .CK(clk_c), .Q(b_inv_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i8.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i9 (.D(b_inv_15__N_17[40]), .CK(clk_c), .Q(b_inv_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i9.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i10 (.D(b_inv_15__N_17[41]), .CK(clk_c), .Q(b_inv_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i10.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i11 (.D(b_inv_15__N_17[42]), .CK(clk_c), .Q(b_inv_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i11.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i12 (.D(b_inv_15__N_17[43]), .CK(clk_c), .Q(b_inv_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i12.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i13 (.D(b_inv_15__N_17[44]), .CK(clk_c), .Q(b_inv_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i13.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i14 (.D(b_inv_15__N_17[45]), .CK(clk_c), .Q(b_inv_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i14.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i15 (.D(b_inv_15__N_17[46]), .CK(clk_c), .Q(b_inv_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i15.GSR = "ENABLED";
    FD1S3AX b_inv_reg_res2_i16 (.D(b_inv_15__N_17[47]), .CK(clk_c), .Q(b_inv_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam b_inv_reg_res2_i16.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i2 (.D(c_inv_15__N_33[33]), .CK(clk_c), .Q(c_inv_c_1));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i2.GSR = "ENABLED";
    LUT4 i1552_2_lut_4_lut (.A(n68_adj_1812), .B(n68_adj_1653), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n42)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1552_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_324_i1_3_lut_rep_83 (.A(n68_adj_2162), .B(n68_adj_2066), .C(n1846), 
         .Z(n13833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_324_i1_3_lut_rep_83.init = 16'hcaca;
    LUT4 i1555_2_lut_4_lut (.A(n68_adj_2162), .B(n68_adj_2066), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n41)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1555_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_325_i1_3_lut_rep_84 (.A(n68_adj_1398), .B(n68_adj_1430), .C(n1846), 
         .Z(n13834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_325_i1_3_lut_rep_84.init = 16'hcaca;
    LUT4 i1558_2_lut_4_lut (.A(n68_adj_1398), .B(n68_adj_1430), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n40)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1558_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_326_i1_3_lut_rep_85 (.A(n68_adj_1335), .B(n68_adj_1367), .C(n1846), 
         .Z(n13835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_326_i1_3_lut_rep_85.init = 16'hcaca;
    LUT4 i1561_2_lut_4_lut (.A(n68_adj_1335), .B(n68_adj_1367), .C(n1846), 
         .D(inv_det_31__N_227), .Z(n39)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1561_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_332_i1_3_lut_rep_86 (.A(n68_adj_890), .B(n68_adj_858), .C(n1410), 
         .Z(n13836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_332_i1_3_lut_rep_86.init = 16'hcaca;
    LUT4 i1567_2_lut_4_lut (.A(n68_adj_890), .B(n68_adj_858), .C(n1410), 
         .D(inv_det_31__N_227), .Z(n37)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1567_2_lut_4_lut.init = 16'h0035;
    LUT4 i714_2_lut_4_lut (.A(n68_adj_890), .B(n68_adj_858), .C(n1410), 
         .D(n1444), .Z(n1813)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i714_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_331_i1_3_lut_rep_87 (.A(n68_adj_954), .B(n68_adj_922), .C(n1410), 
         .Z(n13837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_331_i1_3_lut_rep_87.init = 16'hcaca;
    LUT4 i1570_2_lut_4_lut (.A(n68_adj_954), .B(n68_adj_922), .C(n1410), 
         .D(inv_det_31__N_227), .Z(n36)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1570_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_330_i1_3_lut_rep_88 (.A(n68_adj_1018), .B(n68_adj_986), .C(n1410), 
         .Z(n13838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_330_i1_3_lut_rep_88.init = 16'hcaca;
    CCU2C _add_1_add_4_7 (.A0(n149_adj_1521), .B0(n2583), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1520), .B1(n2583), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12596), .COUT(n12597), .S0(n146_adj_373), 
          .S1(n143_adj_372));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_5 (.A0(n155_adj_1523), .B0(n2583), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1522), .B1(n2583), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12595), .COUT(n12596), .S0(n152_adj_375), 
          .S1(n149_adj_374));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_3 (.A0(n161_adj_1272), .B0(n2583), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1524), .B1(n2583), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12594), .COUT(n12595), .S0(n158_adj_377), 
          .S1(n155_adj_376));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(det_q4_28[0]), .B1(n2583), .C1(det_q4_28[1]), .D1(n1475), 
          .COUT(n12594), .S1(n161_adj_378));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_33 (.A0(n74_adj_1526), .B0(n2516), .C0(n71_adj_348), 
          .D0(n2618), .A1(n71_adj_1525), .B1(n2516), .C1(n68_adj_347), 
          .D1(n2617), .CIN(n12592), .S0(n71), .S1(n2650));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_33.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_33.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_31 (.A0(n80_adj_1528), .B0(n2516), .C0(n77_adj_350), 
          .D0(n2620), .A1(n77_adj_1527), .B1(n2516), .C1(n74_adj_349), 
          .D1(n2619), .CIN(n12591), .COUT(n12592), .S0(n77), .S1(n74));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_29 (.A0(n86_adj_1530), .B0(n2516), .C0(n83_adj_352), 
          .D0(n2622), .A1(n83_adj_1529), .B1(n2516), .C1(n80_adj_351), 
          .D1(n2621), .CIN(n12590), .COUT(n12591), .S0(n83), .S1(n80));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_27 (.A0(n92_adj_1532), .B0(n2516), .C0(n89_adj_354), 
          .D0(n2624), .A1(n89_adj_1531), .B1(n2516), .C1(n86_adj_353), 
          .D1(n2623), .CIN(n12589), .COUT(n12590), .S0(n89), .S1(n86));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_25 (.A0(n98_adj_1534), .B0(n2516), .C0(n95_adj_356), 
          .D0(n2626), .A1(n95_adj_1533), .B1(n2516), .C1(n92_adj_355), 
          .D1(n2625), .CIN(n12588), .COUT(n12589), .S0(n95), .S1(n92));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_23 (.A0(n104_adj_1536), .B0(n2516), .C0(n101_adj_358), 
          .D0(n2628), .A1(n101_adj_1535), .B1(n2516), .C1(n98_adj_357), 
          .D1(n2627), .CIN(n12587), .COUT(n12588), .S0(n101), .S1(n98));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_21 (.A0(n110_adj_1538), .B0(n2516), .C0(n107_adj_360), 
          .D0(n2630), .A1(n107_adj_1537), .B1(n2516), .C1(n104_adj_359), 
          .D1(n2629), .CIN(n12586), .COUT(n12587), .S0(n107), .S1(n104_adj_246));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_19 (.A0(n116_adj_1540), .B0(n2516), .C0(n113_adj_362), 
          .D0(n2632), .A1(n113_adj_1539), .B1(n2516), .C1(n110_adj_361), 
          .D1(n2631), .CIN(n12585), .COUT(n12586), .S0(n113), .S1(n110_adj_247));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_17 (.A0(n122_adj_1542), .B0(n2516), .C0(n119_adj_364), 
          .D0(n2634), .A1(n119_adj_1541), .B1(n2516), .C1(n116_adj_363), 
          .D1(n2633), .CIN(n12584), .COUT(n12585), .S0(n119), .S1(n116_adj_248));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_15 (.A0(n128_adj_1544), .B0(n2516), .C0(n125_adj_366), 
          .D0(n2636), .A1(n125_adj_1543), .B1(n2516), .C1(n122_adj_365), 
          .D1(n2635), .CIN(n12583), .COUT(n12584), .S0(n125), .S1(n122_adj_249));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_13 (.A0(n134_adj_1546), .B0(n2516), .C0(n131_adj_368), 
          .D0(n2638), .A1(n131_adj_1545), .B1(n2516), .C1(n128_adj_367), 
          .D1(n2637), .CIN(n12582), .COUT(n12583), .S0(n131), .S1(n128_adj_250));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_11 (.A0(n140_adj_1548), .B0(n2516), .C0(n137_adj_370), 
          .D0(n2640), .A1(n137_adj_1547), .B1(n2516), .C1(n134_adj_369), 
          .D1(n2639), .CIN(n12581), .COUT(n12582), .S0(n137), .S1(n134));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_9 (.A0(n146_adj_1550), .B0(n2516), .C0(n143_adj_372), 
          .D0(n2642), .A1(n143_adj_1549), .B1(n2516), .C1(n140_adj_371), 
          .D1(n2641), .CIN(n12580), .COUT(n12581), .S0(n143), .S1(n140));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_7 (.A0(n152_adj_1552), .B0(n2516), .C0(n149_adj_374), 
          .D0(n2644), .A1(n149_adj_1551), .B1(n2516), .C1(n146_adj_373), 
          .D1(n2643), .CIN(n12579), .COUT(n12580), .S0(n149), .S1(n146));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_5 (.A0(n158_adj_1554), .B0(n2516), .C0(n155_adj_376), 
          .D0(n2646), .A1(n155_adj_1553), .B1(n2516), .C1(n152_adj_375), 
          .D1(n2645), .CIN(n12578), .COUT(n12579), .S0(n155), .S1(n152));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_565_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_3 (.A0(det_q4_28[0]), .B0(n2516), .C0(n161_adj_378), 
          .D0(n2648), .A1(n161_adj_1555), .B1(n2516), .C1(n158_adj_377), 
          .D1(n2647), .CIN(n12577), .COUT(n12578), .S0(n161), .S1(n158));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_565_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_565_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_565_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2516), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12577));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_565_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_565_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_565_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_565_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_33 (.A0(n1444), .B0(n13832), .C0(n71_adj_1813), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12573), .S0(n68_adj_251));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_394_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_394_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_31 (.A0(n77_adj_1815), .B0(n13832), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1814), .B1(n13832), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12572), .COUT(n12573), .S0(n74_adj_253), 
          .S1(n71_adj_252));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_29 (.A0(n83_adj_1817), .B0(n13832), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1816), .B1(n13832), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12571), .COUT(n12572), .S0(n80_adj_255), 
          .S1(n77_adj_254));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_27 (.A0(n89_adj_1819), .B0(n13832), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1818), .B1(n13832), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12570), .COUT(n12571), .S0(n86_adj_257), 
          .S1(n83_adj_256));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_25 (.A0(n95_adj_1821), .B0(n13832), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1820), .B1(n13832), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12569), .COUT(n12570), .S0(n92_adj_259), 
          .S1(n89_adj_258));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_23 (.A0(n101_adj_1823), .B0(n13832), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1822), .B1(n13832), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12568), .COUT(n12569), .S0(n98_adj_261), 
          .S1(n95_adj_260));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_21 (.A0(n107_adj_1825), .B0(n13832), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1824), .B1(n13832), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12567), .COUT(n12568), .S0(n104_adj_263), 
          .S1(n101_adj_262));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_19 (.A0(n113_adj_1827), .B0(n13832), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1826), .B1(n13832), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12566), .COUT(n12567), .S0(n110_adj_265), 
          .S1(n107_adj_264));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_17 (.A0(n119_adj_1829), .B0(n13832), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1828), .B1(n13832), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12565), .COUT(n12566), .S0(n116_adj_267), 
          .S1(n113_adj_266));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_15 (.A0(n125_adj_1831), .B0(n13832), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1830), .B1(n13832), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12564), .COUT(n12565), .S0(n122_adj_269), 
          .S1(n119_adj_268));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_13 (.A0(n131_adj_1833), .B0(n13832), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1832), .B1(n13832), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12563), .COUT(n12564), .S0(n128_adj_271), 
          .S1(n125_adj_270));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_11 (.A0(n137_adj_1835), .B0(n13832), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1834), .B1(n13832), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12562), .COUT(n12563), .S0(n134_adj_273), 
          .S1(n131_adj_272));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_9 (.A0(n143_adj_1837), .B0(n13832), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1836), .B1(n13832), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12561), .COUT(n12562), .S0(n140_adj_275), 
          .S1(n137_adj_274));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_7 (.A0(n149_adj_1839), .B0(n13832), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1838), .B1(n13832), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12560), .COUT(n12561), .S0(n146_adj_277), 
          .S1(n143_adj_276));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_5 (.A0(n155_adj_1841), .B0(n13832), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1840), .B1(n13832), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12559), .COUT(n12560), .S0(n152_adj_279), 
          .S1(n149_adj_278));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_3 (.A0(n161_adj_1843), .B0(n13832), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1842), .B1(n13832), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12558), .COUT(n12559), .S0(n158_adj_281), 
          .S1(n155_adj_280));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_394_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_394_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13832), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12558), .S1(n161_adj_282));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_394_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_394_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_394_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_394_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_33 (.A0(n1444), .B0(n3454), .C0(n71_adj_380), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12557), .S0(n68_adj_283));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_562_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_562_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_31 (.A0(n77_adj_382), .B0(n3454), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_381), .B1(n3454), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12556), .COUT(n12557), .S0(n74_adj_285), 
          .S1(n71_adj_284));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_29 (.A0(n83_adj_384), .B0(n3454), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_383), .B1(n3454), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12555), .COUT(n12556), .S0(n80_adj_287), 
          .S1(n77_adj_286));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_27 (.A0(n89_adj_386), .B0(n3454), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_385), .B1(n3454), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12554), .COUT(n12555), .S0(n86_adj_289), 
          .S1(n83_adj_288));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_25 (.A0(n95_adj_388), .B0(n3454), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_387), .B1(n3454), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12553), .COUT(n12554), .S0(n92_adj_291), 
          .S1(n89_adj_290));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_23 (.A0(n101_adj_390), .B0(n3454), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_389), .B1(n3454), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12552), .COUT(n12553), .S0(n98_adj_293), 
          .S1(n95_adj_292));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_21 (.A0(n107_adj_392), .B0(n3454), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_391), .B1(n3454), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12551), .COUT(n12552), .S0(n104_adj_295), 
          .S1(n101_adj_294));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_19 (.A0(n113_adj_394), .B0(n3454), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_393), .B1(n3454), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12550), .COUT(n12551), .S0(n110_adj_297), 
          .S1(n107_adj_296));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_17 (.A0(n119_adj_396), .B0(n3454), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_395), .B1(n3454), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12549), .COUT(n12550), .S0(n116_adj_299), 
          .S1(n113_adj_298));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_15 (.A0(n125_adj_398), .B0(n3454), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_397), .B1(n3454), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12548), .COUT(n12549), .S0(n122_adj_301), 
          .S1(n119_adj_300));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_13 (.A0(n131_adj_400), .B0(n3454), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_399), .B1(n3454), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12547), .COUT(n12548), .S0(n128_adj_303), 
          .S1(n125_adj_302));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_11 (.A0(n137_adj_402), .B0(n3454), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_401), .B1(n3454), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12546), .COUT(n12547), .S0(n134_adj_305), 
          .S1(n131_adj_304));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_9 (.A0(n143_adj_404), .B0(n3454), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_403), .B1(n3454), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12545), .COUT(n12546), .S0(n140_adj_307), 
          .S1(n137_adj_306));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_7 (.A0(n149_adj_406), .B0(n3454), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_405), .B1(n3454), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12544), .COUT(n12545), .S0(n146_adj_309), 
          .S1(n143_adj_308));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_5 (.A0(n155_adj_408), .B0(n3454), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_407), .B1(n3454), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12543), .COUT(n12544), .S0(n152_adj_311), 
          .S1(n149_adj_310));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_3 (.A0(n161_adj_410), .B0(n3454), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_409), .B1(n3454), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12542), .COUT(n12543), .S0(n158_adj_313), 
          .S1(n155_adj_312));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_562_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_562_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n3454), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12542), .S1(n161_adj_314));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_562_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_562_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_562_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_562_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_33 (.A0(n1444), .B0(n13818), .C0(n71_adj_443), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12541), .S0(n68_adj_379));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_556_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_556_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_31 (.A0(n77_adj_445), .B0(n13818), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_444), .B1(n13818), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12540), .COUT(n12541), .S0(n74_adj_381), 
          .S1(n71_adj_380));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_29 (.A0(n83_adj_447), .B0(n13818), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_446), .B1(n13818), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12539), .COUT(n12540), .S0(n80_adj_383), 
          .S1(n77_adj_382));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_27 (.A0(n89_adj_449), .B0(n13818), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_448), .B1(n13818), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12538), .COUT(n12539), .S0(n86_adj_385), 
          .S1(n83_adj_384));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_25 (.A0(n95_adj_451), .B0(n13818), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_450), .B1(n13818), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12537), .COUT(n12538), .S0(n92_adj_387), 
          .S1(n89_adj_386));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_23 (.A0(n101_adj_453), .B0(n13818), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_452), .B1(n13818), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12536), .COUT(n12537), .S0(n98_adj_389), 
          .S1(n95_adj_388));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_21 (.A0(n107_adj_455), .B0(n13818), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_454), .B1(n13818), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12535), .COUT(n12536), .S0(n104_adj_391), 
          .S1(n101_adj_390));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_19 (.A0(n113_adj_457), .B0(n13818), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_456), .B1(n13818), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12534), .COUT(n12535), .S0(n110_adj_393), 
          .S1(n107_adj_392));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_17 (.A0(n119_adj_459), .B0(n13818), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_458), .B1(n13818), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12533), .COUT(n12534), .S0(n116_adj_395), 
          .S1(n113_adj_394));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_15 (.A0(n125_adj_461), .B0(n13818), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_460), .B1(n13818), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12532), .COUT(n12533), .S0(n122_adj_397), 
          .S1(n119_adj_396));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_13 (.A0(n131_adj_463), .B0(n13818), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_462), .B1(n13818), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12531), .COUT(n12532), .S0(n128_adj_399), 
          .S1(n125_adj_398));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_11 (.A0(n137_adj_465), .B0(n13818), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_464), .B1(n13818), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12530), .COUT(n12531), .S0(n134_adj_401), 
          .S1(n131_adj_400));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_9 (.A0(n143_adj_467), .B0(n13818), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_466), .B1(n13818), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12529), .COUT(n12530), .S0(n140_adj_403), 
          .S1(n137_adj_402));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_7 (.A0(n149_adj_469), .B0(n13818), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_468), .B1(n13818), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12528), .COUT(n12529), .S0(n146_adj_405), 
          .S1(n143_adj_404));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_5 (.A0(n155_adj_471), .B0(n13818), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_470), .B1(n13818), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12527), .COUT(n12528), .S0(n152_adj_407), 
          .S1(n149_adj_406));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_3 (.A0(n161_adj_473), .B0(n13818), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_472), .B1(n13818), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12526), .COUT(n12527), .S0(n158_adj_409), 
          .S1(n155_adj_408));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_556_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_556_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13818), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12526), .S1(n161_adj_410));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_556_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_556_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_556_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_556_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_33 (.A0(n3422), .B0(n2650), .C0(n74_adj_476), 
          .D0(VCC_net), .A1(n71_adj_475), .B1(n2650), .C1(n68_adj_379), 
          .D1(n3421), .CIN(n12524), .S0(n71_adj_411), .S1(n3454));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_33.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_553_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_33.INJECT1_1 = "NO";
    FD1S3AX c_inv_reg_res1_i3 (.D(c_inv_15__N_33[34]), .CK(clk_c), .Q(c_inv_c_2));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i3.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i4 (.D(c_inv_15__N_33[35]), .CK(clk_c), .Q(c_inv_c_3));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i4.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i5 (.D(c_inv_15__N_33[36]), .CK(clk_c), .Q(c_inv_c_4));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i5.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i6 (.D(c_inv_15__N_33[37]), .CK(clk_c), .Q(c_inv_c_5));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i6.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i7 (.D(c_inv_15__N_33[38]), .CK(clk_c), .Q(c_inv_c_6));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i7.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i8 (.D(c_inv_15__N_33[39]), .CK(clk_c), .Q(c_inv_c_7));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i8.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i9 (.D(c_inv_15__N_33[40]), .CK(clk_c), .Q(c_inv_c_8));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i9.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i10 (.D(c_inv_15__N_33[41]), .CK(clk_c), .Q(c_inv_c_9));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i10.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i11 (.D(c_inv_15__N_33[42]), .CK(clk_c), .Q(c_inv_c_10));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i11.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i12 (.D(c_inv_15__N_33[43]), .CK(clk_c), .Q(c_inv_c_11));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i12.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i13 (.D(c_inv_15__N_33[44]), .CK(clk_c), .Q(c_inv_c_12));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i13.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i14 (.D(c_inv_15__N_33[45]), .CK(clk_c), .Q(c_inv_c_13));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i14.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i15 (.D(c_inv_15__N_33[46]), .CK(clk_c), .Q(c_inv_c_14));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i15.GSR = "ENABLED";
    FD1S3AX c_inv_reg_res1_i16 (.D(c_inv_15__N_33[47]), .CK(clk_c), .Q(c_inv_c_15));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(129[18] 135[12])
    defparam c_inv_reg_res1_i16.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i2 (.D(d1_reg[1]), .CK(clk_c), .Q(n128_adj_232));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i2.GSR = "ENABLED";
    CCU2C _add_1_553_add_4_31 (.A0(n3424), .B0(n2650), .C0(n80_adj_478), 
          .D0(VCC_net), .A1(n3423), .B1(n2650), .C1(n77_adj_477), .D1(VCC_net), 
          .CIN(n12523), .COUT(n12524), .S0(n77_adj_413), .S1(n74_adj_412));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_31.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_31.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_29 (.A0(n3426), .B0(n2650), .C0(n86_adj_480), 
          .D0(VCC_net), .A1(n3425), .B1(n2650), .C1(n83_adj_479), .D1(VCC_net), 
          .CIN(n12522), .COUT(n12523), .S0(n83_adj_415), .S1(n80_adj_414));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_29.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_29.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_27 (.A0(n3428), .B0(n2650), .C0(n92_adj_482), 
          .D0(VCC_net), .A1(n3427), .B1(n2650), .C1(n89_adj_481), .D1(VCC_net), 
          .CIN(n12521), .COUT(n12522), .S0(n89_adj_417), .S1(n86_adj_416));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_27.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_27.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_25 (.A0(n3430), .B0(n2650), .C0(n98_adj_484), 
          .D0(VCC_net), .A1(n3429), .B1(n2650), .C1(n95_adj_483), .D1(VCC_net), 
          .CIN(n12520), .COUT(n12521), .S0(n95_adj_419), .S1(n92_adj_418));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_25.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_25.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_23 (.A0(n3432), .B0(n2650), .C0(n104_adj_486), 
          .D0(VCC_net), .A1(n3431), .B1(n2650), .C1(n101_adj_485), .D1(VCC_net), 
          .CIN(n12519), .COUT(n12520), .S0(n101_adj_421), .S1(n98_adj_420));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_23.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_23.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_21 (.A0(n3434), .B0(n2650), .C0(n110_adj_488), 
          .D0(VCC_net), .A1(n3433), .B1(n2650), .C1(n107_adj_487), .D1(VCC_net), 
          .CIN(n12518), .COUT(n12519), .S0(n107_adj_423), .S1(n104_adj_422));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_21.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_21.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_19 (.A0(n3436), .B0(n2650), .C0(n116_adj_490), 
          .D0(VCC_net), .A1(n3435), .B1(n2650), .C1(n113_adj_489), .D1(VCC_net), 
          .CIN(n12517), .COUT(n12518), .S0(n113_adj_425), .S1(n110_adj_424));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_19.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_19.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_17 (.A0(n3438), .B0(n2650), .C0(n122_adj_492), 
          .D0(VCC_net), .A1(n3437), .B1(n2650), .C1(n119_adj_491), .D1(VCC_net), 
          .CIN(n12516), .COUT(n12517), .S0(n119_adj_427), .S1(n116_adj_426));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_17.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_17.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_15 (.A0(n3440), .B0(n2650), .C0(n128_adj_494), 
          .D0(VCC_net), .A1(n3439), .B1(n2650), .C1(n125_adj_493), .D1(VCC_net), 
          .CIN(n12515), .COUT(n12516), .S0(n125_adj_429), .S1(n122_adj_428));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_15.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_15.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_13 (.A0(n3442), .B0(n2650), .C0(n134_adj_496), 
          .D0(VCC_net), .A1(n3441), .B1(n2650), .C1(n131_adj_495), .D1(VCC_net), 
          .CIN(n12514), .COUT(n12515), .S0(n131_adj_431), .S1(n128_adj_430));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_13.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_13.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_11 (.A0(n3444), .B0(n2650), .C0(n140_adj_498), 
          .D0(VCC_net), .A1(n3443), .B1(n2650), .C1(n137_adj_497), .D1(VCC_net), 
          .CIN(n12513), .COUT(n12514), .S0(n137_adj_433), .S1(n134_adj_432));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_11.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_11.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_9 (.A0(n3446), .B0(n2650), .C0(n146_adj_500), 
          .D0(VCC_net), .A1(n3445), .B1(n2650), .C1(n143_adj_499), .D1(VCC_net), 
          .CIN(n12512), .COUT(n12513), .S0(n143_adj_435), .S1(n140_adj_434));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_9.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_9.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_7 (.A0(n3448), .B0(n2650), .C0(n152_adj_502), 
          .D0(VCC_net), .A1(n3447), .B1(n2650), .C1(n149_adj_501), .D1(VCC_net), 
          .CIN(n12511), .COUT(n12512), .S0(n149_adj_437), .S1(n146_adj_436));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_7.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_7.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_5 (.A0(n3450), .B0(n2650), .C0(n158_adj_504), 
          .D0(VCC_net), .A1(n3449), .B1(n2650), .C1(n155_adj_503), .D1(VCC_net), 
          .CIN(n12510), .COUT(n12511), .S0(n155_adj_439), .S1(n152_adj_438));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_5.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_5.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_3 (.A0(n3452), .B0(n2650), .C0(det_q4_28[0]), 
          .D0(VCC_net), .A1(n3451), .B1(n2650), .C1(n161_adj_505), .D1(VCC_net), 
          .CIN(n12509), .COUT(n12510), .S0(n161_adj_441), .S1(n158_adj_440));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_3.INIT0 = 16'h1212;
    defparam _add_1_553_add_4_3.INIT1 = 16'h1212;
    defparam _add_1_553_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_553_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2650), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12509));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_553_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_553_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_553_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_553_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_33 (.A0(n1444), .B0(n13819), .C0(n71_adj_507), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12505), .S0(n68_adj_442));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_550_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_550_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_31 (.A0(n77_adj_509), .B0(n13819), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_508), .B1(n13819), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12504), .COUT(n12505), .S0(n74_adj_444), 
          .S1(n71_adj_443));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_29 (.A0(n83_adj_511), .B0(n13819), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_510), .B1(n13819), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12503), .COUT(n12504), .S0(n80_adj_446), 
          .S1(n77_adj_445));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_27 (.A0(n89_adj_513), .B0(n13819), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_512), .B1(n13819), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12502), .COUT(n12503), .S0(n86_adj_448), 
          .S1(n83_adj_447));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_25 (.A0(n95_adj_515), .B0(n13819), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_514), .B1(n13819), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12501), .COUT(n12502), .S0(n92_adj_450), 
          .S1(n89_adj_449));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_23 (.A0(n101_adj_517), .B0(n13819), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_516), .B1(n13819), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12500), .COUT(n12501), .S0(n98_adj_452), 
          .S1(n95_adj_451));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_21 (.A0(n107_adj_519), .B0(n13819), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_518), .B1(n13819), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12499), .COUT(n12500), .S0(n104_adj_454), 
          .S1(n101_adj_453));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_19 (.A0(n113_adj_521), .B0(n13819), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_520), .B1(n13819), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12498), .COUT(n12499), .S0(n110_adj_456), 
          .S1(n107_adj_455));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_17 (.A0(n119_adj_523), .B0(n13819), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_522), .B1(n13819), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12497), .COUT(n12498), .S0(n116_adj_458), 
          .S1(n113_adj_457));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_15 (.A0(n125_adj_525), .B0(n13819), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_524), .B1(n13819), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12496), .COUT(n12497), .S0(n122_adj_460), 
          .S1(n119_adj_459));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_13 (.A0(n131_adj_527), .B0(n13819), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_526), .B1(n13819), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12495), .COUT(n12496), .S0(n128_adj_462), 
          .S1(n125_adj_461));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_11 (.A0(n137_adj_529), .B0(n13819), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_528), .B1(n13819), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12494), .COUT(n12495), .S0(n134_adj_464), 
          .S1(n131_adj_463));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_9 (.A0(n143_adj_531), .B0(n13819), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_530), .B1(n13819), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12493), .COUT(n12494), .S0(n140_adj_466), 
          .S1(n137_adj_465));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_7 (.A0(n149_adj_533), .B0(n13819), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_532), .B1(n13819), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12492), .COUT(n12493), .S0(n146_adj_468), 
          .S1(n143_adj_467));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_5 (.A0(n155_adj_535), .B0(n13819), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_534), .B1(n13819), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12491), .COUT(n12492), .S0(n152_adj_470), 
          .S1(n149_adj_469));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_3 (.A0(n161_adj_537), .B0(n13819), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_536), .B1(n13819), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12490), .COUT(n12491), .S0(n158_adj_472), 
          .S1(n155_adj_471));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_550_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_550_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13819), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12490), .S1(n161_adj_473));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_550_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_550_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_550_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_550_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_33 (.A0(n1444), .B0(n13819), .C0(n71_adj_539), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12489), .S0(n68_adj_474));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_547_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_547_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_31 (.A0(n77_adj_541), .B0(n13819), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_540), .B1(n13819), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12488), .COUT(n12489), .S0(n74_adj_476), 
          .S1(n71_adj_475));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_29 (.A0(n83_adj_543), .B0(n13819), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_542), .B1(n13819), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12487), .COUT(n12488), .S0(n80_adj_478), 
          .S1(n77_adj_477));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_27 (.A0(n89_adj_545), .B0(n13819), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_544), .B1(n13819), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12486), .COUT(n12487), .S0(n86_adj_480), 
          .S1(n83_adj_479));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_25 (.A0(n95_adj_547), .B0(n13819), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_546), .B1(n13819), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12485), .COUT(n12486), .S0(n92_adj_482), 
          .S1(n89_adj_481));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_23 (.A0(n101_adj_549), .B0(n13819), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_548), .B1(n13819), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12484), .COUT(n12485), .S0(n98_adj_484), 
          .S1(n95_adj_483));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_21 (.A0(n107_adj_551), .B0(n13819), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_550), .B1(n13819), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12483), .COUT(n12484), .S0(n104_adj_486), 
          .S1(n101_adj_485));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_19 (.A0(n113_adj_553), .B0(n13819), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_552), .B1(n13819), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12482), .COUT(n12483), .S0(n110_adj_488), 
          .S1(n107_adj_487));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_17 (.A0(n119_adj_555), .B0(n13819), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_554), .B1(n13819), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12481), .COUT(n12482), .S0(n116_adj_490), 
          .S1(n113_adj_489));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_15 (.A0(n125_adj_557), .B0(n13819), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_556), .B1(n13819), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12480), .COUT(n12481), .S0(n122_adj_492), 
          .S1(n119_adj_491));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_13 (.A0(n131_adj_559), .B0(n13819), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_558), .B1(n13819), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12479), .COUT(n12480), .S0(n128_adj_494), 
          .S1(n125_adj_493));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_11 (.A0(n137_adj_561), .B0(n13819), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_560), .B1(n13819), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12478), .COUT(n12479), .S0(n134_adj_496), 
          .S1(n131_adj_495));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_9 (.A0(n143_adj_563), .B0(n13819), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_562), .B1(n13819), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12477), .COUT(n12478), .S0(n140_adj_498), 
          .S1(n137_adj_497));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_7 (.A0(n149_adj_565), .B0(n13819), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_564), .B1(n13819), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12476), .COUT(n12477), .S0(n146_adj_500), 
          .S1(n143_adj_499));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_5 (.A0(n155_adj_567), .B0(n13819), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_566), .B1(n13819), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12475), .COUT(n12476), .S0(n152_adj_502), 
          .S1(n149_adj_501));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_3 (.A0(n161_adj_569), .B0(n13819), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_568), .B1(n13819), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12474), .COUT(n12475), .S0(n158_adj_504), 
          .S1(n155_adj_503));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_547_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_547_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13819), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12474), .S1(n161_adj_505));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_547_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_547_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_547_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_547_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_33 (.A0(n1444), .B0(n13820), .C0(n71_adj_571), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12473), .S0(n68_adj_506));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_544_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_544_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_31 (.A0(n77_adj_573), .B0(n13820), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_572), .B1(n13820), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12472), .COUT(n12473), .S0(n74_adj_508), 
          .S1(n71_adj_507));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_29 (.A0(n83_adj_575), .B0(n13820), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_574), .B1(n13820), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12471), .COUT(n12472), .S0(n80_adj_510), 
          .S1(n77_adj_509));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_27 (.A0(n89_adj_577), .B0(n13820), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_576), .B1(n13820), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12470), .COUT(n12471), .S0(n86_adj_512), 
          .S1(n83_adj_511));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_25 (.A0(n95_adj_579), .B0(n13820), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_578), .B1(n13820), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12469), .COUT(n12470), .S0(n92_adj_514), 
          .S1(n89_adj_513));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_23 (.A0(n101_adj_581), .B0(n13820), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_580), .B1(n13820), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12468), .COUT(n12469), .S0(n98_adj_516), 
          .S1(n95_adj_515));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_21 (.A0(n107_adj_583), .B0(n13820), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_582), .B1(n13820), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12467), .COUT(n12468), .S0(n104_adj_518), 
          .S1(n101_adj_517));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_19 (.A0(n113_adj_585), .B0(n13820), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_584), .B1(n13820), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12466), .COUT(n12467), .S0(n110_adj_520), 
          .S1(n107_adj_519));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_17 (.A0(n119_adj_587), .B0(n13820), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_586), .B1(n13820), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12465), .COUT(n12466), .S0(n116_adj_522), 
          .S1(n113_adj_521));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_15 (.A0(n125_adj_589), .B0(n13820), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_588), .B1(n13820), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12464), .COUT(n12465), .S0(n122_adj_524), 
          .S1(n119_adj_523));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_13 (.A0(n131_adj_591), .B0(n13820), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_590), .B1(n13820), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12463), .COUT(n12464), .S0(n128_adj_526), 
          .S1(n125_adj_525));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_11 (.A0(n137_adj_593), .B0(n13820), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_592), .B1(n13820), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12462), .COUT(n12463), .S0(n134_adj_528), 
          .S1(n131_adj_527));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_9 (.A0(n143_adj_595), .B0(n13820), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_594), .B1(n13820), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12461), .COUT(n12462), .S0(n140_adj_530), 
          .S1(n137_adj_529));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_7 (.A0(n149_adj_597), .B0(n13820), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_596), .B1(n13820), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12460), .COUT(n12461), .S0(n146_adj_532), 
          .S1(n143_adj_531));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_5 (.A0(n155_adj_599), .B0(n13820), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_598), .B1(n13820), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12459), .COUT(n12460), .S0(n152_adj_534), 
          .S1(n149_adj_533));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_3 (.A0(n161_adj_601), .B0(n13820), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_600), .B1(n13820), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12458), .COUT(n12459), .S0(n158_adj_536), 
          .S1(n155_adj_535));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_544_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_544_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13820), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12458), .S1(n161_adj_537));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_544_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_544_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_544_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_544_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_33 (.A0(n1444), .B0(n13820), .C0(n71_adj_603), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12457), .S0(n68_adj_538));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_541_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_541_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_31 (.A0(n77_adj_605), .B0(n13820), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_604), .B1(n13820), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12456), .COUT(n12457), .S0(n74_adj_540), 
          .S1(n71_adj_539));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_29 (.A0(n83_adj_607), .B0(n13820), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_606), .B1(n13820), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12455), .COUT(n12456), .S0(n80_adj_542), 
          .S1(n77_adj_541));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_27 (.A0(n89_adj_609), .B0(n13820), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_608), .B1(n13820), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12454), .COUT(n12455), .S0(n86_adj_544), 
          .S1(n83_adj_543));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_25 (.A0(n95_adj_611), .B0(n13820), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_610), .B1(n13820), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12453), .COUT(n12454), .S0(n92_adj_546), 
          .S1(n89_adj_545));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_23 (.A0(n101_adj_613), .B0(n13820), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_612), .B1(n13820), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12452), .COUT(n12453), .S0(n98_adj_548), 
          .S1(n95_adj_547));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_21 (.A0(n107_adj_615), .B0(n13820), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_614), .B1(n13820), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12451), .COUT(n12452), .S0(n104_adj_550), 
          .S1(n101_adj_549));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_19 (.A0(n113_adj_617), .B0(n13820), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_616), .B1(n13820), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12450), .COUT(n12451), .S0(n110_adj_552), 
          .S1(n107_adj_551));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_17 (.A0(n119_adj_619), .B0(n13820), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_618), .B1(n13820), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12449), .COUT(n12450), .S0(n116_adj_554), 
          .S1(n113_adj_553));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_15 (.A0(n125_adj_621), .B0(n13820), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_620), .B1(n13820), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12448), .COUT(n12449), .S0(n122_adj_556), 
          .S1(n119_adj_555));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_13 (.A0(n131_adj_623), .B0(n13820), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_622), .B1(n13820), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12447), .COUT(n12448), .S0(n128_adj_558), 
          .S1(n125_adj_557));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_11 (.A0(n137_adj_625), .B0(n13820), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_624), .B1(n13820), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12446), .COUT(n12447), .S0(n134_adj_560), 
          .S1(n131_adj_559));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_9 (.A0(n143_adj_627), .B0(n13820), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_626), .B1(n13820), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12445), .COUT(n12446), .S0(n140_adj_562), 
          .S1(n137_adj_561));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_7 (.A0(n149_adj_629), .B0(n13820), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_628), .B1(n13820), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12444), .COUT(n12445), .S0(n146_adj_564), 
          .S1(n143_adj_563));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_5 (.A0(n155_adj_631), .B0(n13820), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_630), .B1(n13820), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12443), .COUT(n12444), .S0(n152_adj_566), 
          .S1(n149_adj_565));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_3 (.A0(n161_adj_633), .B0(n13820), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_632), .B1(n13820), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12442), .COUT(n12443), .S0(n158_adj_568), 
          .S1(n155_adj_567));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_541_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_541_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13820), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12442), .S1(n161_adj_569));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_541_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_541_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_541_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_541_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_33 (.A0(n74_adj_412), .B0(n2650), .C0(n71_adj_284), 
          .D0(n3489), .A1(n71_adj_411), .B1(n2650), .C1(n68_adj_283), 
          .D1(n3488), .CIN(n12440), .S0(n71_adj_316), .S1(n68_adj_315));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_33.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_33.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_31 (.A0(n80_adj_414), .B0(n2650), .C0(n77_adj_286), 
          .D0(n3491), .A1(n77_adj_413), .B1(n2650), .C1(n74_adj_285), 
          .D1(n3490), .CIN(n12439), .COUT(n12440), .S0(n77_adj_318), 
          .S1(n74_adj_317));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_29 (.A0(n86_adj_416), .B0(n2650), .C0(n83_adj_288), 
          .D0(n3493), .A1(n83_adj_415), .B1(n2650), .C1(n80_adj_287), 
          .D1(n3492), .CIN(n12438), .COUT(n12439), .S0(n83_adj_320), 
          .S1(n80_adj_319));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_27 (.A0(n92_adj_418), .B0(n2650), .C0(n89_adj_290), 
          .D0(n3495), .A1(n89_adj_417), .B1(n2650), .C1(n86_adj_289), 
          .D1(n3494), .CIN(n12437), .COUT(n12438), .S0(n89_adj_322), 
          .S1(n86_adj_321));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_25 (.A0(n98_adj_420), .B0(n2650), .C0(n95_adj_292), 
          .D0(n3497), .A1(n95_adj_419), .B1(n2650), .C1(n92_adj_291), 
          .D1(n3496), .CIN(n12436), .COUT(n12437), .S0(n95_adj_324), 
          .S1(n92_adj_323));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_23 (.A0(n104_adj_422), .B0(n2650), .C0(n101_adj_294), 
          .D0(n3499), .A1(n101_adj_421), .B1(n2650), .C1(n98_adj_293), 
          .D1(n3498), .CIN(n12435), .COUT(n12436), .S0(n101_adj_326), 
          .S1(n98_adj_325));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_21 (.A0(n110_adj_424), .B0(n2650), .C0(n107_adj_296), 
          .D0(n3501), .A1(n107_adj_423), .B1(n2650), .C1(n104_adj_295), 
          .D1(n3500), .CIN(n12434), .COUT(n12435), .S0(n107_adj_328), 
          .S1(n104_adj_327));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_19 (.A0(n116_adj_426), .B0(n2650), .C0(n113_adj_298), 
          .D0(n3503), .A1(n113_adj_425), .B1(n2650), .C1(n110_adj_297), 
          .D1(n3502), .CIN(n12433), .COUT(n12434), .S0(n113_adj_330), 
          .S1(n110_adj_329));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_17 (.A0(n122_adj_428), .B0(n2650), .C0(n119_adj_300), 
          .D0(n3505), .A1(n119_adj_427), .B1(n2650), .C1(n116_adj_299), 
          .D1(n3504), .CIN(n12432), .COUT(n12433), .S0(n119_adj_332), 
          .S1(n116_adj_331));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_15 (.A0(n128_adj_430), .B0(n2650), .C0(n125_adj_302), 
          .D0(n3507), .A1(n125_adj_429), .B1(n2650), .C1(n122_adj_301), 
          .D1(n3506), .CIN(n12431), .COUT(n12432), .S0(n125_adj_334), 
          .S1(n122_adj_333));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_13 (.A0(n134_adj_432), .B0(n2650), .C0(n131_adj_304), 
          .D0(n3509), .A1(n131_adj_431), .B1(n2650), .C1(n128_adj_303), 
          .D1(n3508), .CIN(n12430), .COUT(n12431), .S0(n131_adj_336), 
          .S1(n128_adj_335));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_11 (.A0(n140_adj_434), .B0(n2650), .C0(n137_adj_306), 
          .D0(n3511), .A1(n137_adj_433), .B1(n2650), .C1(n134_adj_305), 
          .D1(n3510), .CIN(n12429), .COUT(n12430), .S0(n137_adj_338), 
          .S1(n134_adj_337));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_9 (.A0(n146_adj_436), .B0(n2650), .C0(n143_adj_308), 
          .D0(n3513), .A1(n143_adj_435), .B1(n2650), .C1(n140_adj_307), 
          .D1(n3512), .CIN(n12428), .COUT(n12429), .S0(n143_adj_340), 
          .S1(n140_adj_339));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_7 (.A0(n152_adj_438), .B0(n2650), .C0(n149_adj_310), 
          .D0(n3515), .A1(n149_adj_437), .B1(n2650), .C1(n146_adj_309), 
          .D1(n3514), .CIN(n12427), .COUT(n12428), .S0(n149_adj_342), 
          .S1(n146_adj_341));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_5 (.A0(n158_adj_440), .B0(n2650), .C0(n155_adj_312), 
          .D0(n3517), .A1(n155_adj_439), .B1(n2650), .C1(n152_adj_311), 
          .D1(n3516), .CIN(n12426), .COUT(n12427), .S0(n155_adj_344), 
          .S1(n152_adj_343));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_559_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_3 (.A0(det_q4_28[0]), .B0(n2650), .C0(n161_adj_314), 
          .D0(n3519), .A1(n161_adj_441), .B1(n2650), .C1(n158_adj_313), 
          .D1(n3518), .CIN(n12425), .COUT(n12426), .S0(n161_adj_346), 
          .S1(n158_adj_345));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_559_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_559_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_559_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2650), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12425));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_559_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_559_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_559_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_559_add_4_1.INJECT1_1 = "NO";
    CCU2C add_586_add_4_34 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12421), .S0(n1410));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_34.INIT0 = 16'hffff;
    defparam add_586_add_4_34.INIT1 = 16'h0000;
    defparam add_586_add_4_34.INJECT1_0 = "NO";
    defparam add_586_add_4_34.INJECT1_1 = "NO";
    CCU2C add_586_add_4_32 (.A0(det_q4_28[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12420), .COUT(n12421), .S0(n1412), .S1(n1411));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_32.INIT0 = 16'h5555;
    defparam add_586_add_4_32.INIT1 = 16'h5555;
    defparam add_586_add_4_32.INJECT1_0 = "NO";
    defparam add_586_add_4_32.INJECT1_1 = "NO";
    CCU2C add_586_add_4_30 (.A0(det_q4_28[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12419), .COUT(n12420), .S0(n1414), .S1(n1413));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_30.INIT0 = 16'h5555;
    defparam add_586_add_4_30.INIT1 = 16'h5555;
    defparam add_586_add_4_30.INJECT1_0 = "NO";
    defparam add_586_add_4_30.INJECT1_1 = "NO";
    CCU2C add_586_add_4_28 (.A0(det_q4_28[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12418), .COUT(n12419), .S0(n1416), .S1(n1415));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_28.INIT0 = 16'h5555;
    defparam add_586_add_4_28.INIT1 = 16'h5555;
    defparam add_586_add_4_28.INJECT1_0 = "NO";
    defparam add_586_add_4_28.INJECT1_1 = "NO";
    CCU2C add_586_add_4_26 (.A0(det_q4_28[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12417), .COUT(n12418), .S0(n1418), .S1(n1417));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_26.INIT0 = 16'h5555;
    defparam add_586_add_4_26.INIT1 = 16'h5555;
    defparam add_586_add_4_26.INJECT1_0 = "NO";
    defparam add_586_add_4_26.INJECT1_1 = "NO";
    CCU2C add_586_add_4_24 (.A0(det_q4_28[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12416), .COUT(n12417), .S0(n1420), .S1(n1419));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_24.INIT0 = 16'h5555;
    defparam add_586_add_4_24.INIT1 = 16'h5555;
    defparam add_586_add_4_24.INJECT1_0 = "NO";
    defparam add_586_add_4_24.INJECT1_1 = "NO";
    CCU2C add_586_add_4_22 (.A0(det_q4_28[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12415), .COUT(n12416), .S0(n1422), .S1(n1421));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_22.INIT0 = 16'h5555;
    defparam add_586_add_4_22.INIT1 = 16'h5555;
    defparam add_586_add_4_22.INJECT1_0 = "NO";
    defparam add_586_add_4_22.INJECT1_1 = "NO";
    CCU2C add_586_add_4_20 (.A0(det_q4_28[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12414), .COUT(n12415), .S0(n1424), .S1(n1423));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_20.INIT0 = 16'h5555;
    defparam add_586_add_4_20.INIT1 = 16'h5555;
    defparam add_586_add_4_20.INJECT1_0 = "NO";
    defparam add_586_add_4_20.INJECT1_1 = "NO";
    CCU2C add_586_add_4_18 (.A0(det_q4_28[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12413), .COUT(n12414), .S0(n1426), .S1(n1425));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_18.INIT0 = 16'h5555;
    defparam add_586_add_4_18.INIT1 = 16'h5555;
    defparam add_586_add_4_18.INJECT1_0 = "NO";
    defparam add_586_add_4_18.INJECT1_1 = "NO";
    CCU2C add_586_add_4_16 (.A0(det_q4_28[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12412), .COUT(n12413), .S0(n1428), .S1(n1427));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_16.INIT0 = 16'h5555;
    defparam add_586_add_4_16.INIT1 = 16'h5555;
    defparam add_586_add_4_16.INJECT1_0 = "NO";
    defparam add_586_add_4_16.INJECT1_1 = "NO";
    CCU2C add_586_add_4_14 (.A0(det_q4_28[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12411), .COUT(n12412), .S0(n1430), .S1(n1429));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_14.INIT0 = 16'h5555;
    defparam add_586_add_4_14.INIT1 = 16'h5555;
    defparam add_586_add_4_14.INJECT1_0 = "NO";
    defparam add_586_add_4_14.INJECT1_1 = "NO";
    CCU2C add_586_add_4_12 (.A0(det_q4_28[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12410), .COUT(n12411), .S0(n1432), .S1(n1431));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_12.INIT0 = 16'h5555;
    defparam add_586_add_4_12.INIT1 = 16'h5555;
    defparam add_586_add_4_12.INJECT1_0 = "NO";
    defparam add_586_add_4_12.INJECT1_1 = "NO";
    CCU2C add_586_add_4_10 (.A0(det_q4_28[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12409), .COUT(n12410), .S0(n1434), .S1(n1433));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_10.INIT0 = 16'h5555;
    defparam add_586_add_4_10.INIT1 = 16'h5555;
    defparam add_586_add_4_10.INJECT1_0 = "NO";
    defparam add_586_add_4_10.INJECT1_1 = "NO";
    CCU2C add_586_add_4_8 (.A0(det_q4_28[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12408), .COUT(n12409), .S0(n1436), .S1(n1435));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_8.INIT0 = 16'h5555;
    defparam add_586_add_4_8.INIT1 = 16'h5555;
    defparam add_586_add_4_8.INJECT1_0 = "NO";
    defparam add_586_add_4_8.INJECT1_1 = "NO";
    CCU2C add_586_add_4_6 (.A0(det_q4_28[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12407), .COUT(n12408), .S0(n1438), .S1(n1437));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_6.INIT0 = 16'h5555;
    defparam add_586_add_4_6.INIT1 = 16'h5555;
    defparam add_586_add_4_6.INJECT1_0 = "NO";
    defparam add_586_add_4_6.INJECT1_1 = "NO";
    CCU2C add_586_add_4_4 (.A0(det_q4_28[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12406), .COUT(n12407), .S0(n1440), .S1(n1439));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_4.INIT0 = 16'h5555;
    defparam add_586_add_4_4.INIT1 = 16'h5555;
    defparam add_586_add_4_4.INJECT1_0 = "NO";
    defparam add_586_add_4_4.INJECT1_1 = "NO";
    CCU2C add_586_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(det_q4_28[1]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12406), .S1(n1441));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_586_add_4_2.INIT0 = 16'h000f;
    defparam add_586_add_4_2.INIT1 = 16'h5555;
    defparam add_586_add_4_2.INJECT1_0 = "NO";
    defparam add_586_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_33 (.A0(n1444), .B0(n13821), .C0(n71_adj_635), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12405), .S0(n68_adj_570));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_538_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_538_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_31 (.A0(n77_adj_637), .B0(n13821), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_636), .B1(n13821), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12404), .COUT(n12405), .S0(n74_adj_572), 
          .S1(n71_adj_571));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_29 (.A0(n83_adj_639), .B0(n13821), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_638), .B1(n13821), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12403), .COUT(n12404), .S0(n80_adj_574), 
          .S1(n77_adj_573));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_29.INJECT1_1 = "NO";
    FD1S3AX d2_reg_15__I_0_e2__i3 (.D(d1_reg[2]), .CK(clk_c), .Q(n126_adj_233));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i3.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i4 (.D(d1_reg[3]), .CK(clk_c), .Q(n124_adj_234));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i4.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i5 (.D(d1_reg[4]), .CK(clk_c), .Q(n122_adj_235));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i5.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i6 (.D(d1_reg[5]), .CK(clk_c), .Q(n120_adj_236));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i6.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i7 (.D(d1_reg[6]), .CK(clk_c), .Q(n118_adj_237));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i7.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i8 (.D(d1_reg[7]), .CK(clk_c), .Q(n116_adj_238));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i8.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i9 (.D(d1_reg[8]), .CK(clk_c), .Q(n114_adj_239));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i9.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i10 (.D(d1_reg[9]), .CK(clk_c), .Q(n112_adj_240));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i10.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i11 (.D(d1_reg[10]), .CK(clk_c), .Q(n110_adj_241));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i11.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i12 (.D(d1_reg[11]), .CK(clk_c), .Q(n108_adj_242));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i12.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i13 (.D(d1_reg[12]), .CK(clk_c), .Q(n106_adj_230));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i13.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i14 (.D(d1_reg[13]), .CK(clk_c), .Q(n104_adj_243));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i14.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i15 (.D(d1_reg[14]), .CK(clk_c), .Q(n102_adj_244));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i15.GSR = "ENABLED";
    FD1S3AX d2_reg_15__I_0_e2__i16 (.D(d1_reg[15]), .CK(clk_c), .Q(n68_adj_245));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(101[44:57])
    defparam d2_reg_15__I_0_e2__i16.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i2 (.D(a1_reg[1]), .CK(clk_c), .Q(n128));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i2.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i3 (.D(a1_reg[2]), .CK(clk_c), .Q(n126));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i3.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i4 (.D(a1_reg[3]), .CK(clk_c), .Q(n124));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i4.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i5 (.D(a1_reg[4]), .CK(clk_c), .Q(n122));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i5.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i6 (.D(a1_reg[5]), .CK(clk_c), .Q(n120));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i6.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i7 (.D(a1_reg[6]), .CK(clk_c), .Q(n118));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i7.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i8 (.D(a1_reg[7]), .CK(clk_c), .Q(n116));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i8.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i9 (.D(a1_reg[8]), .CK(clk_c), .Q(n114));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i9.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i10 (.D(a1_reg[9]), .CK(clk_c), .Q(n112));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i10.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i11 (.D(a1_reg[10]), .CK(clk_c), .Q(n110));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i11.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i12 (.D(a1_reg[11]), .CK(clk_c), .Q(n108));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i12.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i13 (.D(a1_reg[12]), .CK(clk_c), .Q(n106));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i13.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i14 (.D(a1_reg[13]), .CK(clk_c), .Q(n104));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i14.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i15 (.D(a1_reg[14]), .CK(clk_c), .Q(n102));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i15.GSR = "ENABLED";
    FD1S3AX a2_reg_15__I_0_e2__i16 (.D(a1_reg[15]), .CK(clk_c), .Q(n68));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(104[44:57])
    defparam a2_reg_15__I_0_e2__i16.GSR = "ENABLED";
    FD1S3AX det_q4_28_i5 (.D(det_q4_28_31__N_65[5]), .CK(clk_c), .Q(det_q4_28[5]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(56[18] 65[12])
    defparam det_q4_28_i5.GSR = "ENABLED";
    CCU2C _add_1_538_add_4_27 (.A0(n89_adj_641), .B0(n13821), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_640), .B1(n13821), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12402), .COUT(n12403), .S0(n86_adj_576), 
          .S1(n83_adj_575));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_25 (.A0(n95_adj_643), .B0(n13821), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_642), .B1(n13821), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12401), .COUT(n12402), .S0(n92_adj_578), 
          .S1(n89_adj_577));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_23 (.A0(n101_adj_645), .B0(n13821), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_644), .B1(n13821), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12400), .COUT(n12401), .S0(n98_adj_580), 
          .S1(n95_adj_579));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_21 (.A0(n107_adj_647), .B0(n13821), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_646), .B1(n13821), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12399), .COUT(n12400), .S0(n104_adj_582), 
          .S1(n101_adj_581));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_19 (.A0(n113_adj_649), .B0(n13821), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_648), .B1(n13821), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12398), .COUT(n12399), .S0(n110_adj_584), 
          .S1(n107_adj_583));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_17 (.A0(n119_adj_651), .B0(n13821), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_650), .B1(n13821), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12397), .COUT(n12398), .S0(n116_adj_586), 
          .S1(n113_adj_585));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_15 (.A0(n125_adj_653), .B0(n13821), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_652), .B1(n13821), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12396), .COUT(n12397), .S0(n122_adj_588), 
          .S1(n119_adj_587));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_13 (.A0(n131_adj_655), .B0(n13821), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_654), .B1(n13821), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12395), .COUT(n12396), .S0(n128_adj_590), 
          .S1(n125_adj_589));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_11 (.A0(n137_adj_657), .B0(n13821), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_656), .B1(n13821), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12394), .COUT(n12395), .S0(n134_adj_592), 
          .S1(n131_adj_591));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_9 (.A0(n143_adj_659), .B0(n13821), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_658), .B1(n13821), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12393), .COUT(n12394), .S0(n140_adj_594), 
          .S1(n137_adj_593));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_7 (.A0(n149_adj_661), .B0(n13821), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_660), .B1(n13821), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12392), .COUT(n12393), .S0(n146_adj_596), 
          .S1(n143_adj_595));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_5 (.A0(n155_adj_663), .B0(n13821), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_662), .B1(n13821), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12391), .COUT(n12392), .S0(n152_adj_598), 
          .S1(n149_adj_597));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_3 (.A0(n161_adj_665), .B0(n13821), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_664), .B1(n13821), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12390), .COUT(n12391), .S0(n158_adj_600), 
          .S1(n155_adj_599));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_538_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_538_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13821), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12390), .S1(n161_adj_601));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_538_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_538_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_538_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_538_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_33 (.A0(n1444), .B0(n13821), .C0(n71_adj_667), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12389), .S0(n68_adj_602));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_535_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_535_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_31 (.A0(n77_adj_669), .B0(n13821), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_668), .B1(n13821), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12388), .COUT(n12389), .S0(n74_adj_604), 
          .S1(n71_adj_603));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_29 (.A0(n83_adj_671), .B0(n13821), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_670), .B1(n13821), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12387), .COUT(n12388), .S0(n80_adj_606), 
          .S1(n77_adj_605));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_27 (.A0(n89_adj_673), .B0(n13821), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_672), .B1(n13821), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12386), .COUT(n12387), .S0(n86_adj_608), 
          .S1(n83_adj_607));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_25 (.A0(n95_adj_675), .B0(n13821), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_674), .B1(n13821), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12385), .COUT(n12386), .S0(n92_adj_610), 
          .S1(n89_adj_609));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_23 (.A0(n101_adj_677), .B0(n13821), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_676), .B1(n13821), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12384), .COUT(n12385), .S0(n98_adj_612), 
          .S1(n95_adj_611));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_21 (.A0(n107_adj_679), .B0(n13821), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_678), .B1(n13821), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12383), .COUT(n12384), .S0(n104_adj_614), 
          .S1(n101_adj_613));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_19 (.A0(n113_adj_681), .B0(n13821), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_680), .B1(n13821), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12382), .COUT(n12383), .S0(n110_adj_616), 
          .S1(n107_adj_615));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_17 (.A0(n119_adj_683), .B0(n13821), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_682), .B1(n13821), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12381), .COUT(n12382), .S0(n116_adj_618), 
          .S1(n113_adj_617));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_15 (.A0(n125_adj_685), .B0(n13821), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_684), .B1(n13821), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12380), .COUT(n12381), .S0(n122_adj_620), 
          .S1(n119_adj_619));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_13 (.A0(n131_adj_687), .B0(n13821), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_686), .B1(n13821), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12379), .COUT(n12380), .S0(n128_adj_622), 
          .S1(n125_adj_621));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_11 (.A0(n137_adj_689), .B0(n13821), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_688), .B1(n13821), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12378), .COUT(n12379), .S0(n134_adj_624), 
          .S1(n131_adj_623));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_9 (.A0(n143_adj_691), .B0(n13821), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_690), .B1(n13821), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12377), .COUT(n12378), .S0(n140_adj_626), 
          .S1(n137_adj_625));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_7 (.A0(n149_adj_693), .B0(n13821), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_692), .B1(n13821), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12376), .COUT(n12377), .S0(n146_adj_628), 
          .S1(n143_adj_627));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_5 (.A0(n155_adj_695), .B0(n13821), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_694), .B1(n13821), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12375), .COUT(n12376), .S0(n152_adj_630), 
          .S1(n149_adj_629));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_3 (.A0(n161_adj_697), .B0(n13821), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_696), .B1(n13821), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12374), .COUT(n12375), .S0(n158_adj_632), 
          .S1(n155_adj_631));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_535_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_535_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13821), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12374), .S1(n161_adj_633));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_535_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_535_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_535_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_535_add_4_1.INJECT1_1 = "NO";
    LUT4 i1573_2_lut_4_lut (.A(n68_adj_1018), .B(n68_adj_986), .C(n1410), 
         .D(inv_det_31__N_227), .Z(n35)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1573_2_lut_4_lut.init = 16'h0035;
    LUT4 i1576_2_lut_4_lut (.A(n68_adj_1082), .B(n68_adj_1050), .C(n1410), 
         .D(inv_det_31__N_227), .Z(n34)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1576_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_329_i1_3_lut_rep_89 (.A(n68_adj_1082), .B(n68_adj_1050), .C(n1410), 
         .Z(n13839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_329_i1_3_lut_rep_89.init = 16'hcaca;
    LUT4 mux_328_i1_3_lut_rep_90 (.A(n68_adj_1146), .B(n68_adj_1114), .C(n1410), 
         .Z(n13840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_328_i1_3_lut_rep_90.init = 16'hcaca;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    reciprocal_q16_16 u_recip (.n1474(n1474), .det_q4_28({det_q4_28}), .n13829(n13829), 
            .n2379(n2379), .error_recip(error_recip), .clk_c(clk_c), .inv_det_31__N_227(inv_det_31__N_227), 
            .n1465(n1465), .n13836(n13836), .n1834(n1834), .n1464(n1464), 
            .n1833(n1833), .n1473(n1473), .n2378(n2378), .n1472(n1472), 
            .n2377(n2377), .n1471(n1471), .n2376(n2376), .n1470(n1470), 
            .n2375(n2375), .n1469(n1469), .n2374(n2374), .n1468(n1468), 
            .n2373(n2373), .n1467(n1467), .n2372(n2372), .n1466(n1466), 
            .n2371(n2371), .n2370(n2370), .n2369(n2369), .n1463(n1463), 
            .n2368(n2368), .n1462(n1462), .n2367(n2367), .n1461(n1461), 
            .n2366(n2366), .n1460(n1460), .n2365(n2365), .n1459(n1459), 
            .n2364(n2364), .n1458(n1458), .n2363(n2363), .n1457(n1457), 
            .n2362(n2362), .n1456(n1456), .n2361(n2361), .n1455(n1455), 
            .n2360(n2360), .n1454(n1454), .n2359(n2359), .n1453(n1453), 
            .n2358(n2358), .n1452(n1452), .n2357(n2357), .n1451(n1451), 
            .n2356(n2356), .n1450(n1450), .n2355(n2355), .n1449(n1449), 
            .n2354(n2354), .n1448(n1448), .n2353(n2353), .n1447(n1447), 
            .n2352(n2352), .n1832(n1832), .n1446(n1446), .n2351(n2351), 
            .n1445(n1445), .n2350(n2350), .n1475(n1475), .n1844(n1844), 
            .n1843(n1843), .n1842(n1842), .n1841(n1841), .n1840(n1840), 
            .n1839(n1839), .n1838(n1838), .n1837(n1837), .n1836(n1836), 
            .n1835(n1835), .n1831(n1831), .n1830(n1830), .n1829(n1829), 
            .n1828(n1828), .n1827(n1827), .n2382(n2382), .n46(n46), 
            .n1846(n1846), .n38(n38), .n2583(n2583), .n2616({n2617, 
            n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
            n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
            n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
            n2642, n2643, n2644, n2645, n2646, n2647, n2648}), 
            .n1444(n1444), .n1826(n1826), .n1825(n1825), .n1824(n1824), 
            .n1823(n1823), .n1822(n1822), .n1821(n1821), .n1820(n1820), 
            .n1819(n1819), .n1818(n1818), .n1817(n1817), .n1816(n1816), 
            .n1815(n1815), .n1814(n1814), .n68(n68_adj_1652), .n68_adj_1(n68_adj_1209), 
            .n68_adj_2(n68_adj_315), .n64(n64), .n63(n63), .n13818(n13818), 
            .n3422(n3422), .n3424(n3424), .n3423(n3423), .n3426(n3426), 
            .n3425(n3425), .n3428(n3428), .n3427(n3427), .n3430(n3430), 
            .n3429(n3429), .n3432(n3432), .n3431(n3431), .n3434(n3434), 
            .n3433(n3433), .n3436(n3436), .n3435(n3435), .n3438(n3438), 
            .n3437(n3437), .n3440(n3440), .n3439(n3439), .n3442(n3442), 
            .n3441(n3441), .n3444(n3444), .n3443(n3443), .n3446(n3446), 
            .n3445(n3445), .n3448(n3448), .n3447(n3447), .n3450(n3450), 
            .n3449(n3449), .n3452(n3452), .n3451(n3451), .n3454(n3454), 
            .n3487({n3488, n3489, n3490, n3491, n3492, n3493, n3494, 
            n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
            n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
            n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
            n3519}), .n62(n62), .n2650(n2650), .n50(n50), .n49(n49), 
            .n2449(n2449), .n47(n47), .n2516(n2516), .n48(n48), .GND_net(GND_net), 
            .n2380(n2380), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(86[23] 92[6])
    VLO i1 (.Z(GND_net));
    CCU2C _add_1_532_add_4_27 (.A0(n89_adj_705), .B0(n13822), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_704), .B1(n13822), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12622), .COUT(n12623), .S0(n86_adj_640), 
          .S1(n83_adj_639));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_29 (.A0(n83_adj_703), .B0(n13822), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_702), .B1(n13822), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12623), .COUT(n12624), .S0(n80_adj_638), 
          .S1(n77_adj_637));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_31 (.A0(n77_adj_701), .B0(n13822), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_700), .B1(n13822), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12624), .COUT(n12625), .S0(n74_adj_636), 
          .S1(n71_adj_635));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_532_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_532_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_532_add_4_33 (.A0(n1444), .B0(n13822), .C0(n71_adj_699), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12625), .S0(n68_adj_634));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_532_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_532_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_532_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_532_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13822), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12626), .S1(n161_adj_697));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_529_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_3 (.A0(n161_adj_761), .B0(n13822), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_760), .B1(n13822), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12626), .COUT(n12627), .S0(n158_adj_696), 
          .S1(n155_adj_695));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_5 (.A0(n155_adj_759), .B0(n13822), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_758), .B1(n13822), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12627), .COUT(n12628), .S0(n152_adj_694), 
          .S1(n149_adj_693));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_7 (.A0(n149_adj_757), .B0(n13822), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_756), .B1(n13822), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12628), .COUT(n12629), .S0(n146_adj_692), 
          .S1(n143_adj_691));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_9 (.A0(n143_adj_755), .B0(n13822), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_754), .B1(n13822), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12629), .COUT(n12630), .S0(n140_adj_690), 
          .S1(n137_adj_689));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_11 (.A0(n137_adj_753), .B0(n13822), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_752), .B1(n13822), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12630), .COUT(n12631), .S0(n134_adj_688), 
          .S1(n131_adj_687));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_13 (.A0(n131_adj_751), .B0(n13822), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_750), .B1(n13822), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12631), .COUT(n12632), .S0(n128_adj_686), 
          .S1(n125_adj_685));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_15 (.A0(n125_adj_749), .B0(n13822), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_748), .B1(n13822), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12632), .COUT(n12633), .S0(n122_adj_684), 
          .S1(n119_adj_683));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_17 (.A0(n119_adj_747), .B0(n13822), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_746), .B1(n13822), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12633), .COUT(n12634), .S0(n116_adj_682), 
          .S1(n113_adj_681));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_19 (.A0(n113_adj_745), .B0(n13822), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_744), .B1(n13822), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12634), .COUT(n12635), .S0(n110_adj_680), 
          .S1(n107_adj_679));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_21 (.A0(n107_adj_743), .B0(n13822), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_742), .B1(n13822), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12635), .COUT(n12636), .S0(n104_adj_678), 
          .S1(n101_adj_677));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_23 (.A0(n101_adj_741), .B0(n13822), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_740), .B1(n13822), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12636), .COUT(n12637), .S0(n98_adj_676), 
          .S1(n95_adj_675));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_25 (.A0(n95_adj_739), .B0(n13822), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_738), .B1(n13822), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12637), .COUT(n12638), .S0(n92_adj_674), 
          .S1(n89_adj_673));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_27 (.A0(n89_adj_737), .B0(n13822), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_736), .B1(n13822), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12638), .COUT(n12639), .S0(n86_adj_672), 
          .S1(n83_adj_671));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_29 (.A0(n83_adj_735), .B0(n13822), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_734), .B1(n13822), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12639), .COUT(n12640), .S0(n80_adj_670), 
          .S1(n77_adj_669));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_31 (.A0(n77_adj_733), .B0(n13822), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_732), .B1(n13822), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12640), .COUT(n12641), .S0(n74_adj_668), 
          .S1(n71_adj_667));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_529_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_529_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_529_add_4_33 (.A0(n1444), .B0(n13822), .C0(n71_adj_731), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12641), .S0(n68_adj_666));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_529_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_529_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_529_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_529_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13823), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12642), .S1(n161_adj_729));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_526_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_3 (.A0(n161_adj_793), .B0(n13823), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_792), .B1(n13823), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12642), .COUT(n12643), .S0(n158_adj_728), 
          .S1(n155_adj_727));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_5 (.A0(n155_adj_791), .B0(n13823), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_790), .B1(n13823), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12643), .COUT(n12644), .S0(n152_adj_726), 
          .S1(n149_adj_725));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_7 (.A0(n149_adj_789), .B0(n13823), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_788), .B1(n13823), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12644), .COUT(n12645), .S0(n146_adj_724), 
          .S1(n143_adj_723));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_9 (.A0(n143_adj_787), .B0(n13823), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_786), .B1(n13823), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12645), .COUT(n12646), .S0(n140_adj_722), 
          .S1(n137_adj_721));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_11 (.A0(n137_adj_785), .B0(n13823), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_784), .B1(n13823), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12646), .COUT(n12647), .S0(n134_adj_720), 
          .S1(n131_adj_719));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_13 (.A0(n131_adj_783), .B0(n13823), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_782), .B1(n13823), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12647), .COUT(n12648), .S0(n128_adj_718), 
          .S1(n125_adj_717));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_15 (.A0(n125_adj_781), .B0(n13823), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_780), .B1(n13823), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12648), .COUT(n12649), .S0(n122_adj_716), 
          .S1(n119_adj_715));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_17 (.A0(n119_adj_779), .B0(n13823), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_778), .B1(n13823), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12649), .COUT(n12650), .S0(n116_adj_714), 
          .S1(n113_adj_713));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_19 (.A0(n113_adj_777), .B0(n13823), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_776), .B1(n13823), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12650), .COUT(n12651), .S0(n110_adj_712), 
          .S1(n107_adj_711));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_21 (.A0(n107_adj_775), .B0(n13823), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_774), .B1(n13823), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12651), .COUT(n12652), .S0(n104_adj_710), 
          .S1(n101_adj_709));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_23 (.A0(n101_adj_773), .B0(n13823), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_772), .B1(n13823), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12652), .COUT(n12653), .S0(n98_adj_708), 
          .S1(n95_adj_707));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_25 (.A0(n95_adj_771), .B0(n13823), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_770), .B1(n13823), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12653), .COUT(n12654), .S0(n92_adj_706), 
          .S1(n89_adj_705));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_27 (.A0(n89_adj_769), .B0(n13823), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_768), .B1(n13823), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12654), .COUT(n12655), .S0(n86_adj_704), 
          .S1(n83_adj_703));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_29 (.A0(n83_adj_767), .B0(n13823), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_766), .B1(n13823), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12655), .COUT(n12656), .S0(n80_adj_702), 
          .S1(n77_adj_701));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_31 (.A0(n77_adj_765), .B0(n13823), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_764), .B1(n13823), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12656), .COUT(n12657), .S0(n74_adj_700), 
          .S1(n71_adj_699));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_526_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_526_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_526_add_4_33 (.A0(n1444), .B0(n13823), .C0(n71_adj_763), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12657), .S0(n68_adj_698));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_526_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_526_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_526_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_526_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13823), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12658), .S1(n161_adj_761));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_523_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_3 (.A0(n161_adj_857), .B0(n13823), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_856), .B1(n13823), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12658), .COUT(n12659), .S0(n158_adj_760), 
          .S1(n155_adj_759));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_5 (.A0(n155_adj_855), .B0(n13823), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_854), .B1(n13823), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12659), .COUT(n12660), .S0(n152_adj_758), 
          .S1(n149_adj_757));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_7 (.A0(n149_adj_853), .B0(n13823), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_852), .B1(n13823), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12660), .COUT(n12661), .S0(n146_adj_756), 
          .S1(n143_adj_755));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_9 (.A0(n143_adj_851), .B0(n13823), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_850), .B1(n13823), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12661), .COUT(n12662), .S0(n140_adj_754), 
          .S1(n137_adj_753));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_11 (.A0(n137_adj_849), .B0(n13823), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_848), .B1(n13823), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12662), .COUT(n12663), .S0(n134_adj_752), 
          .S1(n131_adj_751));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_13 (.A0(n131_adj_847), .B0(n13823), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_846), .B1(n13823), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12663), .COUT(n12664), .S0(n128_adj_750), 
          .S1(n125_adj_749));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_15 (.A0(n125_adj_845), .B0(n13823), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_844), .B1(n13823), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12664), .COUT(n12665), .S0(n122_adj_748), 
          .S1(n119_adj_747));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_17 (.A0(n119_adj_843), .B0(n13823), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_842), .B1(n13823), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12665), .COUT(n12666), .S0(n116_adj_746), 
          .S1(n113_adj_745));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_19 (.A0(n113_adj_841), .B0(n13823), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_840), .B1(n13823), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12666), .COUT(n12667), .S0(n110_adj_744), 
          .S1(n107_adj_743));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_21 (.A0(n107_adj_839), .B0(n13823), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_838), .B1(n13823), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12667), .COUT(n12668), .S0(n104_adj_742), 
          .S1(n101_adj_741));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_23 (.A0(n101_adj_837), .B0(n13823), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_836), .B1(n13823), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12668), .COUT(n12669), .S0(n98_adj_740), 
          .S1(n95_adj_739));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_25 (.A0(n95_adj_835), .B0(n13823), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_834), .B1(n13823), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12669), .COUT(n12670), .S0(n92_adj_738), 
          .S1(n89_adj_737));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_27 (.A0(n89_adj_833), .B0(n13823), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_832), .B1(n13823), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12670), .COUT(n12671), .S0(n86_adj_736), 
          .S1(n83_adj_735));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_29 (.A0(n83_adj_831), .B0(n13823), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_830), .B1(n13823), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12671), .COUT(n12672), .S0(n80_adj_734), 
          .S1(n77_adj_733));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_31 (.A0(n77_adj_829), .B0(n13823), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_828), .B1(n13823), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12672), .COUT(n12673), .S0(n74_adj_732), 
          .S1(n71_adj_731));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_523_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_523_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_523_add_4_33 (.A0(n1444), .B0(n13823), .C0(n71_adj_827), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12673), .S0(n68_adj_730));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_523_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_523_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_523_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_523_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13824), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12674), .S1(n161_adj_793));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_520_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_3 (.A0(n161_adj_1716), .B0(n13824), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1715), .B1(n13824), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12674), .COUT(n12675), .S0(n158_adj_792), 
          .S1(n155_adj_791));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_5 (.A0(n155_adj_1714), .B0(n13824), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1713), .B1(n13824), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12675), .COUT(n12676), .S0(n152_adj_790), 
          .S1(n149_adj_789));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_7 (.A0(n149_adj_1712), .B0(n13824), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1711), .B1(n13824), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12676), .COUT(n12677), .S0(n146_adj_788), 
          .S1(n143_adj_787));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_9 (.A0(n143_adj_1710), .B0(n13824), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1709), .B1(n13824), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12677), .COUT(n12678), .S0(n140_adj_786), 
          .S1(n137_adj_785));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_11 (.A0(n137_adj_1708), .B0(n13824), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1707), .B1(n13824), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12678), .COUT(n12679), .S0(n134_adj_784), 
          .S1(n131_adj_783));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_13 (.A0(n131_adj_1706), .B0(n13824), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1705), .B1(n13824), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12679), .COUT(n12680), .S0(n128_adj_782), 
          .S1(n125_adj_781));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_15 (.A0(n125_adj_1704), .B0(n13824), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1703), .B1(n13824), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12680), .COUT(n12681), .S0(n122_adj_780), 
          .S1(n119_adj_779));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_17 (.A0(n119_adj_1702), .B0(n13824), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1701), .B1(n13824), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12681), .COUT(n12682), .S0(n116_adj_778), 
          .S1(n113_adj_777));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_19 (.A0(n113_adj_1700), .B0(n13824), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1699), .B1(n13824), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12682), .COUT(n12683), .S0(n110_adj_776), 
          .S1(n107_adj_775));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_21 (.A0(n107_adj_1698), .B0(n13824), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1697), .B1(n13824), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12683), .COUT(n12684), .S0(n104_adj_774), 
          .S1(n101_adj_773));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_23 (.A0(n101_adj_1696), .B0(n13824), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1695), .B1(n13824), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12684), .COUT(n12685), .S0(n98_adj_772), 
          .S1(n95_adj_771));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_25 (.A0(n95_adj_1694), .B0(n13824), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1693), .B1(n13824), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12685), .COUT(n12686), .S0(n92_adj_770), 
          .S1(n89_adj_769));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_27 (.A0(n89_adj_1692), .B0(n13824), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1691), .B1(n13824), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12686), .COUT(n12687), .S0(n86_adj_768), 
          .S1(n83_adj_767));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_29 (.A0(n83_adj_1690), .B0(n13824), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1689), .B1(n13824), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12687), .COUT(n12688), .S0(n80_adj_766), 
          .S1(n77_adj_765));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_31 (.A0(n77_adj_1688), .B0(n13824), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1687), .B1(n13824), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12688), .COUT(n12689), .S0(n74_adj_764), 
          .S1(n71_adj_763));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_520_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_520_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_520_add_4_33 (.A0(n1444), .B0(n13824), .C0(n71_adj_1686), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12689), .S0(n68_adj_762));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_520_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_520_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_520_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_520_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13831), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12690), .S1(n161_adj_825));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_385_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_3 (.A0(n161_adj_1907), .B0(n13831), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1906), .B1(n13831), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12690), .COUT(n12691), .S0(n158_adj_824), 
          .S1(n155_adj_823));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_5 (.A0(n155_adj_1905), .B0(n13831), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1904), .B1(n13831), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12691), .COUT(n12692), .S0(n152_adj_822), 
          .S1(n149_adj_821));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_7 (.A0(n149_adj_1903), .B0(n13831), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1902), .B1(n13831), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12692), .COUT(n12693), .S0(n146_adj_820), 
          .S1(n143_adj_819));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_9 (.A0(n143_adj_1901), .B0(n13831), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1900), .B1(n13831), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12693), .COUT(n12694), .S0(n140_adj_818), 
          .S1(n137_adj_817));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_11 (.A0(n137_adj_1899), .B0(n13831), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1898), .B1(n13831), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12694), .COUT(n12695), .S0(n134_adj_816), 
          .S1(n131_adj_815));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_13 (.A0(n131_adj_1897), .B0(n13831), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1896), .B1(n13831), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12695), .COUT(n12696), .S0(n128_adj_814), 
          .S1(n125_adj_813));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_15 (.A0(n125_adj_1895), .B0(n13831), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1894), .B1(n13831), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12696), .COUT(n12697), .S0(n122_adj_812), 
          .S1(n119_adj_811));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_17 (.A0(n119_adj_1893), .B0(n13831), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1892), .B1(n13831), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12697), .COUT(n12698), .S0(n116_adj_810), 
          .S1(n113_adj_809));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_19 (.A0(n113_adj_1891), .B0(n13831), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1890), .B1(n13831), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12698), .COUT(n12699), .S0(n110_adj_808), 
          .S1(n107_adj_807));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_21 (.A0(n107_adj_1889), .B0(n13831), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1888), .B1(n13831), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12699), .COUT(n12700), .S0(n104_adj_806), 
          .S1(n101_adj_805));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_23 (.A0(n101_adj_1887), .B0(n13831), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1886), .B1(n13831), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12700), .COUT(n12701), .S0(n98_adj_804), 
          .S1(n95_adj_803));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_25 (.A0(n95_adj_1885), .B0(n13831), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1884), .B1(n13831), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12701), .COUT(n12702), .S0(n92_adj_802), 
          .S1(n89_adj_801));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_27 (.A0(n89_adj_1883), .B0(n13831), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1882), .B1(n13831), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12702), .COUT(n12703), .S0(n86_adj_800), 
          .S1(n83_adj_799));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_29 (.A0(n83_adj_1881), .B0(n13831), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1880), .B1(n13831), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12703), .COUT(n12704), .S0(n80_adj_798), 
          .S1(n77_adj_797));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_31 (.A0(n77_adj_1879), .B0(n13831), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1878), .B1(n13831), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12704), .COUT(n12705), .S0(n74_adj_796), 
          .S1(n71_adj_795));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_385_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_385_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_385_add_4_33 (.A0(n1444), .B0(n13831), .C0(n71_adj_1877), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12705), .S0(n68_adj_794));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_385_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_385_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_385_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_385_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13824), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12706), .S1(n161_adj_857));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_517_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_3 (.A0(n161_adj_1748), .B0(n13824), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1747), .B1(n13824), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12706), .COUT(n12707), .S0(n158_adj_856), 
          .S1(n155_adj_855));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_5 (.A0(n155_adj_1746), .B0(n13824), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1745), .B1(n13824), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12707), .COUT(n12708), .S0(n152_adj_854), 
          .S1(n149_adj_853));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_7 (.A0(n149_adj_1744), .B0(n13824), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1743), .B1(n13824), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12708), .COUT(n12709), .S0(n146_adj_852), 
          .S1(n143_adj_851));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_9 (.A0(n143_adj_1742), .B0(n13824), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1741), .B1(n13824), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12709), .COUT(n12710), .S0(n140_adj_850), 
          .S1(n137_adj_849));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_11 (.A0(n137_adj_1740), .B0(n13824), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1739), .B1(n13824), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12710), .COUT(n12711), .S0(n134_adj_848), 
          .S1(n131_adj_847));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_13 (.A0(n131_adj_1738), .B0(n13824), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1737), .B1(n13824), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12711), .COUT(n12712), .S0(n128_adj_846), 
          .S1(n125_adj_845));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_15 (.A0(n125_adj_1736), .B0(n13824), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1735), .B1(n13824), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12712), .COUT(n12713), .S0(n122_adj_844), 
          .S1(n119_adj_843));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_17 (.A0(n119_adj_1734), .B0(n13824), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1733), .B1(n13824), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12713), .COUT(n12714), .S0(n116_adj_842), 
          .S1(n113_adj_841));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_19 (.A0(n113_adj_1732), .B0(n13824), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1731), .B1(n13824), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12714), .COUT(n12715), .S0(n110_adj_840), 
          .S1(n107_adj_839));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_21 (.A0(n107_adj_1730), .B0(n13824), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1729), .B1(n13824), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12715), .COUT(n12716), .S0(n104_adj_838), 
          .S1(n101_adj_837));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_23 (.A0(n101_adj_1728), .B0(n13824), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1727), .B1(n13824), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12716), .COUT(n12717), .S0(n98_adj_836), 
          .S1(n95_adj_835));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_25 (.A0(n95_adj_1726), .B0(n13824), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1725), .B1(n13824), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12717), .COUT(n12718), .S0(n92_adj_834), 
          .S1(n89_adj_833));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_27 (.A0(n89_adj_1724), .B0(n13824), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1723), .B1(n13824), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12718), .COUT(n12719), .S0(n86_adj_832), 
          .S1(n83_adj_831));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_29 (.A0(n83_adj_1722), .B0(n13824), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1721), .B1(n13824), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12719), .COUT(n12720), .S0(n80_adj_830), 
          .S1(n77_adj_829));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_31 (.A0(n77_adj_1720), .B0(n13824), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1719), .B1(n13824), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12720), .COUT(n12721), .S0(n74_adj_828), 
          .S1(n71_adj_827));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_517_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_517_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_517_add_4_33 (.A0(n1444), .B0(n13824), .C0(n71_adj_1718), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12721), .S0(n68_adj_826));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_517_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_517_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_517_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_517_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13837), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12722), .S1(n161_adj_889));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_478_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_3 (.A0(n161_adj_953), .B0(n13837), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_952), .B1(n13837), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12722), .COUT(n12723), .S0(n158_adj_888), 
          .S1(n155_adj_887));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_5 (.A0(n155_adj_951), .B0(n13837), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_950), .B1(n13837), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12723), .COUT(n12724), .S0(n152_adj_886), 
          .S1(n149_adj_885));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_7 (.A0(n149_adj_949), .B0(n13837), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_948), .B1(n13837), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12724), .COUT(n12725), .S0(n146_adj_884), 
          .S1(n143_adj_883));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_9 (.A0(n143_adj_947), .B0(n13837), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_946), .B1(n13837), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12725), .COUT(n12726), .S0(n140_adj_882), 
          .S1(n137_adj_881));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_11 (.A0(n137_adj_945), .B0(n13837), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_944), .B1(n13837), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12726), .COUT(n12727), .S0(n134_adj_880), 
          .S1(n131_adj_879));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_13 (.A0(n131_adj_943), .B0(n13837), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_942), .B1(n13837), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12727), .COUT(n12728), .S0(n128_adj_878), 
          .S1(n125_adj_877));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_15 (.A0(n125_adj_941), .B0(n13837), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_940), .B1(n13837), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12728), .COUT(n12729), .S0(n122_adj_876), 
          .S1(n119_adj_875));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_17 (.A0(n119_adj_939), .B0(n13837), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_938), .B1(n13837), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12729), .COUT(n12730), .S0(n116_adj_874), 
          .S1(n113_adj_873));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_19 (.A0(n113_adj_937), .B0(n13837), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_936), .B1(n13837), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12730), .COUT(n12731), .S0(n110_adj_872), 
          .S1(n107_adj_871));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_21 (.A0(n107_adj_935), .B0(n13837), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_934), .B1(n13837), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12731), .COUT(n12732), .S0(n104_adj_870), 
          .S1(n101_adj_869));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_23 (.A0(n101_adj_933), .B0(n13837), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_932), .B1(n13837), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12732), .COUT(n12733), .S0(n98_adj_868), 
          .S1(n95_adj_867));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_25 (.A0(n95_adj_931), .B0(n13837), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_930), .B1(n13837), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12733), .COUT(n12734), .S0(n92_adj_866), 
          .S1(n89_adj_865));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_27 (.A0(n89_adj_929), .B0(n13837), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_928), .B1(n13837), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12734), .COUT(n12735), .S0(n86_adj_864), 
          .S1(n83_adj_863));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_29 (.A0(n83_adj_927), .B0(n13837), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_926), .B1(n13837), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12735), .COUT(n12736), .S0(n80_adj_862), 
          .S1(n77_adj_861));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_31 (.A0(n77_adj_925), .B0(n13837), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_924), .B1(n13837), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12736), .COUT(n12737), .S0(n74_adj_860), 
          .S1(n71_adj_859));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_478_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_478_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_478_add_4_33 (.A0(n1444), .B0(n13837), .C0(n71_adj_923), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12737), .S0(n68_adj_858));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_478_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_478_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_478_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_478_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13837), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12738), .S1(n161_adj_921));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_475_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_3 (.A0(n161_adj_985), .B0(n13837), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_984), .B1(n13837), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12738), .COUT(n12739), .S0(n158_adj_920), 
          .S1(n155_adj_919));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_5 (.A0(n155_adj_983), .B0(n13837), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_982), .B1(n13837), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12739), .COUT(n12740), .S0(n152_adj_918), 
          .S1(n149_adj_917));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_7 (.A0(n149_adj_981), .B0(n13837), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_980), .B1(n13837), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12740), .COUT(n12741), .S0(n146_adj_916), 
          .S1(n143_adj_915));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_9 (.A0(n143_adj_979), .B0(n13837), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_978), .B1(n13837), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12741), .COUT(n12742), .S0(n140_adj_914), 
          .S1(n137_adj_913));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_11 (.A0(n137_adj_977), .B0(n13837), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_976), .B1(n13837), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12742), .COUT(n12743), .S0(n134_adj_912), 
          .S1(n131_adj_911));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_13 (.A0(n131_adj_975), .B0(n13837), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_974), .B1(n13837), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12743), .COUT(n12744), .S0(n128_adj_910), 
          .S1(n125_adj_909));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_15 (.A0(n125_adj_973), .B0(n13837), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_972), .B1(n13837), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12744), .COUT(n12745), .S0(n122_adj_908), 
          .S1(n119_adj_907));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_17 (.A0(n119_adj_971), .B0(n13837), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_970), .B1(n13837), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12745), .COUT(n12746), .S0(n116_adj_906), 
          .S1(n113_adj_905));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_19 (.A0(n113_adj_969), .B0(n13837), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_968), .B1(n13837), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12746), .COUT(n12747), .S0(n110_adj_904), 
          .S1(n107_adj_903));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_21 (.A0(n107_adj_967), .B0(n13837), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_966), .B1(n13837), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12747), .COUT(n12748), .S0(n104_adj_902), 
          .S1(n101_adj_901));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_23 (.A0(n101_adj_965), .B0(n13837), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_964), .B1(n13837), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12748), .COUT(n12749), .S0(n98_adj_900), 
          .S1(n95_adj_899));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_25 (.A0(n95_adj_963), .B0(n13837), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_962), .B1(n13837), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12749), .COUT(n12750), .S0(n92_adj_898), 
          .S1(n89_adj_897));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_27 (.A0(n89_adj_961), .B0(n13837), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_960), .B1(n13837), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12750), .COUT(n12751), .S0(n86_adj_896), 
          .S1(n83_adj_895));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_29 (.A0(n83_adj_959), .B0(n13837), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_958), .B1(n13837), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12751), .COUT(n12752), .S0(n80_adj_894), 
          .S1(n77_adj_893));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_31 (.A0(n77_adj_957), .B0(n13837), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_956), .B1(n13837), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12752), .COUT(n12753), .S0(n74_adj_892), 
          .S1(n71_adj_891));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_475_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_475_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_475_add_4_33 (.A0(n1444), .B0(n13837), .C0(n71_adj_955), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12753), .S0(n68_adj_890));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_475_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_475_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_475_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_475_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13838), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12754), .S1(n161_adj_953));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_472_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_3 (.A0(n161_adj_1017), .B0(n13838), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1016), .B1(n13838), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12754), .COUT(n12755), .S0(n158_adj_952), 
          .S1(n155_adj_951));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_5 (.A0(n155_adj_1015), .B0(n13838), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1014), .B1(n13838), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12755), .COUT(n12756), .S0(n152_adj_950), 
          .S1(n149_adj_949));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_7 (.A0(n149_adj_1013), .B0(n13838), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1012), .B1(n13838), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12756), .COUT(n12757), .S0(n146_adj_948), 
          .S1(n143_adj_947));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_9 (.A0(n143_adj_1011), .B0(n13838), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1010), .B1(n13838), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12757), .COUT(n12758), .S0(n140_adj_946), 
          .S1(n137_adj_945));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_11 (.A0(n137_adj_1009), .B0(n13838), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1008), .B1(n13838), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12758), .COUT(n12759), .S0(n134_adj_944), 
          .S1(n131_adj_943));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_13 (.A0(n131_adj_1007), .B0(n13838), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1006), .B1(n13838), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12759), .COUT(n12760), .S0(n128_adj_942), 
          .S1(n125_adj_941));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_15 (.A0(n125_adj_1005), .B0(n13838), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1004), .B1(n13838), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12760), .COUT(n12761), .S0(n122_adj_940), 
          .S1(n119_adj_939));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_17 (.A0(n119_adj_1003), .B0(n13838), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1002), .B1(n13838), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12761), .COUT(n12762), .S0(n116_adj_938), 
          .S1(n113_adj_937));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_19 (.A0(n113_adj_1001), .B0(n13838), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1000), .B1(n13838), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12762), .COUT(n12763), .S0(n110_adj_936), 
          .S1(n107_adj_935));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_21 (.A0(n107_adj_999), .B0(n13838), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_998), .B1(n13838), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12763), .COUT(n12764), .S0(n104_adj_934), 
          .S1(n101_adj_933));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_23 (.A0(n101_adj_997), .B0(n13838), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_996), .B1(n13838), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12764), .COUT(n12765), .S0(n98_adj_932), 
          .S1(n95_adj_931));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_25 (.A0(n95_adj_995), .B0(n13838), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_994), .B1(n13838), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12765), .COUT(n12766), .S0(n92_adj_930), 
          .S1(n89_adj_929));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_27 (.A0(n89_adj_993), .B0(n13838), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_992), .B1(n13838), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12766), .COUT(n12767), .S0(n86_adj_928), 
          .S1(n83_adj_927));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_29 (.A0(n83_adj_991), .B0(n13838), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_990), .B1(n13838), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12767), .COUT(n12768), .S0(n80_adj_926), 
          .S1(n77_adj_925));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_31 (.A0(n77_adj_989), .B0(n13838), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_988), .B1(n13838), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12768), .COUT(n12769), .S0(n74_adj_924), 
          .S1(n71_adj_923));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_472_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_472_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_472_add_4_33 (.A0(n1444), .B0(n13838), .C0(n71_adj_987), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12769), .S0(n68_adj_922));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_472_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_472_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_472_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_472_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13838), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12770), .S1(n161_adj_985));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_469_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_3 (.A0(n161_adj_1049), .B0(n13838), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1048), .B1(n13838), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12770), .COUT(n12771), .S0(n158_adj_984), 
          .S1(n155_adj_983));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_5 (.A0(n155_adj_1047), .B0(n13838), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1046), .B1(n13838), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12771), .COUT(n12772), .S0(n152_adj_982), 
          .S1(n149_adj_981));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_7 (.A0(n149_adj_1045), .B0(n13838), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1044), .B1(n13838), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12772), .COUT(n12773), .S0(n146_adj_980), 
          .S1(n143_adj_979));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_9 (.A0(n143_adj_1043), .B0(n13838), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1042), .B1(n13838), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12773), .COUT(n12774), .S0(n140_adj_978), 
          .S1(n137_adj_977));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_11 (.A0(n137_adj_1041), .B0(n13838), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1040), .B1(n13838), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12774), .COUT(n12775), .S0(n134_adj_976), 
          .S1(n131_adj_975));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_13 (.A0(n131_adj_1039), .B0(n13838), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1038), .B1(n13838), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12775), .COUT(n12776), .S0(n128_adj_974), 
          .S1(n125_adj_973));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_15 (.A0(n125_adj_1037), .B0(n13838), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1036), .B1(n13838), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12776), .COUT(n12777), .S0(n122_adj_972), 
          .S1(n119_adj_971));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_17 (.A0(n119_adj_1035), .B0(n13838), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1034), .B1(n13838), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12777), .COUT(n12778), .S0(n116_adj_970), 
          .S1(n113_adj_969));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_19 (.A0(n113_adj_1033), .B0(n13838), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1032), .B1(n13838), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12778), .COUT(n12779), .S0(n110_adj_968), 
          .S1(n107_adj_967));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_21 (.A0(n107_adj_1031), .B0(n13838), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1030), .B1(n13838), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12779), .COUT(n12780), .S0(n104_adj_966), 
          .S1(n101_adj_965));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_23 (.A0(n101_adj_1029), .B0(n13838), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1028), .B1(n13838), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12780), .COUT(n12781), .S0(n98_adj_964), 
          .S1(n95_adj_963));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_25 (.A0(n95_adj_1027), .B0(n13838), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1026), .B1(n13838), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12781), .COUT(n12782), .S0(n92_adj_962), 
          .S1(n89_adj_961));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_27 (.A0(n89_adj_1025), .B0(n13838), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1024), .B1(n13838), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12782), .COUT(n12783), .S0(n86_adj_960), 
          .S1(n83_adj_959));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_29 (.A0(n83_adj_1023), .B0(n13838), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1022), .B1(n13838), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12783), .COUT(n12784), .S0(n80_adj_958), 
          .S1(n77_adj_957));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_31 (.A0(n77_adj_1021), .B0(n13838), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1020), .B1(n13838), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12784), .COUT(n12785), .S0(n74_adj_956), 
          .S1(n71_adj_955));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_469_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_469_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_469_add_4_33 (.A0(n1444), .B0(n13838), .C0(n71_adj_1019), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12785), .S0(n68_adj_954));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_469_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_469_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_469_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_469_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13839), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12786), .S1(n161_adj_1017));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_466_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_3 (.A0(n161_adj_1081), .B0(n13839), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1080), .B1(n13839), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12786), .COUT(n12787), .S0(n158_adj_1016), 
          .S1(n155_adj_1015));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_5 (.A0(n155_adj_1079), .B0(n13839), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1078), .B1(n13839), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12787), .COUT(n12788), .S0(n152_adj_1014), 
          .S1(n149_adj_1013));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_7 (.A0(n149_adj_1077), .B0(n13839), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1076), .B1(n13839), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12788), .COUT(n12789), .S0(n146_adj_1012), 
          .S1(n143_adj_1011));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_9 (.A0(n143_adj_1075), .B0(n13839), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1074), .B1(n13839), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12789), .COUT(n12790), .S0(n140_adj_1010), 
          .S1(n137_adj_1009));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_11 (.A0(n137_adj_1073), .B0(n13839), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1072), .B1(n13839), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12790), .COUT(n12791), .S0(n134_adj_1008), 
          .S1(n131_adj_1007));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_13 (.A0(n131_adj_1071), .B0(n13839), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1070), .B1(n13839), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12791), .COUT(n12792), .S0(n128_adj_1006), 
          .S1(n125_adj_1005));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_15 (.A0(n125_adj_1069), .B0(n13839), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1068), .B1(n13839), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12792), .COUT(n12793), .S0(n122_adj_1004), 
          .S1(n119_adj_1003));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_17 (.A0(n119_adj_1067), .B0(n13839), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1066), .B1(n13839), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12793), .COUT(n12794), .S0(n116_adj_1002), 
          .S1(n113_adj_1001));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_19 (.A0(n113_adj_1065), .B0(n13839), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1064), .B1(n13839), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12794), .COUT(n12795), .S0(n110_adj_1000), 
          .S1(n107_adj_999));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_21 (.A0(n107_adj_1063), .B0(n13839), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1062), .B1(n13839), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12795), .COUT(n12796), .S0(n104_adj_998), 
          .S1(n101_adj_997));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_23 (.A0(n101_adj_1061), .B0(n13839), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1060), .B1(n13839), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12796), .COUT(n12797), .S0(n98_adj_996), 
          .S1(n95_adj_995));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_25 (.A0(n95_adj_1059), .B0(n13839), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1058), .B1(n13839), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12797), .COUT(n12798), .S0(n92_adj_994), 
          .S1(n89_adj_993));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_27 (.A0(n89_adj_1057), .B0(n13839), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1056), .B1(n13839), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12798), .COUT(n12799), .S0(n86_adj_992), 
          .S1(n83_adj_991));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_29 (.A0(n83_adj_1055), .B0(n13839), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1054), .B1(n13839), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12799), .COUT(n12800), .S0(n80_adj_990), 
          .S1(n77_adj_989));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_31 (.A0(n77_adj_1053), .B0(n13839), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1052), .B1(n13839), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12800), .COUT(n12801), .S0(n74_adj_988), 
          .S1(n71_adj_987));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_466_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_466_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_466_add_4_33 (.A0(n1444), .B0(n13839), .C0(n71_adj_1051), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12801), .S0(n68_adj_986));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_466_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_466_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_466_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_466_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13839), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12802), .S1(n161_adj_1049));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_463_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_3 (.A0(n161_adj_1113), .B0(n13839), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1112), .B1(n13839), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12802), .COUT(n12803), .S0(n158_adj_1048), 
          .S1(n155_adj_1047));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_5 (.A0(n155_adj_1111), .B0(n13839), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1110), .B1(n13839), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12803), .COUT(n12804), .S0(n152_adj_1046), 
          .S1(n149_adj_1045));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_7 (.A0(n149_adj_1109), .B0(n13839), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1108), .B1(n13839), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12804), .COUT(n12805), .S0(n146_adj_1044), 
          .S1(n143_adj_1043));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_9 (.A0(n143_adj_1107), .B0(n13839), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1106), .B1(n13839), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12805), .COUT(n12806), .S0(n140_adj_1042), 
          .S1(n137_adj_1041));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_11 (.A0(n137_adj_1105), .B0(n13839), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1104), .B1(n13839), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12806), .COUT(n12807), .S0(n134_adj_1040), 
          .S1(n131_adj_1039));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_13 (.A0(n131_adj_1103), .B0(n13839), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1102), .B1(n13839), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12807), .COUT(n12808), .S0(n128_adj_1038), 
          .S1(n125_adj_1037));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_15 (.A0(n125_adj_1101), .B0(n13839), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1100), .B1(n13839), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12808), .COUT(n12809), .S0(n122_adj_1036), 
          .S1(n119_adj_1035));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_17 (.A0(n119_adj_1099), .B0(n13839), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1098), .B1(n13839), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12809), .COUT(n12810), .S0(n116_adj_1034), 
          .S1(n113_adj_1033));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_19 (.A0(n113_adj_1097), .B0(n13839), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1096), .B1(n13839), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12810), .COUT(n12811), .S0(n110_adj_1032), 
          .S1(n107_adj_1031));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_21 (.A0(n107_adj_1095), .B0(n13839), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1094), .B1(n13839), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12811), .COUT(n12812), .S0(n104_adj_1030), 
          .S1(n101_adj_1029));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_23 (.A0(n101_adj_1093), .B0(n13839), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1092), .B1(n13839), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12812), .COUT(n12813), .S0(n98_adj_1028), 
          .S1(n95_adj_1027));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_25 (.A0(n95_adj_1091), .B0(n13839), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1090), .B1(n13839), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12813), .COUT(n12814), .S0(n92_adj_1026), 
          .S1(n89_adj_1025));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_27 (.A0(n89_adj_1089), .B0(n13839), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1088), .B1(n13839), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12814), .COUT(n12815), .S0(n86_adj_1024), 
          .S1(n83_adj_1023));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_29 (.A0(n83_adj_1087), .B0(n13839), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1086), .B1(n13839), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12815), .COUT(n12816), .S0(n80_adj_1022), 
          .S1(n77_adj_1021));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_31 (.A0(n77_adj_1085), .B0(n13839), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1084), .B1(n13839), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12816), .COUT(n12817), .S0(n74_adj_1020), 
          .S1(n71_adj_1019));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_463_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_463_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_463_add_4_33 (.A0(n1444), .B0(n13839), .C0(n71_adj_1083), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12817), .S0(n68_adj_1018));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_463_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_463_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_463_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_463_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13840), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12818), .S1(n161_adj_1081));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_460_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_3 (.A0(n161_adj_1145), .B0(n13840), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1144), .B1(n13840), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12818), .COUT(n12819), .S0(n158_adj_1080), 
          .S1(n155_adj_1079));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_5 (.A0(n155_adj_1143), .B0(n13840), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1142), .B1(n13840), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12819), .COUT(n12820), .S0(n152_adj_1078), 
          .S1(n149_adj_1077));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_7 (.A0(n149_adj_1141), .B0(n13840), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1140), .B1(n13840), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12820), .COUT(n12821), .S0(n146_adj_1076), 
          .S1(n143_adj_1075));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_9 (.A0(n143_adj_1139), .B0(n13840), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1138), .B1(n13840), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12821), .COUT(n12822), .S0(n140_adj_1074), 
          .S1(n137_adj_1073));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_11 (.A0(n137_adj_1137), .B0(n13840), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1136), .B1(n13840), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12822), .COUT(n12823), .S0(n134_adj_1072), 
          .S1(n131_adj_1071));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_13 (.A0(n131_adj_1135), .B0(n13840), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1134), .B1(n13840), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12823), .COUT(n12824), .S0(n128_adj_1070), 
          .S1(n125_adj_1069));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_15 (.A0(n125_adj_1133), .B0(n13840), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1132), .B1(n13840), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12824), .COUT(n12825), .S0(n122_adj_1068), 
          .S1(n119_adj_1067));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_17 (.A0(n119_adj_1131), .B0(n13840), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1130), .B1(n13840), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12825), .COUT(n12826), .S0(n116_adj_1066), 
          .S1(n113_adj_1065));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_19 (.A0(n113_adj_1129), .B0(n13840), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1128), .B1(n13840), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12826), .COUT(n12827), .S0(n110_adj_1064), 
          .S1(n107_adj_1063));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_21 (.A0(n107_adj_1127), .B0(n13840), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1126), .B1(n13840), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12827), .COUT(n12828), .S0(n104_adj_1062), 
          .S1(n101_adj_1061));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_23 (.A0(n101_adj_1125), .B0(n13840), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1124), .B1(n13840), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12828), .COUT(n12829), .S0(n98_adj_1060), 
          .S1(n95_adj_1059));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_25 (.A0(n95_adj_1123), .B0(n13840), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1122), .B1(n13840), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12829), .COUT(n12830), .S0(n92_adj_1058), 
          .S1(n89_adj_1057));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_27 (.A0(n89_adj_1121), .B0(n13840), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1120), .B1(n13840), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12830), .COUT(n12831), .S0(n86_adj_1056), 
          .S1(n83_adj_1055));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_29 (.A0(n83_adj_1119), .B0(n13840), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1118), .B1(n13840), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12831), .COUT(n12832), .S0(n80_adj_1054), 
          .S1(n77_adj_1053));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_31 (.A0(n77_adj_1117), .B0(n13840), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1116), .B1(n13840), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12832), .COUT(n12833), .S0(n74_adj_1052), 
          .S1(n71_adj_1051));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_460_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_460_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_460_add_4_33 (.A0(n1444), .B0(n13840), .C0(n71_adj_1115), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12833), .S0(n68_adj_1050));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_460_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_460_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_460_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_460_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13840), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n12834), .S1(n161_adj_1113));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_457_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_3 (.A0(n161_adj_1177), .B0(n13840), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1176), .B1(n13840), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n12834), .COUT(n12835), .S0(n158_adj_1112), 
          .S1(n155_adj_1111));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_5 (.A0(n155_adj_1175), .B0(n13840), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1174), .B1(n13840), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n12835), .COUT(n12836), .S0(n152_adj_1110), 
          .S1(n149_adj_1109));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_7 (.A0(n149_adj_1173), .B0(n13840), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1172), .B1(n13840), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n12836), .COUT(n12837), .S0(n146_adj_1108), 
          .S1(n143_adj_1107));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_9 (.A0(n143_adj_1171), .B0(n13840), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1170), .B1(n13840), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n12837), .COUT(n12838), .S0(n140_adj_1106), 
          .S1(n137_adj_1105));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_11 (.A0(n137_adj_1169), .B0(n13840), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1168), .B1(n13840), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n12838), .COUT(n12839), .S0(n134_adj_1104), 
          .S1(n131_adj_1103));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_13 (.A0(n131_adj_1167), .B0(n13840), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1166), .B1(n13840), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n12839), .COUT(n12840), .S0(n128_adj_1102), 
          .S1(n125_adj_1101));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_15 (.A0(n125_adj_1165), .B0(n13840), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1164), .B1(n13840), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n12840), .COUT(n12841), .S0(n122_adj_1100), 
          .S1(n119_adj_1099));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_17 (.A0(n119_adj_1163), .B0(n13840), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1162), .B1(n13840), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n12841), .COUT(n12842), .S0(n116_adj_1098), 
          .S1(n113_adj_1097));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_19 (.A0(n113_adj_1161), .B0(n13840), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1160), .B1(n13840), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n12842), .COUT(n12843), .S0(n110_adj_1096), 
          .S1(n107_adj_1095));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_21 (.A0(n107_adj_1159), .B0(n13840), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1158), .B1(n13840), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n12843), .COUT(n12844), .S0(n104_adj_1094), 
          .S1(n101_adj_1093));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_23 (.A0(n101_adj_1157), .B0(n13840), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1156), .B1(n13840), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n12844), .COUT(n12845), .S0(n98_adj_1092), 
          .S1(n95_adj_1091));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_25 (.A0(n95_adj_1155), .B0(n13840), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1154), .B1(n13840), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n12845), .COUT(n12846), .S0(n92_adj_1090), 
          .S1(n89_adj_1089));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_27 (.A0(n89_adj_1153), .B0(n13840), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1152), .B1(n13840), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n12846), .COUT(n12847), .S0(n86_adj_1088), 
          .S1(n83_adj_1087));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_29 (.A0(n83_adj_1151), .B0(n13840), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1150), .B1(n13840), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n12847), .COUT(n12848), .S0(n80_adj_1086), 
          .S1(n77_adj_1085));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_31 (.A0(n77_adj_1149), .B0(n13840), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1148), .B1(n13840), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n12848), .COUT(n12849), .S0(n74_adj_1084), 
          .S1(n71_adj_1083));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_457_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_457_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_457_add_4_33 (.A0(n1444), .B0(n13840), .C0(n71_adj_1147), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12849), .S0(n68_adj_1082));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_457_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_457_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_457_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_457_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[1]), .B1(det_q4_28[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12850), .S1(n161_adj_1145));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_454_add_4_1.INIT1 = 16'h999a;
    defparam _add_1_454_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_3 (.A0(det_q4_28[2]), .B0(n1441), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[3]), .B1(n1440), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12850), .COUT(n12851), .S0(n158_adj_1144), 
          .S1(n155_adj_1143));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_3.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_5 (.A0(det_q4_28[4]), .B0(n1439), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[5]), .B1(n1438), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12851), .COUT(n12852), .S0(n152_adj_1142), 
          .S1(n149_adj_1141));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_5.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_5.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_7 (.A0(det_q4_28[6]), .B0(n1437), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[7]), .B1(n1436), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12852), .COUT(n12853), .S0(n146_adj_1140), 
          .S1(n143_adj_1139));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_7.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_7.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_9 (.A0(det_q4_28[8]), .B0(n1435), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[9]), .B1(n1434), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12853), .COUT(n12854), .S0(n140_adj_1138), 
          .S1(n137_adj_1137));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_9.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_9.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_11 (.A0(det_q4_28[10]), .B0(n1433), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[11]), .B1(n1432), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12854), .COUT(n12855), .S0(n134_adj_1136), 
          .S1(n131_adj_1135));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_11.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_11.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_13 (.A0(det_q4_28[12]), .B0(n1431), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[13]), .B1(n1430), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12855), .COUT(n12856), .S0(n128_adj_1134), 
          .S1(n125_adj_1133));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_13.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_13.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_15 (.A0(det_q4_28[14]), .B0(n1429), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[15]), .B1(n1428), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12856), .COUT(n12857), .S0(n122_adj_1132), 
          .S1(n119_adj_1131));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_15.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_15.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_17 (.A0(det_q4_28[16]), .B0(n1427), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[17]), .B1(n1426), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12857), .COUT(n12858), .S0(n116_adj_1130), 
          .S1(n113_adj_1129));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_17.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_17.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_19 (.A0(det_q4_28[18]), .B0(n1425), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[19]), .B1(n1424), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12858), .COUT(n12859), .S0(n110_adj_1128), 
          .S1(n107_adj_1127));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_19.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_19.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_21 (.A0(det_q4_28[20]), .B0(n1423), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[21]), .B1(n1422), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12859), .COUT(n12860), .S0(n104_adj_1126), 
          .S1(n101_adj_1125));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_21.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_21.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_23 (.A0(det_q4_28[22]), .B0(n1421), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[23]), .B1(n1420), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12860), .COUT(n12861), .S0(n98_adj_1124), 
          .S1(n95_adj_1123));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_23.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_23.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_25 (.A0(det_q4_28[24]), .B0(n1419), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[25]), .B1(n1418), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12861), .COUT(n12862), .S0(n92_adj_1122), 
          .S1(n89_adj_1121));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_25.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_25.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_27 (.A0(det_q4_28[26]), .B0(n1417), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[27]), .B1(n1416), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12862), .COUT(n12863), .S0(n86_adj_1120), 
          .S1(n83_adj_1119));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_27.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_27.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_29 (.A0(det_q4_28[28]), .B0(n1415), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[29]), .B1(n1414), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12863), .COUT(n12864), .S0(n80_adj_1118), 
          .S1(n77_adj_1117));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_29.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_29.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_31 (.A0(det_q4_28[30]), .B0(n1413), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[31]), .B1(n1412), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12864), .COUT(n12865), .S0(n74_adj_1116), 
          .S1(n71_adj_1115));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_31.INIT0 = 16'h666a;
    defparam _add_1_454_add_4_31.INIT1 = 16'h666a;
    defparam _add_1_454_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_454_add_4_33 (.A0(n1411), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12865), .S0(n68_adj_1114));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_454_add_4_33.INIT0 = 16'haaa0;
    defparam _add_1_454_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_454_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_454_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n1475), .B1(det_q4_28[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12866), .S1(n161_adj_1177));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_451_add_4_1.INIT1 = 16'h999a;
    defparam _add_1_451_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_3 (.A0(n1474), .B0(n1441), .C0(GND_net), .D0(VCC_net), 
          .A1(n1473), .B1(n1440), .C1(GND_net), .D1(VCC_net), .CIN(n12866), 
          .COUT(n12867), .S0(n158_adj_1176), .S1(n155_adj_1175));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_3.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_5 (.A0(n1472), .B0(n1439), .C0(GND_net), .D0(VCC_net), 
          .A1(n1471), .B1(n1438), .C1(GND_net), .D1(VCC_net), .CIN(n12867), 
          .COUT(n12868), .S0(n152_adj_1174), .S1(n149_adj_1173));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_5.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_5.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_7 (.A0(n1470), .B0(n1437), .C0(GND_net), .D0(VCC_net), 
          .A1(n1469), .B1(n1436), .C1(GND_net), .D1(VCC_net), .CIN(n12868), 
          .COUT(n12869), .S0(n146_adj_1172), .S1(n143_adj_1171));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_7.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_7.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_9 (.A0(n1468), .B0(n1435), .C0(GND_net), .D0(VCC_net), 
          .A1(n1467), .B1(n1434), .C1(GND_net), .D1(VCC_net), .CIN(n12869), 
          .COUT(n12870), .S0(n140_adj_1170), .S1(n137_adj_1169));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_9.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_9.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_11 (.A0(n1466), .B0(n1433), .C0(GND_net), .D0(VCC_net), 
          .A1(n1465), .B1(n1432), .C1(GND_net), .D1(VCC_net), .CIN(n12870), 
          .COUT(n12871), .S0(n134_adj_1168), .S1(n131_adj_1167));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_11.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_11.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_13 (.A0(n1464), .B0(n1431), .C0(GND_net), .D0(VCC_net), 
          .A1(n1463), .B1(n1430), .C1(GND_net), .D1(VCC_net), .CIN(n12871), 
          .COUT(n12872), .S0(n128_adj_1166), .S1(n125_adj_1165));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_13.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_13.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_15 (.A0(n1462), .B0(n1429), .C0(GND_net), .D0(VCC_net), 
          .A1(n1461), .B1(n1428), .C1(GND_net), .D1(VCC_net), .CIN(n12872), 
          .COUT(n12873), .S0(n122_adj_1164), .S1(n119_adj_1163));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_15.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_15.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_17 (.A0(n1460), .B0(n1427), .C0(GND_net), .D0(VCC_net), 
          .A1(n1459), .B1(n1426), .C1(GND_net), .D1(VCC_net), .CIN(n12873), 
          .COUT(n12874), .S0(n116_adj_1162), .S1(n113_adj_1161));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_17.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_17.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_19 (.A0(n1458), .B0(n1425), .C0(GND_net), .D0(VCC_net), 
          .A1(n1457), .B1(n1424), .C1(GND_net), .D1(VCC_net), .CIN(n12874), 
          .COUT(n12875), .S0(n110_adj_1160), .S1(n107_adj_1159));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_19.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_19.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_21 (.A0(n1456), .B0(n1423), .C0(GND_net), .D0(VCC_net), 
          .A1(n1455), .B1(n1422), .C1(GND_net), .D1(VCC_net), .CIN(n12875), 
          .COUT(n12876), .S0(n104_adj_1158), .S1(n101_adj_1157));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_21.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_21.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_23 (.A0(n1454), .B0(n1421), .C0(GND_net), .D0(VCC_net), 
          .A1(n1453), .B1(n1420), .C1(GND_net), .D1(VCC_net), .CIN(n12876), 
          .COUT(n12877), .S0(n98_adj_1156), .S1(n95_adj_1155));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_23.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_23.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_25 (.A0(n1452), .B0(n1419), .C0(GND_net), .D0(VCC_net), 
          .A1(n1451), .B1(n1418), .C1(GND_net), .D1(VCC_net), .CIN(n12877), 
          .COUT(n12878), .S0(n92_adj_1154), .S1(n89_adj_1153));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_25.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_25.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_27 (.A0(n1450), .B0(n1417), .C0(GND_net), .D0(VCC_net), 
          .A1(n1449), .B1(n1416), .C1(GND_net), .D1(VCC_net), .CIN(n12878), 
          .COUT(n12879), .S0(n86_adj_1152), .S1(n83_adj_1151));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_27.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_27.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_29 (.A0(n1448), .B0(n1415), .C0(GND_net), .D0(VCC_net), 
          .A1(n1447), .B1(n1414), .C1(GND_net), .D1(VCC_net), .CIN(n12879), 
          .COUT(n12880), .S0(n80_adj_1150), .S1(n77_adj_1149));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_29.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_29.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_31 (.A0(n1446), .B0(n1413), .C0(GND_net), .D0(VCC_net), 
          .A1(n1445), .B1(n1412), .C1(GND_net), .D1(VCC_net), .CIN(n12880), 
          .COUT(n12881), .S0(n74_adj_1148), .S1(n71_adj_1147));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_31.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_31.INIT1 = 16'h666a;
    defparam _add_1_451_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_451_add_4_33 (.A0(n1444), .B0(n1411), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12881), 
          .S0(n68_adj_1146));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_451_add_4_33.INIT0 = 16'h666a;
    defparam _add_1_451_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_451_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_451_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n1846), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12885));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_448_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_448_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_3 (.A0(det_q4_28[0]), .B0(n1846), .C0(n161_adj_1493), 
          .D0(n2380), .A1(n161_adj_1587), .B1(n1846), .C1(n158_adj_1492), 
          .D1(n2379), .CIN(n12885), .COUT(n12886), .S0(n161_adj_1208), 
          .S1(n158_adj_1207));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_3.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_3.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_5 (.A0(n158_adj_1586), .B0(n1846), .C0(n155_adj_1491), 
          .D0(n2378), .A1(n155_adj_1585), .B1(n1846), .C1(n152_adj_1490), 
          .D1(n2377), .CIN(n12886), .COUT(n12887), .S0(n155_adj_1206), 
          .S1(n152_adj_1205));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_5.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_5.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_7 (.A0(n152_adj_1584), .B0(n1846), .C0(n149_adj_1489), 
          .D0(n2376), .A1(n149_adj_1583), .B1(n1846), .C1(n146_adj_1488), 
          .D1(n2375), .CIN(n12887), .COUT(n12888), .S0(n149_adj_1204), 
          .S1(n146_adj_1203));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_7.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_7.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_9 (.A0(n146_adj_1582), .B0(n1846), .C0(n143_adj_1487), 
          .D0(n2374), .A1(n143_adj_1581), .B1(n1846), .C1(n140_adj_1486), 
          .D1(n2373), .CIN(n12888), .COUT(n12889), .S0(n143_adj_1202), 
          .S1(n140_adj_1201));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_9.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_9.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_11 (.A0(n140_adj_1580), .B0(n1846), .C0(n137_adj_1485), 
          .D0(n2372), .A1(n137_adj_1579), .B1(n1846), .C1(n134_adj_1484), 
          .D1(n2371), .CIN(n12889), .COUT(n12890), .S0(n137_adj_1200), 
          .S1(n134_adj_1199));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_11.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_11.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_13 (.A0(n134_adj_1578), .B0(n1846), .C0(n131_adj_1483), 
          .D0(n2370), .A1(n131_adj_1577), .B1(n1846), .C1(n128_adj_1482), 
          .D1(n2369), .CIN(n12890), .COUT(n12891), .S0(n131_adj_1198), 
          .S1(n128_adj_1197));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_13.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_13.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_15 (.A0(n128_adj_1576), .B0(n1846), .C0(n125_adj_1481), 
          .D0(n2368), .A1(n125_adj_1575), .B1(n1846), .C1(n122_adj_1480), 
          .D1(n2367), .CIN(n12891), .COUT(n12892), .S0(n125_adj_1196), 
          .S1(n122_adj_1195));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_15.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_15.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_17 (.A0(n122_adj_1574), .B0(n1846), .C0(n119_adj_1479), 
          .D0(n2366), .A1(n119_adj_1573), .B1(n1846), .C1(n116_adj_1478), 
          .D1(n2365), .CIN(n12892), .COUT(n12893), .S0(n119_adj_1194), 
          .S1(n116_adj_1193));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_17.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_17.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_19 (.A0(n116_adj_1572), .B0(n1846), .C0(n113_adj_1477), 
          .D0(n2364), .A1(n113_adj_1571), .B1(n1846), .C1(n110_adj_1476), 
          .D1(n2363), .CIN(n12893), .COUT(n12894), .S0(n113_adj_1192), 
          .S1(n110_adj_1191));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_19.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_19.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_21 (.A0(n110_adj_1570), .B0(n1846), .C0(n107_adj_1475), 
          .D0(n2362), .A1(n107_adj_1569), .B1(n1846), .C1(n104_adj_1474), 
          .D1(n2361), .CIN(n12894), .COUT(n12895), .S0(n107_adj_1190), 
          .S1(n104_adj_1189));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_21.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_21.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_23 (.A0(n104_adj_1568), .B0(n1846), .C0(n101_adj_1473), 
          .D0(n2360), .A1(n101_adj_1567), .B1(n1846), .C1(n98_adj_1472), 
          .D1(n2359), .CIN(n12895), .COUT(n12896), .S0(n101_adj_1188), 
          .S1(n98_adj_1187));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_23.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_23.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_25 (.A0(n98_adj_1566), .B0(n1846), .C0(n95_adj_1471), 
          .D0(n2358), .A1(n95_adj_1565), .B1(n1846), .C1(n92_adj_1470), 
          .D1(n2357), .CIN(n12896), .COUT(n12897), .S0(n95_adj_1186), 
          .S1(n92_adj_1185));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_25.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_25.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_27 (.A0(n92_adj_1564), .B0(n1846), .C0(n89_adj_1469), 
          .D0(n2356), .A1(n89_adj_1563), .B1(n1846), .C1(n86_adj_1468), 
          .D1(n2355), .CIN(n12897), .COUT(n12898), .S0(n89_adj_1184), 
          .S1(n86_adj_1183));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_27.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_27.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_29 (.A0(n86_adj_1562), .B0(n1846), .C0(n83_adj_1467), 
          .D0(n2354), .A1(n83_adj_1561), .B1(n1846), .C1(n80_adj_1466), 
          .D1(n2353), .CIN(n12898), .COUT(n12899), .S0(n83_adj_1182), 
          .S1(n80_adj_1181));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_29.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_29.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_31 (.A0(n80_adj_1560), .B0(n1846), .C0(n77_adj_1465), 
          .D0(n2352), .A1(n77_adj_1559), .B1(n1846), .C1(n74_adj_1464), 
          .D1(n2351), .CIN(n12899), .COUT(n12900), .S0(n77_adj_1180), 
          .S1(n74_adj_1179));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_31.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_31.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_448_add_4_33 (.A0(n74_adj_1558), .B0(n1846), .C0(n71_adj_1463), 
          .D0(n2350), .A1(n71_adj_1557), .B1(n1846), .C1(n68_adj_1462), 
          .D1(n2349), .CIN(n12900), .S0(n71_adj_1178), .S1(n2382));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_448_add_4_33.INIT0 = 16'h74b8;
    defparam _add_1_448_add_4_33.INIT1 = 16'h74b8;
    defparam _add_1_448_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_448_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[1]), .B1(det_q4_28[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12902), .S1(n1475));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_445_add_4_1.INIT1 = 16'h6665;
    defparam _add_1_445_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_3 (.A0(det_q4_28[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12902), .COUT(n12903), .S0(n1474), .S1(n1473));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_5 (.A0(det_q4_28[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12903), .COUT(n12904), .S0(n1472), .S1(n1471));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_7 (.A0(det_q4_28[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12904), .COUT(n12905), .S0(n1470), .S1(n1469));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_9 (.A0(det_q4_28[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12905), .COUT(n12906), .S0(n1468), .S1(n1467));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_11 (.A0(det_q4_28[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12906), .COUT(n12907), .S0(n1466), .S1(n1465));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_13 (.A0(det_q4_28[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12907), .COUT(n12908), .S0(n1464), .S1(n1463));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_13.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_15 (.A0(det_q4_28[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12908), .COUT(n12909), .S0(n1462), .S1(n1461));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_15.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_15.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_17 (.A0(det_q4_28[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12909), .COUT(n12910), .S0(n1460), .S1(n1459));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_17.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_17.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_19 (.A0(det_q4_28[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12910), .COUT(n12911), .S0(n1458), .S1(n1457));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_19.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_19.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_21 (.A0(det_q4_28[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12911), .COUT(n12912), .S0(n1456), .S1(n1455));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_21.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_21.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_23 (.A0(det_q4_28[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12912), .COUT(n12913), .S0(n1454), .S1(n1453));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_23.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_23.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_25 (.A0(det_q4_28[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12913), .COUT(n12914), .S0(n1452), .S1(n1451));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_25.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_25.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_27 (.A0(det_q4_28[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12914), .COUT(n12915), .S0(n1450), .S1(n1449));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_27.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_27.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_29 (.A0(det_q4_28[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12915), .COUT(n12916), .S0(n1448), .S1(n1447));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_29.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_29.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_31 (.A0(det_q4_28[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12916), .COUT(n12917), .S0(n1446), .S1(n1445));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_31.INIT0 = 16'h5555;
    defparam _add_1_445_add_4_31.INIT1 = 16'h5555;
    defparam _add_1_445_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_445_add_4_33 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12917), .S0(n1444));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_445_add_4_33.INIT0 = 16'hffff;
    defparam _add_1_445_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_445_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_445_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_2 (.A0(prod_d[15]), .B0(prod_d[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12918));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_442_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_4 (.A0(prod_d[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12918), .COUT(n12919));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_6 (.A0(prod_d[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12919), .COUT(n12920));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_8 (.A0(prod_d[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12920), .COUT(n12921));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_10 (.A0(prod_d[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12921), .COUT(n12922));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_12 (.A0(prod_d[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12922), .COUT(n12923));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_14 (.A0(prod_d[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12923), .COUT(n12924));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_16 (.A0(prod_d[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12924), .COUT(n12925));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_18 (.A0(prod_d[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12925), .COUT(n12926), .S0(d_inv_15__N_49[32]), 
          .S1(d_inv_15__N_49[33]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_20 (.A0(prod_d[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12926), .COUT(n12927), .S0(d_inv_15__N_49[34]), 
          .S1(d_inv_15__N_49[35]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_22 (.A0(prod_d[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12927), .COUT(n12928), .S0(d_inv_15__N_49[36]), 
          .S1(d_inv_15__N_49[37]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_24 (.A0(prod_d[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12928), .COUT(n12929), .S0(d_inv_15__N_49[38]), 
          .S1(d_inv_15__N_49[39]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_26 (.A0(prod_d[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12929), .COUT(n12930), .S0(d_inv_15__N_49[40]), 
          .S1(d_inv_15__N_49[41]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_28 (.A0(prod_d[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12930), .COUT(n12931), .S0(d_inv_15__N_49[42]), 
          .S1(d_inv_15__N_49[43]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_30 (.A0(prod_d[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12931), .COUT(n12932), .S0(d_inv_15__N_49[44]), 
          .S1(d_inv_15__N_49[45]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_442_add_4_32 (.A0(prod_d[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12932), .S0(d_inv_15__N_49[46]), .S1(d_inv_15__N_49[47]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_442_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_442_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_442_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_442_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_2 (.A0(prod_a[15]), .B0(prod_a[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12934));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_439_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_4 (.A0(prod_a[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12934), .COUT(n12935));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_6 (.A0(prod_a[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12935), .COUT(n12936));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_8 (.A0(prod_a[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12936), .COUT(n12937));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_10 (.A0(prod_a[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12937), .COUT(n12938));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_12 (.A0(prod_a[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12938), .COUT(n12939));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_14 (.A0(prod_a[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12939), .COUT(n12940));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_16 (.A0(prod_a[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12940), .COUT(n12941));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_18 (.A0(prod_a[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12941), .COUT(n12942), .S0(a_inv_15__N_1[32]), 
          .S1(a_inv_15__N_1[33]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_20 (.A0(prod_a[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12942), .COUT(n12943), .S0(a_inv_15__N_1[34]), 
          .S1(a_inv_15__N_1[35]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_22 (.A0(prod_a[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12943), .COUT(n12944), .S0(a_inv_15__N_1[36]), 
          .S1(a_inv_15__N_1[37]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_24 (.A0(prod_a[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12944), .COUT(n12945), .S0(a_inv_15__N_1[38]), 
          .S1(a_inv_15__N_1[39]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_26 (.A0(prod_a[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12945), .COUT(n12946), .S0(a_inv_15__N_1[40]), 
          .S1(a_inv_15__N_1[41]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_28 (.A0(prod_a[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12946), .COUT(n12947), .S0(a_inv_15__N_1[42]), 
          .S1(a_inv_15__N_1[43]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_30 (.A0(prod_a[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12947), .COUT(n12948), .S0(a_inv_15__N_1[44]), 
          .S1(a_inv_15__N_1[45]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_439_add_4_32 (.A0(prod_a[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12948), .S0(a_inv_15__N_1[46]), .S1(a_inv_15__N_1[47]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_439_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_439_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_439_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_439_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_2 (.A0(prod_b[15]), .B0(prod_b[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12950));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_436_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_4 (.A0(prod_b[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12950), .COUT(n12951));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_6 (.A0(prod_b[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12951), .COUT(n12952));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_8 (.A0(prod_b[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12952), .COUT(n12953));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_10 (.A0(prod_b[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12953), .COUT(n12954));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_12 (.A0(prod_b[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12954), .COUT(n12955));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_14 (.A0(prod_b[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12955), .COUT(n12956));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_16 (.A0(prod_b[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12956), .COUT(n12957));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_18 (.A0(prod_b[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12957), .COUT(n12958), .S0(b_inv_15__N_17[32]), 
          .S1(b_inv_15__N_17[33]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_20 (.A0(prod_b[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12958), .COUT(n12959), .S0(b_inv_15__N_17[34]), 
          .S1(b_inv_15__N_17[35]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_22 (.A0(prod_b[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12959), .COUT(n12960), .S0(b_inv_15__N_17[36]), 
          .S1(b_inv_15__N_17[37]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_24 (.A0(prod_b[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12960), .COUT(n12961), .S0(b_inv_15__N_17[38]), 
          .S1(b_inv_15__N_17[39]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_26 (.A0(prod_b[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12961), .COUT(n12962), .S0(b_inv_15__N_17[40]), 
          .S1(b_inv_15__N_17[41]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_28 (.A0(prod_b[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12962), .COUT(n12963), .S0(b_inv_15__N_17[42]), 
          .S1(b_inv_15__N_17[43]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_30 (.A0(prod_b[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12963), .COUT(n12964), .S0(b_inv_15__N_17[44]), 
          .S1(b_inv_15__N_17[45]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_436_add_4_32 (.A0(prod_b[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12964), .S0(b_inv_15__N_17[46]), .S1(b_inv_15__N_17[47]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam _add_1_436_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_436_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_436_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_436_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_346), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12966));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_433_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_345), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_344), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12966), .COUT(n12967));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_343), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_342), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12967), .COUT(n12968));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_341), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_340), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12968), .COUT(n12969));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_339), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_338), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12969), .COUT(n12970));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_337), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_336), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12970), .COUT(n12971));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_335), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_334), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12971), .COUT(n12972));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_333), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_332), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12972), .COUT(n12973));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_331), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_330), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12973), .COUT(n12974));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_329), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_328), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12974), .COUT(n12975));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_327), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_326), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12975), .COUT(n12976));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_325), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_324), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12976), .COUT(n12977));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_323), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_322), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12977), .COUT(n12978));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_321), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_320), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12978), .COUT(n12979));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_319), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_318), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12979), .COUT(n12980));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_433_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_433_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_317), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_316), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12980), .S1(n68_adj_1209));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_433_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_433_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_433_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_433_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2449), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12985));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_430_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_430_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_3 (.A0(det_q4_28[0]), .B0(n2449), .C0(n161_adj_1272), 
          .D0(n1475), .A1(n161_adj_1303), .B1(n2449), .C1(n158_adj_1271), 
          .D1(n1474), .CIN(n12985), .COUT(n12986), .S0(n161_adj_1240), 
          .S1(n158_adj_1239));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_5 (.A0(n158_adj_1302), .B0(n2449), .C0(n155_adj_1270), 
          .D0(n1473), .A1(n155_adj_1301), .B1(n2449), .C1(n152_adj_1269), 
          .D1(n1472), .CIN(n12986), .COUT(n12987), .S0(n155_adj_1238), 
          .S1(n152_adj_1237));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_7 (.A0(n152_adj_1300), .B0(n2449), .C0(n149_adj_1268), 
          .D0(n1471), .A1(n149_adj_1299), .B1(n2449), .C1(n146_adj_1267), 
          .D1(n1470), .CIN(n12987), .COUT(n12988), .S0(n149_adj_1236), 
          .S1(n146_adj_1235));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_9 (.A0(n146_adj_1298), .B0(n2449), .C0(n143_adj_1266), 
          .D0(n1469), .A1(n143_adj_1297), .B1(n2449), .C1(n140_adj_1265), 
          .D1(n1468), .CIN(n12988), .COUT(n12989), .S0(n143_adj_1234), 
          .S1(n140_adj_1233));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_11 (.A0(n140_adj_1296), .B0(n2449), .C0(n137_adj_1264), 
          .D0(n1467), .A1(n137_adj_1295), .B1(n2449), .C1(n134_adj_1263), 
          .D1(n1466), .CIN(n12989), .COUT(n12990), .S0(n137_adj_1232), 
          .S1(n134_adj_1231));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_13 (.A0(n134_adj_1294), .B0(n2449), .C0(n131_adj_1262), 
          .D0(n1465), .A1(n131_adj_1293), .B1(n2449), .C1(n128_adj_1261), 
          .D1(n1464), .CIN(n12990), .COUT(n12991), .S0(n131_adj_1230), 
          .S1(n128_adj_1229));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_15 (.A0(n128_adj_1292), .B0(n2449), .C0(n125_adj_1260), 
          .D0(n1463), .A1(n125_adj_1291), .B1(n2449), .C1(n122_adj_1259), 
          .D1(n1462), .CIN(n12991), .COUT(n12992), .S0(n125_adj_1228), 
          .S1(n122_adj_1227));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_17 (.A0(n122_adj_1290), .B0(n2449), .C0(n119_adj_1258), 
          .D0(n1461), .A1(n119_adj_1289), .B1(n2449), .C1(n116_adj_1257), 
          .D1(n1460), .CIN(n12992), .COUT(n12993), .S0(n119_adj_1226), 
          .S1(n116_adj_1225));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_19 (.A0(n116_adj_1288), .B0(n2449), .C0(n113_adj_1256), 
          .D0(n1459), .A1(n113_adj_1287), .B1(n2449), .C1(n110_adj_1255), 
          .D1(n1458), .CIN(n12993), .COUT(n12994), .S0(n113_adj_1224), 
          .S1(n110_adj_1223));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_21 (.A0(n110_adj_1286), .B0(n2449), .C0(n107_adj_1254), 
          .D0(n1457), .A1(n107_adj_1285), .B1(n2449), .C1(n104_adj_1253), 
          .D1(n1456), .CIN(n12994), .COUT(n12995), .S0(n107_adj_1222), 
          .S1(n104_adj_1221));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_23 (.A0(n104_adj_1284), .B0(n2449), .C0(n101_adj_1252), 
          .D0(n1455), .A1(n101_adj_1283), .B1(n2449), .C1(n98_adj_1251), 
          .D1(n1454), .CIN(n12995), .COUT(n12996), .S0(n101_adj_1220), 
          .S1(n98_adj_1219));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_25 (.A0(n98_adj_1282), .B0(n2449), .C0(n95_adj_1250), 
          .D0(n1453), .A1(n95_adj_1281), .B1(n2449), .C1(n92_adj_1249), 
          .D1(n1452), .CIN(n12996), .COUT(n12997), .S0(n95_adj_1218), 
          .S1(n92_adj_1217));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_27 (.A0(n92_adj_1280), .B0(n2449), .C0(n89_adj_1248), 
          .D0(n1451), .A1(n89_adj_1279), .B1(n2449), .C1(n86_adj_1247), 
          .D1(n1450), .CIN(n12997), .COUT(n12998), .S0(n89_adj_1216), 
          .S1(n86_adj_1215));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_29 (.A0(n86_adj_1278), .B0(n2449), .C0(n83_adj_1246), 
          .D0(n1449), .A1(n83_adj_1277), .B1(n2449), .C1(n80_adj_1245), 
          .D1(n1448), .CIN(n12998), .COUT(n12999), .S0(n83_adj_1214), 
          .S1(n80_adj_1213));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_31 (.A0(n80_adj_1276), .B0(n2449), .C0(n77_adj_1244), 
          .D0(n1447), .A1(n77_adj_1275), .B1(n2449), .C1(n74_adj_1243), 
          .D1(n1446), .CIN(n12999), .COUT(n13000), .S0(n77_adj_1212), 
          .S1(n74_adj_1211));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_430_add_4_33 (.A0(n74_adj_1274), .B0(n2449), .C0(n71_adj_1242), 
          .D0(n1445), .A1(n71_adj_1273), .B1(n2449), .C1(n68_adj_1241), 
          .D1(n1444), .CIN(n13000), .S0(n71_adj_1210), .S1(n2516));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_430_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_430_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_430_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_430_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_1303), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13003), .S1(n158_adj_1271));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_427_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_1302), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_1301), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13003), .COUT(n13004), .S0(n155_adj_1270), 
          .S1(n152_adj_1269));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_1300), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_1299), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13004), .COUT(n13005), .S0(n149_adj_1268), 
          .S1(n146_adj_1267));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_1298), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_1297), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13005), .COUT(n13006), .S0(n143_adj_1266), 
          .S1(n140_adj_1265));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_1296), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_1295), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13006), .COUT(n13007), .S0(n137_adj_1264), 
          .S1(n134_adj_1263));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_1294), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_1293), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13007), .COUT(n13008), .S0(n131_adj_1262), 
          .S1(n128_adj_1261));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_1292), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_1291), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13008), .COUT(n13009), .S0(n125_adj_1260), 
          .S1(n122_adj_1259));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_1290), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_1289), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13009), .COUT(n13010), .S0(n119_adj_1258), 
          .S1(n116_adj_1257));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_1288), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_1287), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13010), .COUT(n13011), .S0(n113_adj_1256), 
          .S1(n110_adj_1255));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_1286), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_1285), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13011), .COUT(n13012), .S0(n107_adj_1254), 
          .S1(n104_adj_1253));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_1284), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_1283), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13012), .COUT(n13013), .S0(n101_adj_1252), 
          .S1(n98_adj_1251));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_1282), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_1281), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13013), .COUT(n13014), .S0(n95_adj_1250), 
          .S1(n92_adj_1249));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_1280), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_1279), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13014), .COUT(n13015), .S0(n89_adj_1248), 
          .S1(n86_adj_1247));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_1278), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_1277), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13015), .COUT(n13016), .S0(n83_adj_1246), 
          .S1(n80_adj_1245));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_1276), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_1275), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13016), .COUT(n13017), .S0(n77_adj_1244), 
          .S1(n74_adj_1243));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_427_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_427_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_1274), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_1273), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13017), .S0(n71_adj_1242), .S1(n68_adj_1241));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_427_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_427_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_427_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_427_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2382), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n13022));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_424_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_424_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_3 (.A0(det_q4_28[0]), .B0(n2382), .C0(n161_adj_1272), 
          .D0(n1475), .A1(n161_adj_1208), .B1(n2382), .C1(n158_adj_1334), 
          .D1(n1474), .CIN(n13022), .COUT(n13023), .S0(n161_adj_1303), 
          .S1(n158_adj_1302));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_5 (.A0(n158_adj_1207), .B0(n2382), .C0(n155_adj_1333), 
          .D0(n1473), .A1(n155_adj_1206), .B1(n2382), .C1(n152_adj_1332), 
          .D1(n1472), .CIN(n13023), .COUT(n13024), .S0(n155_adj_1301), 
          .S1(n152_adj_1300));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_7 (.A0(n152_adj_1205), .B0(n2382), .C0(n149_adj_1331), 
          .D0(n1471), .A1(n149_adj_1204), .B1(n2382), .C1(n146_adj_1330), 
          .D1(n1470), .CIN(n13024), .COUT(n13025), .S0(n149_adj_1299), 
          .S1(n146_adj_1298));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_9 (.A0(n146_adj_1203), .B0(n2382), .C0(n143_adj_1329), 
          .D0(n1469), .A1(n143_adj_1202), .B1(n2382), .C1(n140_adj_1328), 
          .D1(n1468), .CIN(n13025), .COUT(n13026), .S0(n143_adj_1297), 
          .S1(n140_adj_1296));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_11 (.A0(n140_adj_1201), .B0(n2382), .C0(n137_adj_1327), 
          .D0(n1467), .A1(n137_adj_1200), .B1(n2382), .C1(n134_adj_1326), 
          .D1(n1466), .CIN(n13026), .COUT(n13027), .S0(n137_adj_1295), 
          .S1(n134_adj_1294));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_13 (.A0(n134_adj_1199), .B0(n2382), .C0(n131_adj_1325), 
          .D0(n1465), .A1(n131_adj_1198), .B1(n2382), .C1(n128_adj_1324), 
          .D1(n1464), .CIN(n13027), .COUT(n13028), .S0(n131_adj_1293), 
          .S1(n128_adj_1292));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_15 (.A0(n128_adj_1197), .B0(n2382), .C0(n125_adj_1323), 
          .D0(n1463), .A1(n125_adj_1196), .B1(n2382), .C1(n122_adj_1322), 
          .D1(n1462), .CIN(n13028), .COUT(n13029), .S0(n125_adj_1291), 
          .S1(n122_adj_1290));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_17 (.A0(n122_adj_1195), .B0(n2382), .C0(n119_adj_1321), 
          .D0(n1461), .A1(n119_adj_1194), .B1(n2382), .C1(n116_adj_1320), 
          .D1(n1460), .CIN(n13029), .COUT(n13030), .S0(n119_adj_1289), 
          .S1(n116_adj_1288));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_19 (.A0(n116_adj_1193), .B0(n2382), .C0(n113_adj_1319), 
          .D0(n1459), .A1(n113_adj_1192), .B1(n2382), .C1(n110_adj_1318), 
          .D1(n1458), .CIN(n13030), .COUT(n13031), .S0(n113_adj_1287), 
          .S1(n110_adj_1286));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_21 (.A0(n110_adj_1191), .B0(n2382), .C0(n107_adj_1317), 
          .D0(n1457), .A1(n107_adj_1190), .B1(n2382), .C1(n104_adj_1316), 
          .D1(n1456), .CIN(n13031), .COUT(n13032), .S0(n107_adj_1285), 
          .S1(n104_adj_1284));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_23 (.A0(n104_adj_1189), .B0(n2382), .C0(n101_adj_1315), 
          .D0(n1455), .A1(n101_adj_1188), .B1(n2382), .C1(n98_adj_1314), 
          .D1(n1454), .CIN(n13032), .COUT(n13033), .S0(n101_adj_1283), 
          .S1(n98_adj_1282));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_25 (.A0(n98_adj_1187), .B0(n2382), .C0(n95_adj_1313), 
          .D0(n1453), .A1(n95_adj_1186), .B1(n2382), .C1(n92_adj_1312), 
          .D1(n1452), .CIN(n13033), .COUT(n13034), .S0(n95_adj_1281), 
          .S1(n92_adj_1280));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_27 (.A0(n92_adj_1185), .B0(n2382), .C0(n89_adj_1311), 
          .D0(n1451), .A1(n89_adj_1184), .B1(n2382), .C1(n86_adj_1310), 
          .D1(n1450), .CIN(n13034), .COUT(n13035), .S0(n89_adj_1279), 
          .S1(n86_adj_1278));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_29 (.A0(n86_adj_1183), .B0(n2382), .C0(n83_adj_1309), 
          .D0(n1449), .A1(n83_adj_1182), .B1(n2382), .C1(n80_adj_1308), 
          .D1(n1448), .CIN(n13035), .COUT(n13036), .S0(n83_adj_1277), 
          .S1(n80_adj_1276));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_31 (.A0(n80_adj_1181), .B0(n2382), .C0(n77_adj_1307), 
          .D0(n1447), .A1(n77_adj_1180), .B1(n2382), .C1(n74_adj_1306), 
          .D1(n1446), .CIN(n13036), .COUT(n13037), .S0(n77_adj_1275), 
          .S1(n74_adj_1274));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_424_add_4_33 (.A0(n74_adj_1179), .B0(n2382), .C0(n71_adj_1305), 
          .D0(n1445), .A1(n71_adj_1178), .B1(n2382), .C1(n68_adj_1304), 
          .D1(n1444), .CIN(n13037), .S0(n71_adj_1273), .S1(n2449));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_424_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_424_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_424_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_424_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_1208), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13040), .S1(n158_adj_1334));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_421_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_1207), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_1206), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13040), .COUT(n13041), .S0(n155_adj_1333), 
          .S1(n152_adj_1332));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_1205), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_1204), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13041), .COUT(n13042), .S0(n149_adj_1331), 
          .S1(n146_adj_1330));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_1203), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_1202), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13042), .COUT(n13043), .S0(n143_adj_1329), 
          .S1(n140_adj_1328));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_1201), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_1200), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13043), .COUT(n13044), .S0(n137_adj_1327), 
          .S1(n134_adj_1326));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_1199), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_1198), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13044), .COUT(n13045), .S0(n131_adj_1325), 
          .S1(n128_adj_1324));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_1197), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_1196), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13045), .COUT(n13046), .S0(n125_adj_1323), 
          .S1(n122_adj_1322));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_1195), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_1194), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13046), .COUT(n13047), .S0(n119_adj_1321), 
          .S1(n116_adj_1320));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_1193), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_1192), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13047), .COUT(n13048), .S0(n113_adj_1319), 
          .S1(n110_adj_1318));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_1191), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_1190), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13048), .COUT(n13049), .S0(n107_adj_1317), 
          .S1(n104_adj_1316));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_1189), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_1188), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13049), .COUT(n13050), .S0(n101_adj_1315), 
          .S1(n98_adj_1314));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_1187), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_1186), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13050), .COUT(n13051), .S0(n95_adj_1313), 
          .S1(n92_adj_1312));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_1185), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_1184), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13051), .COUT(n13052), .S0(n89_adj_1311), 
          .S1(n86_adj_1310));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_1183), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_1182), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13052), .COUT(n13053), .S0(n83_adj_1309), 
          .S1(n80_adj_1308));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_1181), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_1180), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13053), .COUT(n13054), .S0(n77_adj_1307), 
          .S1(n74_adj_1306));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_421_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_421_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_1179), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_1178), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13054), .S0(n71_adj_1305), .S1(n68_adj_1304));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_421_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_421_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_421_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_421_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_2 (.A0(n1475), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1474), .B1(n161_adj_2065), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13057), .S1(n158_adj_1365));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_418_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_4 (.A0(n1473), .B0(n158_adj_2064), .C0(GND_net), 
          .D0(VCC_net), .A1(n1472), .B1(n155_adj_2063), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13057), .COUT(n13058), .S0(n155_adj_1364), 
          .S1(n152_adj_1363));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_6 (.A0(n1471), .B0(n152_adj_2062), .C0(GND_net), 
          .D0(VCC_net), .A1(n1470), .B1(n149_adj_2061), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13058), .COUT(n13059), .S0(n149_adj_1362), 
          .S1(n146_adj_1361));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_8 (.A0(n1469), .B0(n146_adj_2060), .C0(GND_net), 
          .D0(VCC_net), .A1(n1468), .B1(n143_adj_2059), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13059), .COUT(n13060), .S0(n143_adj_1360), 
          .S1(n140_adj_1359));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_10 (.A0(n1467), .B0(n140_adj_2058), .C0(GND_net), 
          .D0(VCC_net), .A1(n1466), .B1(n137_adj_2057), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13060), .COUT(n13061), .S0(n137_adj_1358), 
          .S1(n134_adj_1357));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_12 (.A0(n1465), .B0(n134_adj_2056), .C0(GND_net), 
          .D0(VCC_net), .A1(n1464), .B1(n131_adj_2055), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13061), .COUT(n13062), .S0(n131_adj_1356), 
          .S1(n128_adj_1355));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_14 (.A0(n1463), .B0(n128_adj_2054), .C0(GND_net), 
          .D0(VCC_net), .A1(n1462), .B1(n125_adj_2053), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13062), .COUT(n13063), .S0(n125_adj_1354), 
          .S1(n122_adj_1353));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_16 (.A0(n1461), .B0(n122_adj_2052), .C0(GND_net), 
          .D0(VCC_net), .A1(n1460), .B1(n119_adj_2051), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13063), .COUT(n13064), .S0(n119_adj_1352), 
          .S1(n116_adj_1351));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_18 (.A0(n1459), .B0(n116_adj_2050), .C0(GND_net), 
          .D0(VCC_net), .A1(n1458), .B1(n113_adj_2049), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13064), .COUT(n13065), .S0(n113_adj_1350), 
          .S1(n110_adj_1349));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_20 (.A0(n1457), .B0(n110_adj_2048), .C0(GND_net), 
          .D0(VCC_net), .A1(n1456), .B1(n107_adj_2047), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13065), .COUT(n13066), .S0(n107_adj_1348), 
          .S1(n104_adj_1347));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_22 (.A0(n1455), .B0(n104_adj_2046), .C0(GND_net), 
          .D0(VCC_net), .A1(n1454), .B1(n101_adj_2045), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13066), .COUT(n13067), .S0(n101_adj_1346), 
          .S1(n98_adj_1345));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_24 (.A0(n1453), .B0(n98_adj_2044), .C0(GND_net), 
          .D0(VCC_net), .A1(n1452), .B1(n95_adj_2043), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13067), .COUT(n13068), .S0(n95_adj_1344), 
          .S1(n92_adj_1343));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_26 (.A0(n1451), .B0(n92_adj_2042), .C0(GND_net), 
          .D0(VCC_net), .A1(n1450), .B1(n89_adj_2041), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13068), .COUT(n13069), .S0(n89_adj_1342), 
          .S1(n86_adj_1341));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_28 (.A0(n1449), .B0(n86_adj_2040), .C0(GND_net), 
          .D0(VCC_net), .A1(n1448), .B1(n83_adj_2039), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13069), .COUT(n13070), .S0(n83_adj_1340), 
          .S1(n80_adj_1339));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_30 (.A0(n1447), .B0(n80_adj_2038), .C0(GND_net), 
          .D0(VCC_net), .A1(n1446), .B1(n77_adj_2037), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13070), .COUT(n13071), .S0(n77_adj_1338), 
          .S1(n74_adj_1337));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_418_add_4_32 (.A0(n1445), .B0(n74_adj_2036), .C0(GND_net), 
          .D0(VCC_net), .A1(n1444), .B1(n71_adj_2035), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13071), .S0(n71_adj_1336), .S1(n68_adj_1335));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_418_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_418_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_418_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_418_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_2065), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13074), .S1(n158_adj_1397));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_415_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_2064), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_2063), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13074), .COUT(n13075), .S0(n155_adj_1396), 
          .S1(n152_adj_1395));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_2062), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_2061), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13075), .COUT(n13076), .S0(n149_adj_1394), 
          .S1(n146_adj_1393));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_2060), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_2059), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13076), .COUT(n13077), .S0(n143_adj_1392), 
          .S1(n140_adj_1391));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_2058), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_2057), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13077), .COUT(n13078), .S0(n137_adj_1390), 
          .S1(n134_adj_1389));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_2056), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_2055), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13078), .COUT(n13079), .S0(n131_adj_1388), 
          .S1(n128_adj_1387));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_2054), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_2053), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13079), .COUT(n13080), .S0(n125_adj_1386), 
          .S1(n122_adj_1385));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_2052), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_2051), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13080), .COUT(n13081), .S0(n119_adj_1384), 
          .S1(n116_adj_1383));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_2050), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_2049), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13081), .COUT(n13082), .S0(n113_adj_1382), 
          .S1(n110_adj_1381));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_2048), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_2047), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13082), .COUT(n13083), .S0(n107_adj_1380), 
          .S1(n104_adj_1379));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_2046), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_2045), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13083), .COUT(n13084), .S0(n101_adj_1378), 
          .S1(n98_adj_1377));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_2044), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_2043), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13084), .COUT(n13085), .S0(n95_adj_1376), 
          .S1(n92_adj_1375));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_2042), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_2041), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13085), .COUT(n13086), .S0(n89_adj_1374), 
          .S1(n86_adj_1373));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_2040), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_2039), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13086), .COUT(n13087), .S0(n83_adj_1372), 
          .S1(n80_adj_1371));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_2038), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_2037), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13087), .COUT(n13088), .S0(n77_adj_1370), 
          .S1(n74_adj_1369));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_415_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_415_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_2036), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_2035), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13088), .S0(n71_adj_1368), .S1(n68_adj_1367));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_415_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_415_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_415_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_415_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13835), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13090), .S1(n161_adj_1429));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_412_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_3 (.A0(n161_adj_1366), .B0(n13835), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1365), .B1(n13835), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13090), .COUT(n13091), .S0(n158_adj_1428), 
          .S1(n155_adj_1427));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_5 (.A0(n155_adj_1364), .B0(n13835), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1363), .B1(n13835), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13091), .COUT(n13092), .S0(n152_adj_1426), 
          .S1(n149_adj_1425));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_7 (.A0(n149_adj_1362), .B0(n13835), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1361), .B1(n13835), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13092), .COUT(n13093), .S0(n146_adj_1424), 
          .S1(n143_adj_1423));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_9 (.A0(n143_adj_1360), .B0(n13835), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1359), .B1(n13835), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13093), .COUT(n13094), .S0(n140_adj_1422), 
          .S1(n137_adj_1421));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_11 (.A0(n137_adj_1358), .B0(n13835), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1357), .B1(n13835), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13094), .COUT(n13095), .S0(n134_adj_1420), 
          .S1(n131_adj_1419));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_13 (.A0(n131_adj_1356), .B0(n13835), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1355), .B1(n13835), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13095), .COUT(n13096), .S0(n128_adj_1418), 
          .S1(n125_adj_1417));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_15 (.A0(n125_adj_1354), .B0(n13835), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1353), .B1(n13835), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13096), .COUT(n13097), .S0(n122_adj_1416), 
          .S1(n119_adj_1415));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_17 (.A0(n119_adj_1352), .B0(n13835), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1351), .B1(n13835), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13097), .COUT(n13098), .S0(n116_adj_1414), 
          .S1(n113_adj_1413));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_19 (.A0(n113_adj_1350), .B0(n13835), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1349), .B1(n13835), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13098), .COUT(n13099), .S0(n110_adj_1412), 
          .S1(n107_adj_1411));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_21 (.A0(n107_adj_1348), .B0(n13835), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1347), .B1(n13835), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13099), .COUT(n13100), .S0(n104_adj_1410), 
          .S1(n101_adj_1409));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_23 (.A0(n101_adj_1346), .B0(n13835), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1345), .B1(n13835), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13100), .COUT(n13101), .S0(n98_adj_1408), 
          .S1(n95_adj_1407));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_25 (.A0(n95_adj_1344), .B0(n13835), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1343), .B1(n13835), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13101), .COUT(n13102), .S0(n92_adj_1406), 
          .S1(n89_adj_1405));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_27 (.A0(n89_adj_1342), .B0(n13835), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1341), .B1(n13835), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13102), .COUT(n13103), .S0(n86_adj_1404), 
          .S1(n83_adj_1403));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_29 (.A0(n83_adj_1340), .B0(n13835), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1339), .B1(n13835), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13103), .COUT(n13104), .S0(n80_adj_1402), 
          .S1(n77_adj_1401));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_31 (.A0(n77_adj_1338), .B0(n13835), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1337), .B1(n13835), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13104), .COUT(n13105), .S0(n74_adj_1400), 
          .S1(n71_adj_1399));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_412_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_412_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_412_add_4_33 (.A0(n1444), .B0(n13835), .C0(n71_adj_1336), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13105), .S0(n68_adj_1398));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_412_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_412_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_412_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_412_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13835), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13106), .S1(n161_adj_1461));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_409_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_3 (.A0(n161_adj_1272), .B0(n13835), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1397), .B1(n13835), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13106), .COUT(n13107), .S0(n158_adj_1460), 
          .S1(n155_adj_1459));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_5 (.A0(n155_adj_1396), .B0(n13835), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1395), .B1(n13835), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13107), .COUT(n13108), .S0(n152_adj_1458), 
          .S1(n149_adj_1457));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_7 (.A0(n149_adj_1394), .B0(n13835), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1393), .B1(n13835), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13108), .COUT(n13109), .S0(n146_adj_1456), 
          .S1(n143_adj_1455));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_9 (.A0(n143_adj_1392), .B0(n13835), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1391), .B1(n13835), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13109), .COUT(n13110), .S0(n140_adj_1454), 
          .S1(n137_adj_1453));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_11 (.A0(n137_adj_1390), .B0(n13835), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1389), .B1(n13835), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13110), .COUT(n13111), .S0(n134_adj_1452), 
          .S1(n131_adj_1451));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_13 (.A0(n131_adj_1388), .B0(n13835), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1387), .B1(n13835), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13111), .COUT(n13112), .S0(n128_adj_1450), 
          .S1(n125_adj_1449));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_15 (.A0(n125_adj_1386), .B0(n13835), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1385), .B1(n13835), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13112), .COUT(n13113), .S0(n122_adj_1448), 
          .S1(n119_adj_1447));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_17 (.A0(n119_adj_1384), .B0(n13835), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1383), .B1(n13835), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13113), .COUT(n13114), .S0(n116_adj_1446), 
          .S1(n113_adj_1445));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_19 (.A0(n113_adj_1382), .B0(n13835), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1381), .B1(n13835), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13114), .COUT(n13115), .S0(n110_adj_1444), 
          .S1(n107_adj_1443));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_21 (.A0(n107_adj_1380), .B0(n13835), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1379), .B1(n13835), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13115), .COUT(n13116), .S0(n104_adj_1442), 
          .S1(n101_adj_1441));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_23 (.A0(n101_adj_1378), .B0(n13835), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1377), .B1(n13835), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13116), .COUT(n13117), .S0(n98_adj_1440), 
          .S1(n95_adj_1439));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_25 (.A0(n95_adj_1376), .B0(n13835), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1375), .B1(n13835), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13117), .COUT(n13118), .S0(n92_adj_1438), 
          .S1(n89_adj_1437));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_27 (.A0(n89_adj_1374), .B0(n13835), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1373), .B1(n13835), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13118), .COUT(n13119), .S0(n86_adj_1436), 
          .S1(n83_adj_1435));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_29 (.A0(n83_adj_1372), .B0(n13835), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1371), .B1(n13835), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13119), .COUT(n13120), .S0(n80_adj_1434), 
          .S1(n77_adj_1433));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_31 (.A0(n77_adj_1370), .B0(n13835), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1369), .B1(n13835), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13120), .COUT(n13121), .S0(n74_adj_1432), 
          .S1(n71_adj_1431));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_409_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_409_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_409_add_4_33 (.A0(n1444), .B0(n13835), .C0(n71_adj_1368), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13121), .S0(n68_adj_1430));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_409_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_409_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_409_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_409_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13829), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13122), .S1(n161_adj_1493));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_361_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_3 (.A0(n161_adj_1619), .B0(n13829), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1618), .B1(n13829), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13122), .COUT(n13123), .S0(n158_adj_1492), 
          .S1(n155_adj_1491));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_5 (.A0(n155_adj_1617), .B0(n13829), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1616), .B1(n13829), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13123), .COUT(n13124), .S0(n152_adj_1490), 
          .S1(n149_adj_1489));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_7 (.A0(n149_adj_1615), .B0(n13829), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1614), .B1(n13829), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13124), .COUT(n13125), .S0(n146_adj_1488), 
          .S1(n143_adj_1487));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_9 (.A0(n143_adj_1613), .B0(n13829), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1612), .B1(n13829), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13125), .COUT(n13126), .S0(n140_adj_1486), 
          .S1(n137_adj_1485));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_11 (.A0(n137_adj_1611), .B0(n13829), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1610), .B1(n13829), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13126), .COUT(n13127), .S0(n134_adj_1484), 
          .S1(n131_adj_1483));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_13 (.A0(n131_adj_1609), .B0(n13829), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1608), .B1(n13829), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13127), .COUT(n13128), .S0(n128_adj_1482), 
          .S1(n125_adj_1481));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_15 (.A0(n125_adj_1607), .B0(n13829), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1606), .B1(n13829), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13128), .COUT(n13129), .S0(n122_adj_1480), 
          .S1(n119_adj_1479));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_17 (.A0(n119_adj_1605), .B0(n13829), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1604), .B1(n13829), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13129), .COUT(n13130), .S0(n116_adj_1478), 
          .S1(n113_adj_1477));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_19 (.A0(n113_adj_1603), .B0(n13829), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1602), .B1(n13829), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13130), .COUT(n13131), .S0(n110_adj_1476), 
          .S1(n107_adj_1475));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_21 (.A0(n107_adj_1601), .B0(n13829), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1600), .B1(n13829), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13131), .COUT(n13132), .S0(n104_adj_1474), 
          .S1(n101_adj_1473));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_23 (.A0(n101_adj_1599), .B0(n13829), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1598), .B1(n13829), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13132), .COUT(n13133), .S0(n98_adj_1472), 
          .S1(n95_adj_1471));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_25 (.A0(n95_adj_1597), .B0(n13829), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1596), .B1(n13829), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13133), .COUT(n13134), .S0(n92_adj_1470), 
          .S1(n89_adj_1469));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_27 (.A0(n89_adj_1595), .B0(n13829), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1594), .B1(n13829), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13134), .COUT(n13135), .S0(n86_adj_1468), 
          .S1(n83_adj_1467));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_29 (.A0(n83_adj_1593), .B0(n13829), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1592), .B1(n13829), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13135), .COUT(n13136), .S0(n80_adj_1466), 
          .S1(n77_adj_1465));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_31 (.A0(n77_adj_1591), .B0(n13829), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1590), .B1(n13829), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13136), .COUT(n13137), .S0(n74_adj_1464), 
          .S1(n71_adj_1463));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_361_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_361_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_361_add_4_33 (.A0(n1444), .B0(n13829), .C0(n71_adj_1589), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13137), .S0(n68_adj_1462));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_361_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_361_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_361_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_361_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13138), .S1(c_s[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_370_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_370_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_3 (.A0(c2_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13138), .COUT(n13139), .S0(c_s[1]), .S1(c_s[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_5 (.A0(c2_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13139), .COUT(n13140), .S0(c_s[3]), .S1(c_s[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_7 (.A0(c2_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13140), .COUT(n13141), .S0(c_s[5]), .S1(c_s[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_9 (.A0(c2_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13141), .COUT(n13142), .S0(c_s[7]), .S1(c_s[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_11 (.A0(c2_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13142), .COUT(n13143), .S0(c_s[9]), .S1(c_s[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_13 (.A0(c2_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13143), .COUT(n13144), .S0(c_s[11]), .S1(c_s[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_13.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_15 (.A0(c2_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13144), .COUT(n13145), .S0(c_s[13]), .S1(c_s[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_15.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_15.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_370_add_4_17 (.A0(c2_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c2_reg[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13145), .S0(c_s[15]), .S1(c_s[16]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(97[30:59])
    defparam _add_1_370_add_4_17.INIT0 = 16'h5555;
    defparam _add_1_370_add_4_17.INIT1 = 16'h5555;
    defparam _add_1_370_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_370_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_1240), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13148), .S1(n158_adj_1524));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_373_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_1239), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_1238), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13148), .COUT(n13149), .S0(n155_adj_1523), 
          .S1(n152_adj_1522));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_1237), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_1236), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13149), .COUT(n13150), .S0(n149_adj_1521), 
          .S1(n146_adj_1520));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_1235), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_1234), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13150), .COUT(n13151), .S0(n143_adj_1519), 
          .S1(n140_adj_1518));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_1233), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_1232), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13151), .COUT(n13152), .S0(n137_adj_1517), 
          .S1(n134_adj_1516));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_1231), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_1230), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13152), .COUT(n13153), .S0(n131_adj_1515), 
          .S1(n128_adj_1514));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_1229), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_1228), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13153), .COUT(n13154), .S0(n125_adj_1513), 
          .S1(n122_adj_1512));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_1227), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_1226), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13154), .COUT(n13155), .S0(n119_adj_1511), 
          .S1(n116_adj_1510));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_1225), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_1224), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13155), .COUT(n13156), .S0(n113_adj_1509), 
          .S1(n110_adj_1508));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_1223), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_1222), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13156), .COUT(n13157), .S0(n107_adj_1507), 
          .S1(n104_adj_1506));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_1221), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_1220), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13157), .COUT(n13158), .S0(n101_adj_1505), 
          .S1(n98_adj_1504));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_1219), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_1218), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13158), .COUT(n13159), .S0(n95_adj_1503), 
          .S1(n92_adj_1502));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_1217), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_1216), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13159), .COUT(n13160), .S0(n89_adj_1501), 
          .S1(n86_adj_1500));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_1215), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_1214), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13160), .COUT(n13161), .S0(n83_adj_1499), 
          .S1(n80_adj_1498));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_1213), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_1212), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13161), .COUT(n13162), .S0(n77_adj_1497), 
          .S1(n74_adj_1496));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_373_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_373_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_1211), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_1210), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13162), .S0(n71_adj_1495), .S1(n68_adj_1494));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_373_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_373_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_373_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_373_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2516), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n13167));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_376_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_376_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_3 (.A0(n1475), .B0(n2516), .C0(det_q4_28[0]), 
          .D0(VCC_net), .A1(n1474), .B1(n2516), .C1(n161_adj_1240), 
          .D1(VCC_net), .CIN(n13167), .COUT(n13168), .S0(n161_adj_1555), 
          .S1(n158_adj_1554));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_3.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_3.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_5 (.A0(n1473), .B0(n2516), .C0(n158_adj_1239), 
          .D0(VCC_net), .A1(n1472), .B1(n2516), .C1(n155_adj_1238), 
          .D1(VCC_net), .CIN(n13168), .COUT(n13169), .S0(n155_adj_1553), 
          .S1(n152_adj_1552));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_5.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_5.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_7 (.A0(n1471), .B0(n2516), .C0(n152_adj_1237), 
          .D0(VCC_net), .A1(n1470), .B1(n2516), .C1(n149_adj_1236), 
          .D1(VCC_net), .CIN(n13169), .COUT(n13170), .S0(n149_adj_1551), 
          .S1(n146_adj_1550));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_7.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_7.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_9 (.A0(n1469), .B0(n2516), .C0(n146_adj_1235), 
          .D0(VCC_net), .A1(n1468), .B1(n2516), .C1(n143_adj_1234), 
          .D1(VCC_net), .CIN(n13170), .COUT(n13171), .S0(n143_adj_1549), 
          .S1(n140_adj_1548));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_9.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_9.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_11 (.A0(n1467), .B0(n2516), .C0(n140_adj_1233), 
          .D0(VCC_net), .A1(n1466), .B1(n2516), .C1(n137_adj_1232), 
          .D1(VCC_net), .CIN(n13171), .COUT(n13172), .S0(n137_adj_1547), 
          .S1(n134_adj_1546));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_11.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_11.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_13 (.A0(n1465), .B0(n2516), .C0(n134_adj_1231), 
          .D0(VCC_net), .A1(n1464), .B1(n2516), .C1(n131_adj_1230), 
          .D1(VCC_net), .CIN(n13172), .COUT(n13173), .S0(n131_adj_1545), 
          .S1(n128_adj_1544));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_13.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_13.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_15 (.A0(n1463), .B0(n2516), .C0(n128_adj_1229), 
          .D0(VCC_net), .A1(n1462), .B1(n2516), .C1(n125_adj_1228), 
          .D1(VCC_net), .CIN(n13173), .COUT(n13174), .S0(n125_adj_1543), 
          .S1(n122_adj_1542));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_15.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_15.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_17 (.A0(n1461), .B0(n2516), .C0(n122_adj_1227), 
          .D0(VCC_net), .A1(n1460), .B1(n2516), .C1(n119_adj_1226), 
          .D1(VCC_net), .CIN(n13174), .COUT(n13175), .S0(n119_adj_1541), 
          .S1(n116_adj_1540));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_17.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_17.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_19 (.A0(n1459), .B0(n2516), .C0(n116_adj_1225), 
          .D0(VCC_net), .A1(n1458), .B1(n2516), .C1(n113_adj_1224), 
          .D1(VCC_net), .CIN(n13175), .COUT(n13176), .S0(n113_adj_1539), 
          .S1(n110_adj_1538));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_19.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_19.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_21 (.A0(n1457), .B0(n2516), .C0(n110_adj_1223), 
          .D0(VCC_net), .A1(n1456), .B1(n2516), .C1(n107_adj_1222), 
          .D1(VCC_net), .CIN(n13176), .COUT(n13177), .S0(n107_adj_1537), 
          .S1(n104_adj_1536));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_21.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_21.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_23 (.A0(n1455), .B0(n2516), .C0(n104_adj_1221), 
          .D0(VCC_net), .A1(n1454), .B1(n2516), .C1(n101_adj_1220), 
          .D1(VCC_net), .CIN(n13177), .COUT(n13178), .S0(n101_adj_1535), 
          .S1(n98_adj_1534));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_23.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_23.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_25 (.A0(n1453), .B0(n2516), .C0(n98_adj_1219), 
          .D0(VCC_net), .A1(n1452), .B1(n2516), .C1(n95_adj_1218), .D1(VCC_net), 
          .CIN(n13178), .COUT(n13179), .S0(n95_adj_1533), .S1(n92_adj_1532));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_25.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_25.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_27 (.A0(n1451), .B0(n2516), .C0(n92_adj_1217), 
          .D0(VCC_net), .A1(n1450), .B1(n2516), .C1(n89_adj_1216), .D1(VCC_net), 
          .CIN(n13179), .COUT(n13180), .S0(n89_adj_1531), .S1(n86_adj_1530));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_27.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_27.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_29 (.A0(n1449), .B0(n2516), .C0(n86_adj_1215), 
          .D0(VCC_net), .A1(n1448), .B1(n2516), .C1(n83_adj_1214), .D1(VCC_net), 
          .CIN(n13180), .COUT(n13181), .S0(n83_adj_1529), .S1(n80_adj_1528));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_29.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_29.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_31 (.A0(n1447), .B0(n2516), .C0(n80_adj_1213), 
          .D0(VCC_net), .A1(n1446), .B1(n2516), .C1(n77_adj_1212), .D1(VCC_net), 
          .CIN(n13181), .COUT(n13182), .S0(n77_adj_1527), .S1(n74_adj_1526));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_31.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_31.INIT1 = 16'h1212;
    defparam _add_1_376_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_376_add_4_33 (.A0(n1445), .B0(n2516), .C0(n74_adj_1211), 
          .D0(VCC_net), .A1(n71_adj_1210), .B1(n2516), .C1(n68_adj_1494), 
          .D1(n1444), .CIN(n13182), .S0(n71_adj_1525), .S1(n2583));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_376_add_4_33.INIT0 = 16'h1212;
    defparam _add_1_376_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_376_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_376_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13830), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13184), .S1(n161_adj_1587));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_379_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_3 (.A0(n161_adj_825), .B0(n13830), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_824), .B1(n13830), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13184), .COUT(n13185), .S0(n158_adj_1586), 
          .S1(n155_adj_1585));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_5 (.A0(n155_adj_823), .B0(n13830), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_822), .B1(n13830), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13185), .COUT(n13186), .S0(n152_adj_1584), 
          .S1(n149_adj_1583));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_7 (.A0(n149_adj_821), .B0(n13830), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_820), .B1(n13830), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13186), .COUT(n13187), .S0(n146_adj_1582), 
          .S1(n143_adj_1581));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_9 (.A0(n143_adj_819), .B0(n13830), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_818), .B1(n13830), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13187), .COUT(n13188), .S0(n140_adj_1580), 
          .S1(n137_adj_1579));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_11 (.A0(n137_adj_817), .B0(n13830), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_816), .B1(n13830), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13188), .COUT(n13189), .S0(n134_adj_1578), 
          .S1(n131_adj_1577));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_13 (.A0(n131_adj_815), .B0(n13830), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_814), .B1(n13830), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13189), .COUT(n13190), .S0(n128_adj_1576), 
          .S1(n125_adj_1575));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_15 (.A0(n125_adj_813), .B0(n13830), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_812), .B1(n13830), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13190), .COUT(n13191), .S0(n122_adj_1574), 
          .S1(n119_adj_1573));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_17 (.A0(n119_adj_811), .B0(n13830), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_810), .B1(n13830), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13191), .COUT(n13192), .S0(n116_adj_1572), 
          .S1(n113_adj_1571));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_19 (.A0(n113_adj_809), .B0(n13830), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_808), .B1(n13830), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13192), .COUT(n13193), .S0(n110_adj_1570), 
          .S1(n107_adj_1569));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_21 (.A0(n107_adj_807), .B0(n13830), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_806), .B1(n13830), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13193), .COUT(n13194), .S0(n104_adj_1568), 
          .S1(n101_adj_1567));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_23 (.A0(n101_adj_805), .B0(n13830), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_804), .B1(n13830), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13194), .COUT(n13195), .S0(n98_adj_1566), 
          .S1(n95_adj_1565));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_25 (.A0(n95_adj_803), .B0(n13830), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_802), .B1(n13830), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13195), .COUT(n13196), .S0(n92_adj_1564), 
          .S1(n89_adj_1563));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_27 (.A0(n89_adj_801), .B0(n13830), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_800), .B1(n13830), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13196), .COUT(n13197), .S0(n86_adj_1562), 
          .S1(n83_adj_1561));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_29 (.A0(n83_adj_799), .B0(n13830), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_798), .B1(n13830), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13197), .COUT(n13198), .S0(n80_adj_1560), 
          .S1(n77_adj_1559));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_31 (.A0(n77_adj_797), .B0(n13830), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_796), .B1(n13830), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13198), .COUT(n13199), .S0(n74_adj_1558), 
          .S1(n71_adj_1557));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_379_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_379_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_379_add_4_33 (.A0(n1444), .B0(n13830), .C0(n71_adj_795), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13199), .S0(n68_adj_1556));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_379_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_379_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_379_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_379_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13830), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13200), .S1(n161_adj_1619));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_382_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_3 (.A0(n161_adj_1811), .B0(n13830), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1810), .B1(n13830), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13200), .COUT(n13201), .S0(n158_adj_1618), 
          .S1(n155_adj_1617));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_5 (.A0(n155_adj_1809), .B0(n13830), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1808), .B1(n13830), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13201), .COUT(n13202), .S0(n152_adj_1616), 
          .S1(n149_adj_1615));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_7 (.A0(n149_adj_1807), .B0(n13830), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1806), .B1(n13830), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13202), .COUT(n13203), .S0(n146_adj_1614), 
          .S1(n143_adj_1613));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_9 (.A0(n143_adj_1805), .B0(n13830), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1804), .B1(n13830), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13203), .COUT(n13204), .S0(n140_adj_1612), 
          .S1(n137_adj_1611));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_11 (.A0(n137_adj_1803), .B0(n13830), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1802), .B1(n13830), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13204), .COUT(n13205), .S0(n134_adj_1610), 
          .S1(n131_adj_1609));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_13 (.A0(n131_adj_1801), .B0(n13830), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1800), .B1(n13830), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13205), .COUT(n13206), .S0(n128_adj_1608), 
          .S1(n125_adj_1607));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_15 (.A0(n125_adj_1799), .B0(n13830), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1798), .B1(n13830), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13206), .COUT(n13207), .S0(n122_adj_1606), 
          .S1(n119_adj_1605));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_17 (.A0(n119_adj_1797), .B0(n13830), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1796), .B1(n13830), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13207), .COUT(n13208), .S0(n116_adj_1604), 
          .S1(n113_adj_1603));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_19 (.A0(n113_adj_1795), .B0(n13830), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1794), .B1(n13830), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13208), .COUT(n13209), .S0(n110_adj_1602), 
          .S1(n107_adj_1601));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_21 (.A0(n107_adj_1793), .B0(n13830), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1792), .B1(n13830), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13209), .COUT(n13210), .S0(n104_adj_1600), 
          .S1(n101_adj_1599));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_23 (.A0(n101_adj_1791), .B0(n13830), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1790), .B1(n13830), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13210), .COUT(n13211), .S0(n98_adj_1598), 
          .S1(n95_adj_1597));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_25 (.A0(n95_adj_1789), .B0(n13830), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1788), .B1(n13830), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13211), .COUT(n13212), .S0(n92_adj_1596), 
          .S1(n89_adj_1595));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_27 (.A0(n89_adj_1787), .B0(n13830), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1786), .B1(n13830), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13212), .COUT(n13213), .S0(n86_adj_1594), 
          .S1(n83_adj_1593));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_29 (.A0(n83_adj_1785), .B0(n13830), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1784), .B1(n13830), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13213), .COUT(n13214), .S0(n80_adj_1592), 
          .S1(n77_adj_1591));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_31 (.A0(n77_adj_1783), .B0(n13830), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1782), .B1(n13830), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13214), .COUT(n13215), .S0(n74_adj_1590), 
          .S1(n71_adj_1589));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_382_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_382_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_382_add_4_33 (.A0(n1444), .B0(n13830), .C0(n71_adj_1781), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13215), .S0(n68_adj_1588));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_382_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_382_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_382_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_382_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13828), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13216), .S1(n161_adj_1651));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_493_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_3 (.A0(n161_adj_1366), .B0(n13828), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1970), .B1(n13828), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13216), .COUT(n13217), .S0(n158_adj_1650), 
          .S1(n155_adj_1649));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_5 (.A0(n155_adj_1969), .B0(n13828), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1968), .B1(n13828), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13217), .COUT(n13218), .S0(n152_adj_1648), 
          .S1(n149_adj_1647));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_7 (.A0(n149_adj_1967), .B0(n13828), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1966), .B1(n13828), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13218), .COUT(n13219), .S0(n146_adj_1646), 
          .S1(n143_adj_1645));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_9 (.A0(n143_adj_1965), .B0(n13828), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1964), .B1(n13828), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13219), .COUT(n13220), .S0(n140_adj_1644), 
          .S1(n137_adj_1643));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_11 (.A0(n137_adj_1963), .B0(n13828), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1962), .B1(n13828), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13220), .COUT(n13221), .S0(n134_adj_1642), 
          .S1(n131_adj_1641));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_13 (.A0(n131_adj_1961), .B0(n13828), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1960), .B1(n13828), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13221), .COUT(n13222), .S0(n128_adj_1640), 
          .S1(n125_adj_1639));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_15 (.A0(n125_adj_1959), .B0(n13828), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1958), .B1(n13828), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13222), .COUT(n13223), .S0(n122_adj_1638), 
          .S1(n119_adj_1637));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_17 (.A0(n119_adj_1957), .B0(n13828), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1956), .B1(n13828), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13223), .COUT(n13224), .S0(n116_adj_1636), 
          .S1(n113_adj_1635));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_19 (.A0(n113_adj_1955), .B0(n13828), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1954), .B1(n13828), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13224), .COUT(n13225), .S0(n110_adj_1634), 
          .S1(n107_adj_1633));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_21 (.A0(n107_adj_1953), .B0(n13828), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1952), .B1(n13828), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13225), .COUT(n13226), .S0(n104_adj_1632), 
          .S1(n101_adj_1631));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_23 (.A0(n101_adj_1951), .B0(n13828), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1950), .B1(n13828), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13226), .COUT(n13227), .S0(n98_adj_1630), 
          .S1(n95_adj_1629));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_25 (.A0(n95_adj_1949), .B0(n13828), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1948), .B1(n13828), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13227), .COUT(n13228), .S0(n92_adj_1628), 
          .S1(n89_adj_1627));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_27 (.A0(n89_adj_1947), .B0(n13828), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1946), .B1(n13828), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13228), .COUT(n13229), .S0(n86_adj_1626), 
          .S1(n83_adj_1625));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_29 (.A0(n83_adj_1945), .B0(n13828), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1944), .B1(n13828), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13229), .COUT(n13230), .S0(n80_adj_1624), 
          .S1(n77_adj_1623));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_31 (.A0(n77_adj_1943), .B0(n13828), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1942), .B1(n13828), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13230), .COUT(n13231), .S0(n74_adj_1622), 
          .S1(n71_adj_1621));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_493_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_493_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_493_add_4_33 (.A0(n1444), .B0(n13828), .C0(n71_adj_1941), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13231), .S0(n68_adj_1620));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_493_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_493_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_493_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_493_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_2 (.A0(n1475), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1474), .B1(n161_adj_346), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13232));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_355_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_4 (.A0(n1473), .B0(n158_adj_345), .C0(GND_net), 
          .D0(VCC_net), .A1(n1472), .B1(n155_adj_344), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13232), .COUT(n13233));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_6 (.A0(n1471), .B0(n152_adj_343), .C0(GND_net), 
          .D0(VCC_net), .A1(n1470), .B1(n149_adj_342), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13233), .COUT(n13234));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_8 (.A0(n1469), .B0(n146_adj_341), .C0(GND_net), 
          .D0(VCC_net), .A1(n1468), .B1(n143_adj_340), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13234), .COUT(n13235));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_10 (.A0(n1467), .B0(n140_adj_339), .C0(GND_net), 
          .D0(VCC_net), .A1(n1466), .B1(n137_adj_338), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13235), .COUT(n13236));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_12 (.A0(n1465), .B0(n134_adj_337), .C0(GND_net), 
          .D0(VCC_net), .A1(n1464), .B1(n131_adj_336), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13236), .COUT(n13237));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_14 (.A0(n1463), .B0(n128_adj_335), .C0(GND_net), 
          .D0(VCC_net), .A1(n1462), .B1(n125_adj_334), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13237), .COUT(n13238));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_16 (.A0(n1461), .B0(n122_adj_333), .C0(GND_net), 
          .D0(VCC_net), .A1(n1460), .B1(n119_adj_332), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13238), .COUT(n13239));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_18 (.A0(n1459), .B0(n116_adj_331), .C0(GND_net), 
          .D0(VCC_net), .A1(n1458), .B1(n113_adj_330), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13239), .COUT(n13240));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_20 (.A0(n1457), .B0(n110_adj_329), .C0(GND_net), 
          .D0(VCC_net), .A1(n1456), .B1(n107_adj_328), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13240), .COUT(n13241));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_22 (.A0(n1455), .B0(n104_adj_327), .C0(GND_net), 
          .D0(VCC_net), .A1(n1454), .B1(n101_adj_326), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13241), .COUT(n13242));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_24 (.A0(n1453), .B0(n98_adj_325), .C0(GND_net), 
          .D0(VCC_net), .A1(n1452), .B1(n95_adj_324), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13242), .COUT(n13243));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_26 (.A0(n1451), .B0(n92_adj_323), .C0(GND_net), 
          .D0(VCC_net), .A1(n1450), .B1(n89_adj_322), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13243), .COUT(n13244));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_28 (.A0(n1449), .B0(n86_adj_321), .C0(GND_net), 
          .D0(VCC_net), .A1(n1448), .B1(n83_adj_320), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13244), .COUT(n13245));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_30 (.A0(n1447), .B0(n80_adj_319), .C0(GND_net), 
          .D0(VCC_net), .A1(n1446), .B1(n77_adj_318), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13245), .COUT(n13246));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_355_add_4_32 (.A0(n1445), .B0(n74_adj_317), .C0(GND_net), 
          .D0(VCC_net), .A1(n1444), .B1(n71_adj_316), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13246), .S1(n68_adj_1652));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_355_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_355_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_355_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_355_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13833), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13248), .S1(n161_adj_1684));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_397_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_3 (.A0(n161_adj_2097), .B0(n13833), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_2096), .B1(n13833), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13248), .COUT(n13249), .S0(n158_adj_1683), 
          .S1(n155_adj_1682));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_5 (.A0(n155_adj_2095), .B0(n13833), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_2094), .B1(n13833), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13249), .COUT(n13250), .S0(n152_adj_1681), 
          .S1(n149_adj_1680));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_7 (.A0(n149_adj_2093), .B0(n13833), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_2092), .B1(n13833), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13250), .COUT(n13251), .S0(n146_adj_1679), 
          .S1(n143_adj_1678));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_9 (.A0(n143_adj_2091), .B0(n13833), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_2090), .B1(n13833), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13251), .COUT(n13252), .S0(n140_adj_1677), 
          .S1(n137_adj_1676));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_11 (.A0(n137_adj_2089), .B0(n13833), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_2088), .B1(n13833), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13252), .COUT(n13253), .S0(n134_adj_1675), 
          .S1(n131_adj_1674));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_13 (.A0(n131_adj_2087), .B0(n13833), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_2086), .B1(n13833), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13253), .COUT(n13254), .S0(n128_adj_1673), 
          .S1(n125_adj_1672));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_15 (.A0(n125_adj_2085), .B0(n13833), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_2084), .B1(n13833), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13254), .COUT(n13255), .S0(n122_adj_1671), 
          .S1(n119_adj_1670));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_17 (.A0(n119_adj_2083), .B0(n13833), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_2082), .B1(n13833), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13255), .COUT(n13256), .S0(n116_adj_1669), 
          .S1(n113_adj_1668));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_19 (.A0(n113_adj_2081), .B0(n13833), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_2080), .B1(n13833), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13256), .COUT(n13257), .S0(n110_adj_1667), 
          .S1(n107_adj_1666));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_21 (.A0(n107_adj_2079), .B0(n13833), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_2078), .B1(n13833), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13257), .COUT(n13258), .S0(n104_adj_1665), 
          .S1(n101_adj_1664));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_23 (.A0(n101_adj_2077), .B0(n13833), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_2076), .B1(n13833), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13258), .COUT(n13259), .S0(n98_adj_1663), 
          .S1(n95_adj_1662));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_25 (.A0(n95_adj_2075), .B0(n13833), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_2074), .B1(n13833), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13259), .COUT(n13260), .S0(n92_adj_1661), 
          .S1(n89_adj_1660));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_27 (.A0(n89_adj_2073), .B0(n13833), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_2072), .B1(n13833), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13260), .COUT(n13261), .S0(n86_adj_1659), 
          .S1(n83_adj_1658));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_29 (.A0(n83_adj_2071), .B0(n13833), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_2070), .B1(n13833), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13261), .COUT(n13262), .S0(n80_adj_1657), 
          .S1(n77_adj_1656));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_31 (.A0(n77_adj_2069), .B0(n13833), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_2068), .B1(n13833), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13262), .COUT(n13263), .S0(n74_adj_1655), 
          .S1(n71_adj_1654));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_397_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_397_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_397_add_4_33 (.A0(n1444), .B0(n13833), .C0(n71_adj_2067), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13263), .S0(n68_adj_1653));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_397_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_397_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_397_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_397_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13825), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13264), .S1(n161_adj_1716));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_514_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_3 (.A0(n161_adj_1875), .B0(n13825), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1874), .B1(n13825), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13264), .COUT(n13265), .S0(n158_adj_1715), 
          .S1(n155_adj_1714));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_5 (.A0(n155_adj_1873), .B0(n13825), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1872), .B1(n13825), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13265), .COUT(n13266), .S0(n152_adj_1713), 
          .S1(n149_adj_1712));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_7 (.A0(n149_adj_1871), .B0(n13825), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1870), .B1(n13825), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13266), .COUT(n13267), .S0(n146_adj_1711), 
          .S1(n143_adj_1710));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_9 (.A0(n143_adj_1869), .B0(n13825), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1868), .B1(n13825), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13267), .COUT(n13268), .S0(n140_adj_1709), 
          .S1(n137_adj_1708));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_11 (.A0(n137_adj_1867), .B0(n13825), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1866), .B1(n13825), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13268), .COUT(n13269), .S0(n134_adj_1707), 
          .S1(n131_adj_1706));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_13 (.A0(n131_adj_1865), .B0(n13825), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1864), .B1(n13825), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13269), .COUT(n13270), .S0(n128_adj_1705), 
          .S1(n125_adj_1704));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_15 (.A0(n125_adj_1863), .B0(n13825), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1862), .B1(n13825), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13270), .COUT(n13271), .S0(n122_adj_1703), 
          .S1(n119_adj_1702));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_17 (.A0(n119_adj_1861), .B0(n13825), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1860), .B1(n13825), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13271), .COUT(n13272), .S0(n116_adj_1701), 
          .S1(n113_adj_1700));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_19 (.A0(n113_adj_1859), .B0(n13825), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1858), .B1(n13825), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13272), .COUT(n13273), .S0(n110_adj_1699), 
          .S1(n107_adj_1698));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_21 (.A0(n107_adj_1857), .B0(n13825), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1856), .B1(n13825), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13273), .COUT(n13274), .S0(n104_adj_1697), 
          .S1(n101_adj_1696));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_23 (.A0(n101_adj_1855), .B0(n13825), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1854), .B1(n13825), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13274), .COUT(n13275), .S0(n98_adj_1695), 
          .S1(n95_adj_1694));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_25 (.A0(n95_adj_1853), .B0(n13825), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1852), .B1(n13825), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13275), .COUT(n13276), .S0(n92_adj_1693), 
          .S1(n89_adj_1692));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_27 (.A0(n89_adj_1851), .B0(n13825), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1850), .B1(n13825), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13276), .COUT(n13277), .S0(n86_adj_1691), 
          .S1(n83_adj_1690));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_29 (.A0(n83_adj_1849), .B0(n13825), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1848), .B1(n13825), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13277), .COUT(n13278), .S0(n80_adj_1689), 
          .S1(n77_adj_1688));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_31 (.A0(n77_adj_1847), .B0(n13825), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1846), .B1(n13825), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13278), .COUT(n13279), .S0(n74_adj_1687), 
          .S1(n71_adj_1686));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_514_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_514_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_514_add_4_33 (.A0(n1444), .B0(n13825), .C0(n71_adj_1845), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13279), .S0(n68_adj_1685));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_514_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_514_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_514_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_514_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13825), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13280), .S1(n161_adj_1748));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_511_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_3 (.A0(n161_adj_1939), .B0(n13825), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1938), .B1(n13825), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13280), .COUT(n13281), .S0(n158_adj_1747), 
          .S1(n155_adj_1746));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_5 (.A0(n155_adj_1937), .B0(n13825), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1936), .B1(n13825), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13281), .COUT(n13282), .S0(n152_adj_1745), 
          .S1(n149_adj_1744));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_7 (.A0(n149_adj_1935), .B0(n13825), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1934), .B1(n13825), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13282), .COUT(n13283), .S0(n146_adj_1743), 
          .S1(n143_adj_1742));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_9 (.A0(n143_adj_1933), .B0(n13825), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1932), .B1(n13825), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13283), .COUT(n13284), .S0(n140_adj_1741), 
          .S1(n137_adj_1740));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_11 (.A0(n137_adj_1931), .B0(n13825), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1930), .B1(n13825), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13284), .COUT(n13285), .S0(n134_adj_1739), 
          .S1(n131_adj_1738));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_13 (.A0(n131_adj_1929), .B0(n13825), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1928), .B1(n13825), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13285), .COUT(n13286), .S0(n128_adj_1737), 
          .S1(n125_adj_1736));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_15 (.A0(n125_adj_1927), .B0(n13825), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1926), .B1(n13825), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13286), .COUT(n13287), .S0(n122_adj_1735), 
          .S1(n119_adj_1734));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_17 (.A0(n119_adj_1925), .B0(n13825), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1924), .B1(n13825), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13287), .COUT(n13288), .S0(n116_adj_1733), 
          .S1(n113_adj_1732));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_19 (.A0(n113_adj_1923), .B0(n13825), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1922), .B1(n13825), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13288), .COUT(n13289), .S0(n110_adj_1731), 
          .S1(n107_adj_1730));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_21 (.A0(n107_adj_1921), .B0(n13825), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1920), .B1(n13825), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13289), .COUT(n13290), .S0(n104_adj_1729), 
          .S1(n101_adj_1728));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_23 (.A0(n101_adj_1919), .B0(n13825), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1918), .B1(n13825), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13290), .COUT(n13291), .S0(n98_adj_1727), 
          .S1(n95_adj_1726));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_25 (.A0(n95_adj_1917), .B0(n13825), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1916), .B1(n13825), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13291), .COUT(n13292), .S0(n92_adj_1725), 
          .S1(n89_adj_1724));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_27 (.A0(n89_adj_1915), .B0(n13825), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1914), .B1(n13825), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13292), .COUT(n13293), .S0(n86_adj_1723), 
          .S1(n83_adj_1722));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_29 (.A0(n83_adj_1913), .B0(n13825), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1912), .B1(n13825), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13293), .COUT(n13294), .S0(n80_adj_1721), 
          .S1(n77_adj_1720));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_31 (.A0(n77_adj_1911), .B0(n13825), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1910), .B1(n13825), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13294), .COUT(n13295), .S0(n74_adj_1719), 
          .S1(n71_adj_1718));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_511_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_511_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_511_add_4_33 (.A0(n1444), .B0(n13825), .C0(n71_adj_1909), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13295), .S0(n68_adj_1717));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_511_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_511_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_511_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_511_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13297), .S1(n158_adj_1779));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_490_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_4 (.A0(det_q4_28[3]), .B0(n158), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13297), .COUT(n13298), .S0(n155_adj_1778), 
          .S1(n152_adj_1777));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_6 (.A0(det_q4_28[5]), .B0(n152), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13298), .COUT(n13299), .S0(n149_adj_1776), 
          .S1(n146_adj_1775));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_8 (.A0(det_q4_28[7]), .B0(n146), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13299), .COUT(n13300), .S0(n143_adj_1774), 
          .S1(n140_adj_1773));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_10 (.A0(det_q4_28[9]), .B0(n140), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13300), .COUT(n13301), .S0(n137_adj_1772), 
          .S1(n134_adj_1771));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_12 (.A0(det_q4_28[11]), .B0(n134), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13301), .COUT(n13302), .S0(n131_adj_1770), 
          .S1(n128_adj_1769));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_250), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13302), .COUT(n13303), .S0(n125_adj_1768), 
          .S1(n122_adj_1767));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_249), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13303), .COUT(n13304), .S0(n119_adj_1766), 
          .S1(n116_adj_1765));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_248), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13304), .COUT(n13305), .S0(n113_adj_1764), 
          .S1(n110_adj_1763));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_247), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13305), .COUT(n13306), .S0(n107_adj_1762), 
          .S1(n104_adj_1761));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_246), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13306), .COUT(n13307), .S0(n101_adj_1760), 
          .S1(n98_adj_1759));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_24 (.A0(det_q4_28[23]), .B0(n98), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13307), .COUT(n13308), .S0(n95_adj_1758), 
          .S1(n92_adj_1757));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_26 (.A0(det_q4_28[25]), .B0(n92), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13308), .COUT(n13309), .S0(n89_adj_1756), 
          .S1(n86_adj_1755));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_28 (.A0(det_q4_28[27]), .B0(n86), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13309), .COUT(n13310), .S0(n83_adj_1754), 
          .S1(n80_adj_1753));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_30 (.A0(det_q4_28[29]), .B0(n80), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13310), .COUT(n13311), .S0(n77_adj_1752), 
          .S1(n74_adj_1751));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_490_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_490_add_4_32 (.A0(det_q4_28[31]), .B0(n74), .C0(GND_net), 
          .D0(VCC_net), .A1(n71), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13311), .S0(n71_adj_1750), .S1(n68_adj_1749));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_490_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_490_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_490_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_490_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13831), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13313), .S1(n161_adj_1811));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_388_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_3 (.A0(n161_adj_282), .B0(n13831), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_281), .B1(n13831), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13313), .COUT(n13314), .S0(n158_adj_1810), 
          .S1(n155_adj_1809));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_5 (.A0(n155_adj_280), .B0(n13831), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_279), .B1(n13831), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13314), .COUT(n13315), .S0(n152_adj_1808), 
          .S1(n149_adj_1807));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_7 (.A0(n149_adj_278), .B0(n13831), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_277), .B1(n13831), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13315), .COUT(n13316), .S0(n146_adj_1806), 
          .S1(n143_adj_1805));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_9 (.A0(n143_adj_276), .B0(n13831), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_275), .B1(n13831), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13316), .COUT(n13317), .S0(n140_adj_1804), 
          .S1(n137_adj_1803));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_11 (.A0(n137_adj_274), .B0(n13831), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_273), .B1(n13831), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13317), .COUT(n13318), .S0(n134_adj_1802), 
          .S1(n131_adj_1801));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_13 (.A0(n131_adj_272), .B0(n13831), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_271), .B1(n13831), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13318), .COUT(n13319), .S0(n128_adj_1800), 
          .S1(n125_adj_1799));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_15 (.A0(n125_adj_270), .B0(n13831), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_269), .B1(n13831), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13319), .COUT(n13320), .S0(n122_adj_1798), 
          .S1(n119_adj_1797));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_17 (.A0(n119_adj_268), .B0(n13831), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_267), .B1(n13831), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13320), .COUT(n13321), .S0(n116_adj_1796), 
          .S1(n113_adj_1795));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_19 (.A0(n113_adj_266), .B0(n13831), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_265), .B1(n13831), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13321), .COUT(n13322), .S0(n110_adj_1794), 
          .S1(n107_adj_1793));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_21 (.A0(n107_adj_264), .B0(n13831), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_263), .B1(n13831), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13322), .COUT(n13323), .S0(n104_adj_1792), 
          .S1(n101_adj_1791));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_23 (.A0(n101_adj_262), .B0(n13831), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_261), .B1(n13831), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13323), .COUT(n13324), .S0(n98_adj_1790), 
          .S1(n95_adj_1789));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_25 (.A0(n95_adj_260), .B0(n13831), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_259), .B1(n13831), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13324), .COUT(n13325), .S0(n92_adj_1788), 
          .S1(n89_adj_1787));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_27 (.A0(n89_adj_258), .B0(n13831), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_257), .B1(n13831), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13325), .COUT(n13326), .S0(n86_adj_1786), 
          .S1(n83_adj_1785));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_29 (.A0(n83_adj_256), .B0(n13831), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_255), .B1(n13831), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13326), .COUT(n13327), .S0(n80_adj_1784), 
          .S1(n77_adj_1783));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_31 (.A0(n77_adj_254), .B0(n13831), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_253), .B1(n13831), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13327), .COUT(n13328), .S0(n74_adj_1782), 
          .S1(n71_adj_1781));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_388_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_388_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_388_add_4_33 (.A0(n1444), .B0(n13831), .C0(n71_adj_252), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13328), .S0(n68_adj_1780));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_388_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_388_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_388_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_388_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13833), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13329), .S1(n161_adj_1843));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_400_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_3 (.A0(n161_adj_2193), .B0(n13833), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_2192), .B1(n13833), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13329), .COUT(n13330), .S0(n158_adj_1842), 
          .S1(n155_adj_1841));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_5 (.A0(n155_adj_2191), .B0(n13833), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_2190), .B1(n13833), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13330), .COUT(n13331), .S0(n152_adj_1840), 
          .S1(n149_adj_1839));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_7 (.A0(n149_adj_2189), .B0(n13833), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_2188), .B1(n13833), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13331), .COUT(n13332), .S0(n146_adj_1838), 
          .S1(n143_adj_1837));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_9 (.A0(n143_adj_2187), .B0(n13833), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_2186), .B1(n13833), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13332), .COUT(n13333), .S0(n140_adj_1836), 
          .S1(n137_adj_1835));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_11 (.A0(n137_adj_2185), .B0(n13833), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_2184), .B1(n13833), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13333), .COUT(n13334), .S0(n134_adj_1834), 
          .S1(n131_adj_1833));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_13 (.A0(n131_adj_2183), .B0(n13833), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_2182), .B1(n13833), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13334), .COUT(n13335), .S0(n128_adj_1832), 
          .S1(n125_adj_1831));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_15 (.A0(n125_adj_2181), .B0(n13833), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_2180), .B1(n13833), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13335), .COUT(n13336), .S0(n122_adj_1830), 
          .S1(n119_adj_1829));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_17 (.A0(n119_adj_2179), .B0(n13833), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_2178), .B1(n13833), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13336), .COUT(n13337), .S0(n116_adj_1828), 
          .S1(n113_adj_1827));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_19 (.A0(n113_adj_2177), .B0(n13833), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_2176), .B1(n13833), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13337), .COUT(n13338), .S0(n110_adj_1826), 
          .S1(n107_adj_1825));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_21 (.A0(n107_adj_2175), .B0(n13833), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_2174), .B1(n13833), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13338), .COUT(n13339), .S0(n104_adj_1824), 
          .S1(n101_adj_1823));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_23 (.A0(n101_adj_2173), .B0(n13833), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_2172), .B1(n13833), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13339), .COUT(n13340), .S0(n98_adj_1822), 
          .S1(n95_adj_1821));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_25 (.A0(n95_adj_2171), .B0(n13833), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_2170), .B1(n13833), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13340), .COUT(n13341), .S0(n92_adj_1820), 
          .S1(n89_adj_1819));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_27 (.A0(n89_adj_2169), .B0(n13833), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_2168), .B1(n13833), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13341), .COUT(n13342), .S0(n86_adj_1818), 
          .S1(n83_adj_1817));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_29 (.A0(n83_adj_2167), .B0(n13833), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_2166), .B1(n13833), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13342), .COUT(n13343), .S0(n80_adj_1816), 
          .S1(n77_adj_1815));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_31 (.A0(n77_adj_2165), .B0(n13833), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_2164), .B1(n13833), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13343), .COUT(n13344), .S0(n74_adj_1814), 
          .S1(n71_adj_1813));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_400_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_400_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_400_add_4_33 (.A0(n1444), .B0(n13833), .C0(n71_adj_2163), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13344), .S0(n68_adj_1812));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_400_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_400_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_400_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_400_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13826), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13345), .S1(n161_adj_1875));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_508_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_3 (.A0(n161_adj_2002), .B0(n13826), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_2001), .B1(n13826), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13345), .COUT(n13346), .S0(n158_adj_1874), 
          .S1(n155_adj_1873));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_5 (.A0(n155_adj_2000), .B0(n13826), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1999), .B1(n13826), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13346), .COUT(n13347), .S0(n152_adj_1872), 
          .S1(n149_adj_1871));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_7 (.A0(n149_adj_1998), .B0(n13826), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1997), .B1(n13826), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13347), .COUT(n13348), .S0(n146_adj_1870), 
          .S1(n143_adj_1869));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_9 (.A0(n143_adj_1996), .B0(n13826), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1995), .B1(n13826), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13348), .COUT(n13349), .S0(n140_adj_1868), 
          .S1(n137_adj_1867));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_11 (.A0(n137_adj_1994), .B0(n13826), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1993), .B1(n13826), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13349), .COUT(n13350), .S0(n134_adj_1866), 
          .S1(n131_adj_1865));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_13 (.A0(n131_adj_1992), .B0(n13826), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1991), .B1(n13826), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13350), .COUT(n13351), .S0(n128_adj_1864), 
          .S1(n125_adj_1863));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_15 (.A0(n125_adj_1990), .B0(n13826), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1989), .B1(n13826), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13351), .COUT(n13352), .S0(n122_adj_1862), 
          .S1(n119_adj_1861));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_17 (.A0(n119_adj_1988), .B0(n13826), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1987), .B1(n13826), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13352), .COUT(n13353), .S0(n116_adj_1860), 
          .S1(n113_adj_1859));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_19 (.A0(n113_adj_1986), .B0(n13826), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1985), .B1(n13826), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13353), .COUT(n13354), .S0(n110_adj_1858), 
          .S1(n107_adj_1857));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_21 (.A0(n107_adj_1984), .B0(n13826), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1983), .B1(n13826), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13354), .COUT(n13355), .S0(n104_adj_1856), 
          .S1(n101_adj_1855));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_23 (.A0(n101_adj_1982), .B0(n13826), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1981), .B1(n13826), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13355), .COUT(n13356), .S0(n98_adj_1854), 
          .S1(n95_adj_1853));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_25 (.A0(n95_adj_1980), .B0(n13826), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1979), .B1(n13826), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13356), .COUT(n13357), .S0(n92_adj_1852), 
          .S1(n89_adj_1851));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_27 (.A0(n89_adj_1978), .B0(n13826), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1977), .B1(n13826), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13357), .COUT(n13358), .S0(n86_adj_1850), 
          .S1(n83_adj_1849));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_29 (.A0(n83_adj_1976), .B0(n13826), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1975), .B1(n13826), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13358), .COUT(n13359), .S0(n80_adj_1848), 
          .S1(n77_adj_1847));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_31 (.A0(n77_adj_1974), .B0(n13826), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1973), .B1(n13826), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13359), .COUT(n13360), .S0(n74_adj_1846), 
          .S1(n71_adj_1845));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_508_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_508_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_508_add_4_33 (.A0(n1444), .B0(n13826), .C0(n71_adj_1972), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13360), .S0(n68_adj_1844));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_508_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_508_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_508_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_508_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13832), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13361), .S1(n161_adj_1907));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_391_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_3 (.A0(n161_adj_1684), .B0(n13832), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1683), .B1(n13832), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13361), .COUT(n13362), .S0(n158_adj_1906), 
          .S1(n155_adj_1905));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_5 (.A0(n155_adj_1682), .B0(n13832), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1681), .B1(n13832), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13362), .COUT(n13363), .S0(n152_adj_1904), 
          .S1(n149_adj_1903));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_7 (.A0(n149_adj_1680), .B0(n13832), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1679), .B1(n13832), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13363), .COUT(n13364), .S0(n146_adj_1902), 
          .S1(n143_adj_1901));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_9 (.A0(n143_adj_1678), .B0(n13832), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1677), .B1(n13832), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13364), .COUT(n13365), .S0(n140_adj_1900), 
          .S1(n137_adj_1899));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_11 (.A0(n137_adj_1676), .B0(n13832), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1675), .B1(n13832), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13365), .COUT(n13366), .S0(n134_adj_1898), 
          .S1(n131_adj_1897));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_13 (.A0(n131_adj_1674), .B0(n13832), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1673), .B1(n13832), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13366), .COUT(n13367), .S0(n128_adj_1896), 
          .S1(n125_adj_1895));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_15 (.A0(n125_adj_1672), .B0(n13832), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1671), .B1(n13832), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13367), .COUT(n13368), .S0(n122_adj_1894), 
          .S1(n119_adj_1893));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_17 (.A0(n119_adj_1670), .B0(n13832), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1669), .B1(n13832), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13368), .COUT(n13369), .S0(n116_adj_1892), 
          .S1(n113_adj_1891));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_19 (.A0(n113_adj_1668), .B0(n13832), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1667), .B1(n13832), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13369), .COUT(n13370), .S0(n110_adj_1890), 
          .S1(n107_adj_1889));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_21 (.A0(n107_adj_1666), .B0(n13832), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1665), .B1(n13832), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13370), .COUT(n13371), .S0(n104_adj_1888), 
          .S1(n101_adj_1887));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_23 (.A0(n101_adj_1664), .B0(n13832), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1663), .B1(n13832), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13371), .COUT(n13372), .S0(n98_adj_1886), 
          .S1(n95_adj_1885));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_25 (.A0(n95_adj_1662), .B0(n13832), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1661), .B1(n13832), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13372), .COUT(n13373), .S0(n92_adj_1884), 
          .S1(n89_adj_1883));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_27 (.A0(n89_adj_1660), .B0(n13832), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1659), .B1(n13832), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13373), .COUT(n13374), .S0(n86_adj_1882), 
          .S1(n83_adj_1881));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_29 (.A0(n83_adj_1658), .B0(n13832), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1657), .B1(n13832), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13374), .COUT(n13375), .S0(n80_adj_1880), 
          .S1(n77_adj_1879));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_31 (.A0(n77_adj_1656), .B0(n13832), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1655), .B1(n13832), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13375), .COUT(n13376), .S0(n74_adj_1878), 
          .S1(n71_adj_1877));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_391_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_391_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_391_add_4_33 (.A0(n1444), .B0(n13832), .C0(n71_adj_1654), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13376), .S0(n68_adj_1876));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_391_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_391_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_391_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_391_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13826), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13377), .S1(n161_adj_1939));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_505_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_3 (.A0(n161_adj_2034), .B0(n13826), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_2033), .B1(n13826), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13377), .COUT(n13378), .S0(n158_adj_1938), 
          .S1(n155_adj_1937));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_5 (.A0(n155_adj_2032), .B0(n13826), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_2031), .B1(n13826), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13378), .COUT(n13379), .S0(n152_adj_1936), 
          .S1(n149_adj_1935));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_7 (.A0(n149_adj_2030), .B0(n13826), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_2029), .B1(n13826), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13379), .COUT(n13380), .S0(n146_adj_1934), 
          .S1(n143_adj_1933));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_9 (.A0(n143_adj_2028), .B0(n13826), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_2027), .B1(n13826), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13380), .COUT(n13381), .S0(n140_adj_1932), 
          .S1(n137_adj_1931));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_11 (.A0(n137_adj_2026), .B0(n13826), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_2025), .B1(n13826), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13381), .COUT(n13382), .S0(n134_adj_1930), 
          .S1(n131_adj_1929));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_13 (.A0(n131_adj_2024), .B0(n13826), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_2023), .B1(n13826), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13382), .COUT(n13383), .S0(n128_adj_1928), 
          .S1(n125_adj_1927));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_15 (.A0(n125_adj_2022), .B0(n13826), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_2021), .B1(n13826), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13383), .COUT(n13384), .S0(n122_adj_1926), 
          .S1(n119_adj_1925));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_17 (.A0(n119_adj_2020), .B0(n13826), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_2019), .B1(n13826), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13384), .COUT(n13385), .S0(n116_adj_1924), 
          .S1(n113_adj_1923));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_19 (.A0(n113_adj_2018), .B0(n13826), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_2017), .B1(n13826), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13385), .COUT(n13386), .S0(n110_adj_1922), 
          .S1(n107_adj_1921));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_21 (.A0(n107_adj_2016), .B0(n13826), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_2015), .B1(n13826), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13386), .COUT(n13387), .S0(n104_adj_1920), 
          .S1(n101_adj_1919));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_23 (.A0(n101_adj_2014), .B0(n13826), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_2013), .B1(n13826), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13387), .COUT(n13388), .S0(n98_adj_1918), 
          .S1(n95_adj_1917));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_25 (.A0(n95_adj_2012), .B0(n13826), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_2011), .B1(n13826), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13388), .COUT(n13389), .S0(n92_adj_1916), 
          .S1(n89_adj_1915));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_27 (.A0(n89_adj_2010), .B0(n13826), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_2009), .B1(n13826), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13389), .COUT(n13390), .S0(n86_adj_1914), 
          .S1(n83_adj_1913));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_29 (.A0(n83_adj_2008), .B0(n13826), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_2007), .B1(n13826), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13390), .COUT(n13391), .S0(n80_adj_1912), 
          .S1(n77_adj_1911));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_31 (.A0(n77_adj_2006), .B0(n13826), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_2005), .B1(n13826), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13391), .COUT(n13392), .S0(n74_adj_1910), 
          .S1(n71_adj_1909));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_505_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_505_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_505_add_4_33 (.A0(n1444), .B0(n13826), .C0(n71_adj_2004), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13392), .S0(n68_adj_1908));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_505_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_505_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_505_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_505_add_4_33.INJECT1_1 = "NO";
    LUT4 i1579_2_lut_4_lut (.A(n68_adj_1146), .B(n68_adj_1114), .C(n1410), 
         .D(inv_det_31__N_227), .Z(n33)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1579_2_lut_4_lut.init = 16'h0035;
    CCU2C _add_1_487_add_4_2 (.A0(n1475), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1474), .B1(n161), .C1(GND_net), .D1(VCC_net), 
          .COUT(n13394), .S1(n158_adj_1970));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_487_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_4 (.A0(n1473), .B0(n158), .C0(GND_net), .D0(VCC_net), 
          .A1(n1472), .B1(n155), .C1(GND_net), .D1(VCC_net), .CIN(n13394), 
          .COUT(n13395), .S0(n155_adj_1969), .S1(n152_adj_1968));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_6 (.A0(n1471), .B0(n152), .C0(GND_net), .D0(VCC_net), 
          .A1(n1470), .B1(n149), .C1(GND_net), .D1(VCC_net), .CIN(n13395), 
          .COUT(n13396), .S0(n149_adj_1967), .S1(n146_adj_1966));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_8 (.A0(n1469), .B0(n146), .C0(GND_net), .D0(VCC_net), 
          .A1(n1468), .B1(n143), .C1(GND_net), .D1(VCC_net), .CIN(n13396), 
          .COUT(n13397), .S0(n143_adj_1965), .S1(n140_adj_1964));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_10 (.A0(n1467), .B0(n140), .C0(GND_net), .D0(VCC_net), 
          .A1(n1466), .B1(n137), .C1(GND_net), .D1(VCC_net), .CIN(n13397), 
          .COUT(n13398), .S0(n137_adj_1963), .S1(n134_adj_1962));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_12 (.A0(n1465), .B0(n134), .C0(GND_net), .D0(VCC_net), 
          .A1(n1464), .B1(n131), .C1(GND_net), .D1(VCC_net), .CIN(n13398), 
          .COUT(n13399), .S0(n131_adj_1961), .S1(n128_adj_1960));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_14 (.A0(n1463), .B0(n128_adj_250), .C0(GND_net), 
          .D0(VCC_net), .A1(n1462), .B1(n125), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13399), .COUT(n13400), .S0(n125_adj_1959), .S1(n122_adj_1958));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_16 (.A0(n1461), .B0(n122_adj_249), .C0(GND_net), 
          .D0(VCC_net), .A1(n1460), .B1(n119), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13400), .COUT(n13401), .S0(n119_adj_1957), .S1(n116_adj_1956));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_18 (.A0(n1459), .B0(n116_adj_248), .C0(GND_net), 
          .D0(VCC_net), .A1(n1458), .B1(n113), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13401), .COUT(n13402), .S0(n113_adj_1955), .S1(n110_adj_1954));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_20 (.A0(n1457), .B0(n110_adj_247), .C0(GND_net), 
          .D0(VCC_net), .A1(n1456), .B1(n107), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13402), .COUT(n13403), .S0(n107_adj_1953), .S1(n104_adj_1952));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_22 (.A0(n1455), .B0(n104_adj_246), .C0(GND_net), 
          .D0(VCC_net), .A1(n1454), .B1(n101), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13403), .COUT(n13404), .S0(n101_adj_1951), .S1(n98_adj_1950));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_24 (.A0(n1453), .B0(n98), .C0(GND_net), .D0(VCC_net), 
          .A1(n1452), .B1(n95), .C1(GND_net), .D1(VCC_net), .CIN(n13404), 
          .COUT(n13405), .S0(n95_adj_1949), .S1(n92_adj_1948));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_26 (.A0(n1451), .B0(n92), .C0(GND_net), .D0(VCC_net), 
          .A1(n1450), .B1(n89), .C1(GND_net), .D1(VCC_net), .CIN(n13405), 
          .COUT(n13406), .S0(n89_adj_1947), .S1(n86_adj_1946));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_28 (.A0(n1449), .B0(n86), .C0(GND_net), .D0(VCC_net), 
          .A1(n1448), .B1(n83), .C1(GND_net), .D1(VCC_net), .CIN(n13406), 
          .COUT(n13407), .S0(n83_adj_1945), .S1(n80_adj_1944));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_30 (.A0(n1447), .B0(n80), .C0(GND_net), .D0(VCC_net), 
          .A1(n1446), .B1(n77), .C1(GND_net), .D1(VCC_net), .CIN(n13407), 
          .COUT(n13408), .S0(n77_adj_1943), .S1(n74_adj_1942));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_487_add_4_32 (.A0(n1445), .B0(n74), .C0(GND_net), .D0(VCC_net), 
          .A1(n1444), .B1(n71), .C1(GND_net), .D1(VCC_net), .CIN(n13408), 
          .S0(n71_adj_1941), .S1(n68_adj_1940));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_487_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_487_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_487_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_487_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n13410), .S1(b_s[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_358_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_358_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_3 (.A0(b2_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13410), .COUT(n13411), .S0(b_s[1]), .S1(b_s[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_5 (.A0(b2_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13411), .COUT(n13412), .S0(b_s[3]), .S1(b_s[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_7 (.A0(b2_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13412), .COUT(n13413), .S0(b_s[5]), .S1(b_s[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_9 (.A0(b2_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13413), .COUT(n13414), .S0(b_s[7]), .S1(b_s[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_11 (.A0(b2_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13414), .COUT(n13415), .S0(b_s[9]), .S1(b_s[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_13 (.A0(b2_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13415), .COUT(n13416), .S0(b_s[11]), .S1(b_s[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_13.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_15 (.A0(b2_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13416), .COUT(n13417), .S0(b_s[13]), .S1(b_s[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_15.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_15.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_358_add_4_17 (.A0(b2_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b2_reg[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n13417), .S0(b_s[15]), .S1(b_s[16]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(96[30:59])
    defparam _add_1_358_add_4_17.INIT0 = 16'h5555;
    defparam _add_1_358_add_4_17.INIT1 = 16'h5555;
    defparam _add_1_358_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_358_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13827), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13419), .S1(n161_adj_2002));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_502_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_3 (.A0(n161_adj_2129), .B0(n13827), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_2128), .B1(n13827), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13419), .COUT(n13420), .S0(n158_adj_2001), 
          .S1(n155_adj_2000));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_5 (.A0(n155_adj_2127), .B0(n13827), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_2126), .B1(n13827), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13420), .COUT(n13421), .S0(n152_adj_1999), 
          .S1(n149_adj_1998));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_7 (.A0(n149_adj_2125), .B0(n13827), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_2124), .B1(n13827), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13421), .COUT(n13422), .S0(n146_adj_1997), 
          .S1(n143_adj_1996));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_9 (.A0(n143_adj_2123), .B0(n13827), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_2122), .B1(n13827), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13422), .COUT(n13423), .S0(n140_adj_1995), 
          .S1(n137_adj_1994));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_11 (.A0(n137_adj_2121), .B0(n13827), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_2120), .B1(n13827), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13423), .COUT(n13424), .S0(n134_adj_1993), 
          .S1(n131_adj_1992));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_13 (.A0(n131_adj_2119), .B0(n13827), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_2118), .B1(n13827), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13424), .COUT(n13425), .S0(n128_adj_1991), 
          .S1(n125_adj_1990));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_15 (.A0(n125_adj_2117), .B0(n13827), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_2116), .B1(n13827), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13425), .COUT(n13426), .S0(n122_adj_1989), 
          .S1(n119_adj_1988));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_17 (.A0(n119_adj_2115), .B0(n13827), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_2114), .B1(n13827), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13426), .COUT(n13427), .S0(n116_adj_1987), 
          .S1(n113_adj_1986));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_19 (.A0(n113_adj_2113), .B0(n13827), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_2112), .B1(n13827), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13427), .COUT(n13428), .S0(n110_adj_1985), 
          .S1(n107_adj_1984));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_21 (.A0(n107_adj_2111), .B0(n13827), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_2110), .B1(n13827), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13428), .COUT(n13429), .S0(n104_adj_1983), 
          .S1(n101_adj_1982));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_23 (.A0(n101_adj_2109), .B0(n13827), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_2108), .B1(n13827), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13429), .COUT(n13430), .S0(n98_adj_1981), 
          .S1(n95_adj_1980));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_25 (.A0(n95_adj_2107), .B0(n13827), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_2106), .B1(n13827), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13430), .COUT(n13431), .S0(n92_adj_1979), 
          .S1(n89_adj_1978));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_27 (.A0(n89_adj_2105), .B0(n13827), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_2104), .B1(n13827), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13431), .COUT(n13432), .S0(n86_adj_1977), 
          .S1(n83_adj_1976));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_29 (.A0(n83_adj_2103), .B0(n13827), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_2102), .B1(n13827), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13432), .COUT(n13433), .S0(n80_adj_1975), 
          .S1(n77_adj_1974));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_31 (.A0(n77_adj_2101), .B0(n13827), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_2100), .B1(n13827), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13433), .COUT(n13434), .S0(n74_adj_1973), 
          .S1(n71_adj_1972));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_502_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_502_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_502_add_4_33 (.A0(n1444), .B0(n13827), .C0(n71_adj_2099), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13434), .S0(n68_adj_1971));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_502_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_502_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_502_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_502_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13827), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13435), .S1(n161_adj_2034));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_499_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_3 (.A0(n161_adj_1651), .B0(n13827), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1650), .B1(n13827), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13435), .COUT(n13436), .S0(n158_adj_2033), 
          .S1(n155_adj_2032));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_5 (.A0(n155_adj_1649), .B0(n13827), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1648), .B1(n13827), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13436), .COUT(n13437), .S0(n152_adj_2031), 
          .S1(n149_adj_2030));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_7 (.A0(n149_adj_1647), .B0(n13827), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1646), .B1(n13827), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13437), .COUT(n13438), .S0(n146_adj_2029), 
          .S1(n143_adj_2028));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_9 (.A0(n143_adj_1645), .B0(n13827), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1644), .B1(n13827), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13438), .COUT(n13439), .S0(n140_adj_2027), 
          .S1(n137_adj_2026));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_11 (.A0(n137_adj_1643), .B0(n13827), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1642), .B1(n13827), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13439), .COUT(n13440), .S0(n134_adj_2025), 
          .S1(n131_adj_2024));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_13 (.A0(n131_adj_1641), .B0(n13827), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1640), .B1(n13827), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13440), .COUT(n13441), .S0(n128_adj_2023), 
          .S1(n125_adj_2022));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_15 (.A0(n125_adj_1639), .B0(n13827), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1638), .B1(n13827), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13441), .COUT(n13442), .S0(n122_adj_2021), 
          .S1(n119_adj_2020));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_17 (.A0(n119_adj_1637), .B0(n13827), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1636), .B1(n13827), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13442), .COUT(n13443), .S0(n116_adj_2019), 
          .S1(n113_adj_2018));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_19 (.A0(n113_adj_1635), .B0(n13827), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1634), .B1(n13827), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13443), .COUT(n13444), .S0(n110_adj_2017), 
          .S1(n107_adj_2016));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_21 (.A0(n107_adj_1633), .B0(n13827), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1632), .B1(n13827), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13444), .COUT(n13445), .S0(n104_adj_2015), 
          .S1(n101_adj_2014));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_23 (.A0(n101_adj_1631), .B0(n13827), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1630), .B1(n13827), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13445), .COUT(n13446), .S0(n98_adj_2013), 
          .S1(n95_adj_2012));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_25 (.A0(n95_adj_1629), .B0(n13827), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1628), .B1(n13827), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13446), .COUT(n13447), .S0(n92_adj_2011), 
          .S1(n89_adj_2010));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_27 (.A0(n89_adj_1627), .B0(n13827), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1626), .B1(n13827), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13447), .COUT(n13448), .S0(n86_adj_2009), 
          .S1(n83_adj_2008));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_29 (.A0(n83_adj_1625), .B0(n13827), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1624), .B1(n13827), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13448), .COUT(n13449), .S0(n80_adj_2007), 
          .S1(n77_adj_2006));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_31 (.A0(n77_adj_1623), .B0(n13827), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1622), .B1(n13827), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13449), .COUT(n13450), .S0(n74_adj_2005), 
          .S1(n71_adj_2004));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_499_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_499_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_499_add_4_33 (.A0(n1444), .B0(n13827), .C0(n71_adj_1621), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13450), .S0(n68_adj_2003));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_499_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_499_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_499_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_499_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n1410), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n13454));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_484_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_484_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_3 (.A0(det_q4_28[0]), .B0(n1410), .C0(n161_adj_2161), 
          .D0(n1844), .A1(n161_adj_889), .B1(n1410), .C1(n158_adj_2160), 
          .D1(n1843), .CIN(n13454), .COUT(n13455), .S0(n161_adj_2065), 
          .S1(n158_adj_2064));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_3.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_3.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_5 (.A0(n158_adj_888), .B0(n1410), .C0(n155_adj_2159), 
          .D0(n1842), .A1(n155_adj_887), .B1(n1410), .C1(n152_adj_2158), 
          .D1(n1841), .CIN(n13455), .COUT(n13456), .S0(n155_adj_2063), 
          .S1(n152_adj_2062));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_5.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_5.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_7 (.A0(n152_adj_886), .B0(n1410), .C0(n149_adj_2157), 
          .D0(n1840), .A1(n149_adj_885), .B1(n1410), .C1(n146_adj_2156), 
          .D1(n1839), .CIN(n13456), .COUT(n13457), .S0(n149_adj_2061), 
          .S1(n146_adj_2060));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_7.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_7.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_9 (.A0(n146_adj_884), .B0(n1410), .C0(n143_adj_2155), 
          .D0(n1838), .A1(n143_adj_883), .B1(n1410), .C1(n140_adj_2154), 
          .D1(n1837), .CIN(n13457), .COUT(n13458), .S0(n143_adj_2059), 
          .S1(n140_adj_2058));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_9.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_9.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_11 (.A0(n140_adj_882), .B0(n1410), .C0(n137_adj_2153), 
          .D0(n1836), .A1(n137_adj_881), .B1(n1410), .C1(n134_adj_2152), 
          .D1(n1835), .CIN(n13458), .COUT(n13459), .S0(n137_adj_2057), 
          .S1(n134_adj_2056));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_11.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_11.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_13 (.A0(n134_adj_880), .B0(n1410), .C0(n131_adj_2151), 
          .D0(n1834), .A1(n131_adj_879), .B1(n1410), .C1(n128_adj_2150), 
          .D1(n1833), .CIN(n13459), .COUT(n13460), .S0(n131_adj_2055), 
          .S1(n128_adj_2054));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_13.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_13.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_15 (.A0(n128_adj_878), .B0(n1410), .C0(n125_adj_2149), 
          .D0(n1832), .A1(n125_adj_877), .B1(n1410), .C1(n122_adj_2148), 
          .D1(n1831), .CIN(n13460), .COUT(n13461), .S0(n125_adj_2053), 
          .S1(n122_adj_2052));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_15.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_15.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_17 (.A0(n122_adj_876), .B0(n1410), .C0(n119_adj_2147), 
          .D0(n1830), .A1(n119_adj_875), .B1(n1410), .C1(n116_adj_2146), 
          .D1(n1829), .CIN(n13461), .COUT(n13462), .S0(n119_adj_2051), 
          .S1(n116_adj_2050));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_17.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_17.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_19 (.A0(n116_adj_874), .B0(n1410), .C0(n113_adj_2145), 
          .D0(n1828), .A1(n113_adj_873), .B1(n1410), .C1(n110_adj_2144), 
          .D1(n1827), .CIN(n13462), .COUT(n13463), .S0(n113_adj_2049), 
          .S1(n110_adj_2048));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_19.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_19.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_21 (.A0(n110_adj_872), .B0(n1410), .C0(n107_adj_2143), 
          .D0(n1826), .A1(n107_adj_871), .B1(n1410), .C1(n104_adj_2142), 
          .D1(n1825), .CIN(n13463), .COUT(n13464), .S0(n107_adj_2047), 
          .S1(n104_adj_2046));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_21.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_21.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_23 (.A0(n104_adj_870), .B0(n1410), .C0(n101_adj_2141), 
          .D0(n1824), .A1(n101_adj_869), .B1(n1410), .C1(n98_adj_2140), 
          .D1(n1823), .CIN(n13464), .COUT(n13465), .S0(n101_adj_2045), 
          .S1(n98_adj_2044));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_23.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_23.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_25 (.A0(n98_adj_868), .B0(n1410), .C0(n95_adj_2139), 
          .D0(n1822), .A1(n95_adj_867), .B1(n1410), .C1(n92_adj_2138), 
          .D1(n1821), .CIN(n13465), .COUT(n13466), .S0(n95_adj_2043), 
          .S1(n92_adj_2042));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_25.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_25.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_27 (.A0(n92_adj_866), .B0(n1410), .C0(n89_adj_2137), 
          .D0(n1820), .A1(n89_adj_865), .B1(n1410), .C1(n86_adj_2136), 
          .D1(n1819), .CIN(n13466), .COUT(n13467), .S0(n89_adj_2041), 
          .S1(n86_adj_2040));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_27.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_27.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_29 (.A0(n86_adj_864), .B0(n1410), .C0(n83_adj_2135), 
          .D0(n1818), .A1(n83_adj_863), .B1(n1410), .C1(n80_adj_2134), 
          .D1(n1817), .CIN(n13467), .COUT(n13468), .S0(n83_adj_2039), 
          .S1(n80_adj_2038));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_29.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_29.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_31 (.A0(n80_adj_862), .B0(n1410), .C0(n77_adj_2133), 
          .D0(n1816), .A1(n77_adj_861), .B1(n1410), .C1(n74_adj_2132), 
          .D1(n1815), .CIN(n13468), .COUT(n13469), .S0(n77_adj_2037), 
          .S1(n74_adj_2036));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_31.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_31.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_484_add_4_33 (.A0(n74_adj_860), .B0(n1410), .C0(n71_adj_2131), 
          .D0(n1814), .A1(n71_adj_859), .B1(n1410), .C1(n68_adj_2130), 
          .D1(n1813), .CIN(n13469), .S0(n71_adj_2035), .S1(n1846));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_484_add_4_33.INIT0 = 16'h74b8;
    defparam _add_1_484_add_4_33.INIT1 = 16'h74b8;
    defparam _add_1_484_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_484_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13834), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13471), .S1(n161_adj_2097));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_403_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_3 (.A0(n161_adj_1461), .B0(n13834), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1460), .B1(n13834), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13471), .COUT(n13472), .S0(n158_adj_2096), 
          .S1(n155_adj_2095));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_5 (.A0(n155_adj_1459), .B0(n13834), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1458), .B1(n13834), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13472), .COUT(n13473), .S0(n152_adj_2094), 
          .S1(n149_adj_2093));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_7 (.A0(n149_adj_1457), .B0(n13834), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1456), .B1(n13834), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13473), .COUT(n13474), .S0(n146_adj_2092), 
          .S1(n143_adj_2091));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_9 (.A0(n143_adj_1455), .B0(n13834), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1454), .B1(n13834), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13474), .COUT(n13475), .S0(n140_adj_2090), 
          .S1(n137_adj_2089));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_11 (.A0(n137_adj_1453), .B0(n13834), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1452), .B1(n13834), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13475), .COUT(n13476), .S0(n134_adj_2088), 
          .S1(n131_adj_2087));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_13 (.A0(n131_adj_1451), .B0(n13834), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1450), .B1(n13834), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13476), .COUT(n13477), .S0(n128_adj_2086), 
          .S1(n125_adj_2085));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_15 (.A0(n125_adj_1449), .B0(n13834), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1448), .B1(n13834), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13477), .COUT(n13478), .S0(n122_adj_2084), 
          .S1(n119_adj_2083));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_17 (.A0(n119_adj_1447), .B0(n13834), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1446), .B1(n13834), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13478), .COUT(n13479), .S0(n116_adj_2082), 
          .S1(n113_adj_2081));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_19 (.A0(n113_adj_1445), .B0(n13834), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1444), .B1(n13834), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13479), .COUT(n13480), .S0(n110_adj_2080), 
          .S1(n107_adj_2079));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_21 (.A0(n107_adj_1443), .B0(n13834), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1442), .B1(n13834), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13480), .COUT(n13481), .S0(n104_adj_2078), 
          .S1(n101_adj_2077));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_23 (.A0(n101_adj_1441), .B0(n13834), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1440), .B1(n13834), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13481), .COUT(n13482), .S0(n98_adj_2076), 
          .S1(n95_adj_2075));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_25 (.A0(n95_adj_1439), .B0(n13834), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1438), .B1(n13834), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13482), .COUT(n13483), .S0(n92_adj_2074), 
          .S1(n89_adj_2073));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_27 (.A0(n89_adj_1437), .B0(n13834), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1436), .B1(n13834), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13483), .COUT(n13484), .S0(n86_adj_2072), 
          .S1(n83_adj_2071));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_29 (.A0(n83_adj_1435), .B0(n13834), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1434), .B1(n13834), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13484), .COUT(n13485), .S0(n80_adj_2070), 
          .S1(n77_adj_2069));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_31 (.A0(n77_adj_1433), .B0(n13834), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1432), .B1(n13834), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13485), .COUT(n13486), .S0(n74_adj_2068), 
          .S1(n71_adj_2067));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_403_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_403_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_403_add_4_33 (.A0(n1444), .B0(n13834), .C0(n71_adj_1431), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13486), .S0(n68_adj_2066));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_403_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_403_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_403_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_403_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13828), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13487), .S1(n161_adj_2129));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_496_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_3 (.A0(n161_adj_1272), .B0(n13828), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1779), .B1(n13828), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13487), .COUT(n13488), .S0(n158_adj_2128), 
          .S1(n155_adj_2127));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_5 (.A0(n155_adj_1778), .B0(n13828), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1777), .B1(n13828), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13488), .COUT(n13489), .S0(n152_adj_2126), 
          .S1(n149_adj_2125));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_7 (.A0(n149_adj_1776), .B0(n13828), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1775), .B1(n13828), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13489), .COUT(n13490), .S0(n146_adj_2124), 
          .S1(n143_adj_2123));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_9 (.A0(n143_adj_1774), .B0(n13828), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1773), .B1(n13828), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13490), .COUT(n13491), .S0(n140_adj_2122), 
          .S1(n137_adj_2121));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_11 (.A0(n137_adj_1772), .B0(n13828), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1771), .B1(n13828), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13491), .COUT(n13492), .S0(n134_adj_2120), 
          .S1(n131_adj_2119));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_13 (.A0(n131_adj_1770), .B0(n13828), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1769), .B1(n13828), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13492), .COUT(n13493), .S0(n128_adj_2118), 
          .S1(n125_adj_2117));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_15 (.A0(n125_adj_1768), .B0(n13828), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1767), .B1(n13828), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13493), .COUT(n13494), .S0(n122_adj_2116), 
          .S1(n119_adj_2115));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_17 (.A0(n119_adj_1766), .B0(n13828), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1765), .B1(n13828), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13494), .COUT(n13495), .S0(n116_adj_2114), 
          .S1(n113_adj_2113));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_19 (.A0(n113_adj_1764), .B0(n13828), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1763), .B1(n13828), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13495), .COUT(n13496), .S0(n110_adj_2112), 
          .S1(n107_adj_2111));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_21 (.A0(n107_adj_1762), .B0(n13828), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1761), .B1(n13828), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13496), .COUT(n13497), .S0(n104_adj_2110), 
          .S1(n101_adj_2109));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_23 (.A0(n101_adj_1760), .B0(n13828), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1759), .B1(n13828), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13497), .COUT(n13498), .S0(n98_adj_2108), 
          .S1(n95_adj_2107));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_25 (.A0(n95_adj_1758), .B0(n13828), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1757), .B1(n13828), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13498), .COUT(n13499), .S0(n92_adj_2106), 
          .S1(n89_adj_2105));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_27 (.A0(n89_adj_1756), .B0(n13828), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1755), .B1(n13828), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13499), .COUT(n13500), .S0(n86_adj_2104), 
          .S1(n83_adj_2103));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_29 (.A0(n83_adj_1754), .B0(n13828), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1753), .B1(n13828), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13500), .COUT(n13501), .S0(n80_adj_2102), 
          .S1(n77_adj_2101));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_31 (.A0(n77_adj_1752), .B0(n13828), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1751), .B1(n13828), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13501), .COUT(n13502), .S0(n74_adj_2100), 
          .S1(n71_adj_2099));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_496_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_496_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_496_add_4_33 (.A0(n1444), .B0(n13828), .C0(n71_adj_1750), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13502), .S0(n68_adj_2098));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_496_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_496_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_496_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_496_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13836), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13503), .S1(n161_adj_2161));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_481_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_3 (.A0(n161_adj_921), .B0(n13836), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_920), .B1(n13836), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13503), .COUT(n13504), .S0(n158_adj_2160), 
          .S1(n155_adj_2159));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_5 (.A0(n155_adj_919), .B0(n13836), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_918), .B1(n13836), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13504), .COUT(n13505), .S0(n152_adj_2158), 
          .S1(n149_adj_2157));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_7 (.A0(n149_adj_917), .B0(n13836), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_916), .B1(n13836), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13505), .COUT(n13506), .S0(n146_adj_2156), 
          .S1(n143_adj_2155));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_9 (.A0(n143_adj_915), .B0(n13836), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_914), .B1(n13836), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13506), .COUT(n13507), .S0(n140_adj_2154), 
          .S1(n137_adj_2153));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_11 (.A0(n137_adj_913), .B0(n13836), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_912), .B1(n13836), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13507), .COUT(n13508), .S0(n134_adj_2152), 
          .S1(n131_adj_2151));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_13 (.A0(n131_adj_911), .B0(n13836), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_910), .B1(n13836), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13508), .COUT(n13509), .S0(n128_adj_2150), 
          .S1(n125_adj_2149));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_15 (.A0(n125_adj_909), .B0(n13836), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_908), .B1(n13836), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13509), .COUT(n13510), .S0(n122_adj_2148), 
          .S1(n119_adj_2147));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_17 (.A0(n119_adj_907), .B0(n13836), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_906), .B1(n13836), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13510), .COUT(n13511), .S0(n116_adj_2146), 
          .S1(n113_adj_2145));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_19 (.A0(n113_adj_905), .B0(n13836), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_904), .B1(n13836), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13511), .COUT(n13512), .S0(n110_adj_2144), 
          .S1(n107_adj_2143));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_21 (.A0(n107_adj_903), .B0(n13836), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_902), .B1(n13836), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13512), .COUT(n13513), .S0(n104_adj_2142), 
          .S1(n101_adj_2141));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_23 (.A0(n101_adj_901), .B0(n13836), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_900), .B1(n13836), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13513), .COUT(n13514), .S0(n98_adj_2140), 
          .S1(n95_adj_2139));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_25 (.A0(n95_adj_899), .B0(n13836), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_898), .B1(n13836), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13514), .COUT(n13515), .S0(n92_adj_2138), 
          .S1(n89_adj_2137));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_27 (.A0(n89_adj_897), .B0(n13836), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_896), .B1(n13836), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13515), .COUT(n13516), .S0(n86_adj_2136), 
          .S1(n83_adj_2135));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_29 (.A0(n83_adj_895), .B0(n13836), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_894), .B1(n13836), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13516), .COUT(n13517), .S0(n80_adj_2134), 
          .S1(n77_adj_2133));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_31 (.A0(n77_adj_893), .B0(n13836), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_892), .B1(n13836), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13517), .COUT(n13518), .S0(n74_adj_2132), 
          .S1(n71_adj_2131));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_481_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_481_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_481_add_4_33 (.A0(n1444), .B0(n13836), .C0(n71_adj_891), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13518), .S0(n68_adj_2130));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_481_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_481_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_481_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_481_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13834), .C1(det_q4_28[1]), 
          .D1(n1475), .COUT(n13519), .S1(n161_adj_2193));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_406_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_3 (.A0(n161_adj_1429), .B0(n13834), .C0(det_q4_28[2]), 
          .D0(n1474), .A1(n158_adj_1428), .B1(n13834), .C1(det_q4_28[3]), 
          .D1(n1473), .CIN(n13519), .COUT(n13520), .S0(n158_adj_2192), 
          .S1(n155_adj_2191));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_5 (.A0(n155_adj_1427), .B0(n13834), .C0(det_q4_28[4]), 
          .D0(n1472), .A1(n152_adj_1426), .B1(n13834), .C1(det_q4_28[5]), 
          .D1(n1471), .CIN(n13520), .COUT(n13521), .S0(n152_adj_2190), 
          .S1(n149_adj_2189));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_7 (.A0(n149_adj_1425), .B0(n13834), .C0(det_q4_28[6]), 
          .D0(n1470), .A1(n146_adj_1424), .B1(n13834), .C1(det_q4_28[7]), 
          .D1(n1469), .CIN(n13521), .COUT(n13522), .S0(n146_adj_2188), 
          .S1(n143_adj_2187));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_9 (.A0(n143_adj_1423), .B0(n13834), .C0(det_q4_28[8]), 
          .D0(n1468), .A1(n140_adj_1422), .B1(n13834), .C1(det_q4_28[9]), 
          .D1(n1467), .CIN(n13522), .COUT(n13523), .S0(n140_adj_2186), 
          .S1(n137_adj_2185));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_11 (.A0(n137_adj_1421), .B0(n13834), .C0(det_q4_28[10]), 
          .D0(n1466), .A1(n134_adj_1420), .B1(n13834), .C1(det_q4_28[11]), 
          .D1(n1465), .CIN(n13523), .COUT(n13524), .S0(n134_adj_2184), 
          .S1(n131_adj_2183));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_13 (.A0(n131_adj_1419), .B0(n13834), .C0(det_q4_28[12]), 
          .D0(n1464), .A1(n128_adj_1418), .B1(n13834), .C1(det_q4_28[13]), 
          .D1(n1463), .CIN(n13524), .COUT(n13525), .S0(n128_adj_2182), 
          .S1(n125_adj_2181));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_15 (.A0(n125_adj_1417), .B0(n13834), .C0(det_q4_28[14]), 
          .D0(n1462), .A1(n122_adj_1416), .B1(n13834), .C1(det_q4_28[15]), 
          .D1(n1461), .CIN(n13525), .COUT(n13526), .S0(n122_adj_2180), 
          .S1(n119_adj_2179));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_17 (.A0(n119_adj_1415), .B0(n13834), .C0(det_q4_28[16]), 
          .D0(n1460), .A1(n116_adj_1414), .B1(n13834), .C1(det_q4_28[17]), 
          .D1(n1459), .CIN(n13526), .COUT(n13527), .S0(n116_adj_2178), 
          .S1(n113_adj_2177));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_19 (.A0(n113_adj_1413), .B0(n13834), .C0(det_q4_28[18]), 
          .D0(n1458), .A1(n110_adj_1412), .B1(n13834), .C1(det_q4_28[19]), 
          .D1(n1457), .CIN(n13527), .COUT(n13528), .S0(n110_adj_2176), 
          .S1(n107_adj_2175));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_21 (.A0(n107_adj_1411), .B0(n13834), .C0(det_q4_28[20]), 
          .D0(n1456), .A1(n104_adj_1410), .B1(n13834), .C1(det_q4_28[21]), 
          .D1(n1455), .CIN(n13528), .COUT(n13529), .S0(n104_adj_2174), 
          .S1(n101_adj_2173));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_23 (.A0(n101_adj_1409), .B0(n13834), .C0(det_q4_28[22]), 
          .D0(n1454), .A1(n98_adj_1408), .B1(n13834), .C1(det_q4_28[23]), 
          .D1(n1453), .CIN(n13529), .COUT(n13530), .S0(n98_adj_2172), 
          .S1(n95_adj_2171));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_25 (.A0(n95_adj_1407), .B0(n13834), .C0(det_q4_28[24]), 
          .D0(n1452), .A1(n92_adj_1406), .B1(n13834), .C1(det_q4_28[25]), 
          .D1(n1451), .CIN(n13530), .COUT(n13531), .S0(n92_adj_2170), 
          .S1(n89_adj_2169));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_27 (.A0(n89_adj_1405), .B0(n13834), .C0(det_q4_28[26]), 
          .D0(n1450), .A1(n86_adj_1404), .B1(n13834), .C1(det_q4_28[27]), 
          .D1(n1449), .CIN(n13531), .COUT(n13532), .S0(n86_adj_2168), 
          .S1(n83_adj_2167));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_29 (.A0(n83_adj_1403), .B0(n13834), .C0(det_q4_28[28]), 
          .D0(n1448), .A1(n80_adj_1402), .B1(n13834), .C1(det_q4_28[29]), 
          .D1(n1447), .CIN(n13532), .COUT(n13533), .S0(n80_adj_2166), 
          .S1(n77_adj_2165));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_31 (.A0(n77_adj_1401), .B0(n13834), .C0(det_q4_28[30]), 
          .D0(n1446), .A1(n74_adj_1400), .B1(n13834), .C1(det_q4_28[31]), 
          .D1(n1445), .CIN(n13533), .COUT(n13534), .S0(n74_adj_2164), 
          .S1(n71_adj_2163));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_406_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_406_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_406_add_4_33 (.A0(n1444), .B0(n13834), .C0(n71_adj_1399), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13534), .S0(n68_adj_2162));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_406_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_406_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_406_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_406_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28_31__N_129[0]), .B1(det_q4_28_31__N_97[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n13535), .S1(det_q4_28_31__N_65[0]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_352_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_4 (.A0(det_q4_28_31__N_129[1]), .B0(det_q4_28_31__N_97[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[2]), .B1(det_q4_28_31__N_97[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13535), .COUT(n13536), .S0(det_q4_28_31__N_65[1]), 
          .S1(det_q4_28_31__N_65[2]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_6 (.A0(det_q4_28_31__N_129[3]), .B0(det_q4_28_31__N_97[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[4]), .B1(det_q4_28_31__N_97[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13536), .COUT(n13537), .S0(det_q4_28_31__N_65[3]), 
          .S1(det_q4_28_31__N_65[4]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_8 (.A0(det_q4_28_31__N_129[5]), .B0(det_q4_28_31__N_97[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[6]), .B1(det_q4_28_31__N_97[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13537), .COUT(n13538), .S0(det_q4_28_31__N_65[5]), 
          .S1(det_q4_28_31__N_65[6]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_10 (.A0(det_q4_28_31__N_129[7]), .B0(det_q4_28_31__N_97[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[8]), .B1(det_q4_28_31__N_97[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13538), .COUT(n13539), .S0(det_q4_28_31__N_65[7]), 
          .S1(det_q4_28_31__N_65[8]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_12 (.A0(det_q4_28_31__N_129[9]), .B0(det_q4_28_31__N_97[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[10]), .B1(det_q4_28_31__N_97[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13539), .COUT(n13540), .S0(det_q4_28_31__N_65[9]), 
          .S1(det_q4_28_31__N_65[10]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_14 (.A0(det_q4_28_31__N_129[11]), .B0(det_q4_28_31__N_97[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[12]), .B1(det_q4_28_31__N_97[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13540), .COUT(n13541), .S0(det_q4_28_31__N_65[11]), 
          .S1(det_q4_28_31__N_65[12]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_16 (.A0(det_q4_28_31__N_129[13]), .B0(det_q4_28_31__N_97[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[14]), .B1(det_q4_28_31__N_97[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13541), .COUT(n13542), .S0(det_q4_28_31__N_65[13]), 
          .S1(det_q4_28_31__N_65[14]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_18 (.A0(det_q4_28_31__N_129[15]), .B0(det_q4_28_31__N_97[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[16]), .B1(det_q4_28_31__N_97[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13542), .COUT(n13543), .S0(det_q4_28_31__N_65[15]), 
          .S1(det_q4_28_31__N_65[16]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_20 (.A0(det_q4_28_31__N_129[17]), .B0(det_q4_28_31__N_97[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[18]), .B1(det_q4_28_31__N_97[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13543), .COUT(n13544), .S0(det_q4_28_31__N_65[17]), 
          .S1(det_q4_28_31__N_65[18]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_22 (.A0(det_q4_28_31__N_129[19]), .B0(det_q4_28_31__N_97[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[20]), .B1(det_q4_28_31__N_97[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13544), .COUT(n13545), .S0(det_q4_28_31__N_65[19]), 
          .S1(det_q4_28_31__N_65[20]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_24 (.A0(det_q4_28_31__N_129[21]), .B0(det_q4_28_31__N_97[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[22]), .B1(det_q4_28_31__N_97[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13545), .COUT(n13546), .S0(det_q4_28_31__N_65[21]), 
          .S1(det_q4_28_31__N_65[22]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_26 (.A0(det_q4_28_31__N_129[23]), .B0(det_q4_28_31__N_97[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[24]), .B1(det_q4_28_31__N_97[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13546), .COUT(n13547), .S0(det_q4_28_31__N_65[23]), 
          .S1(det_q4_28_31__N_65[24]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_28 (.A0(det_q4_28_31__N_129[25]), .B0(det_q4_28_31__N_97[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[26]), .B1(det_q4_28_31__N_97[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13547), .COUT(n13548), .S0(det_q4_28_31__N_65[25]), 
          .S1(det_q4_28_31__N_65[26]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_30 (.A0(det_q4_28_31__N_129[27]), .B0(det_q4_28_31__N_97[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[28]), .B1(det_q4_28_31__N_97[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13548), .COUT(n13549), .S0(det_q4_28_31__N_65[27]), 
          .S1(det_q4_28_31__N_65[28]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_32 (.A0(det_q4_28_31__N_129[29]), .B0(det_q4_28_31__N_97[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_129[30]), .B1(det_q4_28_31__N_97[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n13549), .COUT(n13550), .S0(det_q4_28_31__N_65[29]), 
          .S1(det_q4_28_31__N_65[30]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_352_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_352_add_4_34 (.A0(det_q4_28_31__N_129[31]), .B0(det_q4_28_31__N_97[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n13550), .S0(det_q4_28_31__N_65[31]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(58[26:43])
    defparam _add_1_352_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_352_add_4_34.INIT1 = 16'h0000;
    defparam _add_1_352_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_352_add_4_34.INJECT1_1 = "NO";
    CCU2C add_807_2 (.A0(prod_c[15]), .B0(prod_c[16]), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n13551));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_2.INIT0 = 16'h0008;
    defparam add_807_2.INIT1 = 16'haaa0;
    defparam add_807_2.INJECT1_0 = "NO";
    defparam add_807_2.INJECT1_1 = "NO";
    CCU2C add_807_4 (.A0(prod_c[18]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[19]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13551), .COUT(n13552));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_4.INIT0 = 16'haaa0;
    defparam add_807_4.INIT1 = 16'haaa0;
    defparam add_807_4.INJECT1_0 = "NO";
    defparam add_807_4.INJECT1_1 = "NO";
    CCU2C add_807_6 (.A0(prod_c[20]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[21]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13552), .COUT(n13553));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_6.INIT0 = 16'haaa0;
    defparam add_807_6.INIT1 = 16'haaa0;
    defparam add_807_6.INJECT1_0 = "NO";
    defparam add_807_6.INJECT1_1 = "NO";
    CCU2C add_807_8 (.A0(prod_c[22]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[23]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13553), .COUT(n13554));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_8.INIT0 = 16'haaa0;
    defparam add_807_8.INIT1 = 16'haaa0;
    defparam add_807_8.INJECT1_0 = "NO";
    defparam add_807_8.INJECT1_1 = "NO";
    CCU2C add_807_10 (.A0(prod_c[24]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[25]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13554), .COUT(n13555));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_10.INIT0 = 16'haaa0;
    defparam add_807_10.INIT1 = 16'haaa0;
    defparam add_807_10.INJECT1_0 = "NO";
    defparam add_807_10.INJECT1_1 = "NO";
    CCU2C add_807_12 (.A0(prod_c[26]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[27]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13555), .COUT(n13556));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_12.INIT0 = 16'haaa0;
    defparam add_807_12.INIT1 = 16'haaa0;
    defparam add_807_12.INJECT1_0 = "NO";
    defparam add_807_12.INJECT1_1 = "NO";
    CCU2C add_807_14 (.A0(prod_c[28]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[29]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13556), .COUT(n13557));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_14.INIT0 = 16'haaa0;
    defparam add_807_14.INIT1 = 16'haaa0;
    defparam add_807_14.INJECT1_0 = "NO";
    defparam add_807_14.INJECT1_1 = "NO";
    CCU2C add_807_16 (.A0(prod_c[30]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[31]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13557), .COUT(n13558));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_16.INIT0 = 16'haaa0;
    defparam add_807_16.INIT1 = 16'haaa0;
    defparam add_807_16.INJECT1_0 = "NO";
    defparam add_807_16.INJECT1_1 = "NO";
    CCU2C add_807_18 (.A0(prod_c[32]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[33]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13558), .COUT(n13559), .S0(c_inv_15__N_33[32]), .S1(c_inv_15__N_33[33]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_18.INIT0 = 16'haaa0;
    defparam add_807_18.INIT1 = 16'haaa0;
    defparam add_807_18.INJECT1_0 = "NO";
    defparam add_807_18.INJECT1_1 = "NO";
    CCU2C add_807_20 (.A0(prod_c[34]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[35]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13559), .COUT(n13560), .S0(c_inv_15__N_33[34]), .S1(c_inv_15__N_33[35]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_20.INIT0 = 16'haaa0;
    defparam add_807_20.INIT1 = 16'haaa0;
    defparam add_807_20.INJECT1_0 = "NO";
    defparam add_807_20.INJECT1_1 = "NO";
    CCU2C add_807_22 (.A0(prod_c[36]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[37]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13560), .COUT(n13561), .S0(c_inv_15__N_33[36]), .S1(c_inv_15__N_33[37]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_22.INIT0 = 16'haaa0;
    defparam add_807_22.INIT1 = 16'haaa0;
    defparam add_807_22.INJECT1_0 = "NO";
    defparam add_807_22.INJECT1_1 = "NO";
    CCU2C add_807_24 (.A0(prod_c[38]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[39]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13561), .COUT(n13562), .S0(c_inv_15__N_33[38]), .S1(c_inv_15__N_33[39]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_24.INIT0 = 16'haaa0;
    defparam add_807_24.INIT1 = 16'haaa0;
    defparam add_807_24.INJECT1_0 = "NO";
    defparam add_807_24.INJECT1_1 = "NO";
    CCU2C add_807_26 (.A0(prod_c[40]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[41]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13562), .COUT(n13563), .S0(c_inv_15__N_33[40]), .S1(c_inv_15__N_33[41]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_26.INIT0 = 16'haaa0;
    defparam add_807_26.INIT1 = 16'haaa0;
    defparam add_807_26.INJECT1_0 = "NO";
    defparam add_807_26.INJECT1_1 = "NO";
    CCU2C add_807_28 (.A0(prod_c[42]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[43]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13563), .COUT(n13564), .S0(c_inv_15__N_33[42]), .S1(c_inv_15__N_33[43]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_28.INIT0 = 16'haaa0;
    defparam add_807_28.INIT1 = 16'haaa0;
    defparam add_807_28.INJECT1_0 = "NO";
    defparam add_807_28.INJECT1_1 = "NO";
    CCU2C add_807_30 (.A0(prod_c[44]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[45]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13564), .COUT(n13565), .S0(c_inv_15__N_33[44]), .S1(c_inv_15__N_33[45]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_30.INIT0 = 16'haaa0;
    defparam add_807_30.INIT1 = 16'haaa0;
    defparam add_807_30.INJECT1_0 = "NO";
    defparam add_807_30.INJECT1_1 = "NO";
    CCU2C add_807_32 (.A0(prod_c[46]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(prod_c[47]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n13565), .S0(c_inv_15__N_33[46]), .S1(c_inv_15__N_33[47]));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(116[19:38])
    defparam add_807_32.INIT0 = 16'haaa0;
    defparam add_807_32.INIT1 = 16'haaa0;
    defparam add_807_32.INJECT1_0 = "NO";
    defparam add_807_32.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module reciprocal_q16_16
//

module reciprocal_q16_16 (n1474, det_q4_28, n13829, n2379, error_recip, 
            clk_c, inv_det_31__N_227, n1465, n13836, n1834, n1464, 
            n1833, n1473, n2378, n1472, n2377, n1471, n2376, n1470, 
            n2375, n1469, n2374, n1468, n2373, n1467, n2372, n1466, 
            n2371, n2370, n2369, n1463, n2368, n1462, n2367, n1461, 
            n2366, n1460, n2365, n1459, n2364, n1458, n2363, n1457, 
            n2362, n1456, n2361, n1455, n2360, n1454, n2359, n1453, 
            n2358, n1452, n2357, n1451, n2356, n1450, n2355, n1449, 
            n2354, n1448, n2353, n1447, n2352, n1832, n1446, n2351, 
            n1445, n2350, n1475, n1844, n1843, n1842, n1841, n1840, 
            n1839, n1838, n1837, n1836, n1835, n1831, n1830, n1829, 
            n1828, n1827, n2382, n46, n1846, n38, n2583, n2616, 
            n1444, n1826, n1825, n1824, n1823, n1822, n1821, n1820, 
            n1819, n1818, n1817, n1816, n1815, n1814, n68, n68_adj_1, 
            n68_adj_2, n64, n63, n13818, n3422, n3424, n3423, 
            n3426, n3425, n3428, n3427, n3430, n3429, n3432, n3431, 
            n3434, n3433, n3436, n3435, n3438, n3437, n3440, n3439, 
            n3442, n3441, n3444, n3443, n3446, n3445, n3448, n3447, 
            n3450, n3449, n3452, n3451, n3454, n3487, n62, n2650, 
            n50, n49, n2449, n47, n2516, n48, GND_net, n2380, 
            VCC_net) /* synthesis syn_module_defined=1 */ ;
    input n1474;
    input [31:0]det_q4_28;
    input n13829;
    output n2379;
    output error_recip;
    input clk_c;
    output inv_det_31__N_227;
    input n1465;
    input n13836;
    output n1834;
    input n1464;
    output n1833;
    input n1473;
    output n2378;
    input n1472;
    output n2377;
    input n1471;
    output n2376;
    input n1470;
    output n2375;
    input n1469;
    output n2374;
    input n1468;
    output n2373;
    input n1467;
    output n2372;
    input n1466;
    output n2371;
    output n2370;
    output n2369;
    input n1463;
    output n2368;
    input n1462;
    output n2367;
    input n1461;
    output n2366;
    input n1460;
    output n2365;
    input n1459;
    output n2364;
    input n1458;
    output n2363;
    input n1457;
    output n2362;
    input n1456;
    output n2361;
    input n1455;
    output n2360;
    input n1454;
    output n2359;
    input n1453;
    output n2358;
    input n1452;
    output n2357;
    input n1451;
    output n2356;
    input n1450;
    output n2355;
    input n1449;
    output n2354;
    input n1448;
    output n2353;
    input n1447;
    output n2352;
    output n1832;
    input n1446;
    output n2351;
    input n1445;
    output n2350;
    input n1475;
    output n1844;
    output n1843;
    output n1842;
    output n1841;
    output n1840;
    output n1839;
    output n1838;
    output n1837;
    output n1836;
    output n1835;
    output n1831;
    output n1830;
    output n1829;
    output n1828;
    output n1827;
    input n2382;
    output n46;
    input n1846;
    output n38;
    input n2583;
    output [31:0]n2616;
    input n1444;
    output n1826;
    output n1825;
    output n1824;
    output n1823;
    output n1822;
    output n1821;
    output n1820;
    output n1819;
    output n1818;
    output n1817;
    output n1816;
    output n1815;
    output n1814;
    input n68;
    input n68_adj_1;
    input n68_adj_2;
    output n64;
    output n63;
    input n13818;
    output n3422;
    output n3424;
    output n3423;
    output n3426;
    output n3425;
    output n3428;
    output n3427;
    output n3430;
    output n3429;
    output n3432;
    output n3431;
    output n3434;
    output n3433;
    output n3436;
    output n3435;
    output n3438;
    output n3437;
    output n3440;
    output n3439;
    output n3442;
    output n3441;
    output n3444;
    output n3443;
    output n3446;
    output n3445;
    output n3448;
    output n3447;
    output n3450;
    output n3449;
    output n3452;
    output n3451;
    input n3454;
    output [31:0]n3487;
    output n62;
    input n2650;
    output n50;
    output n49;
    input n2449;
    output n47;
    input n2516;
    output n48;
    input GND_net;
    output n2380;
    input VCC_net;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/inverterv1.v(16[20:23])
    
    wire n13634, n13633, n13632, n13631;
    
    LUT4 mux_90_i2_3_lut (.A(n1474), .B(det_q4_28[2]), .C(n13829), .Z(n2379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i2_3_lut.init = 16'hcaca;
    FD1S3AX error_10 (.D(inv_det_31__N_227), .CK(clk_c), .Q(error_recip)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=23, LSE_RCOL=6, LSE_LLINE=86, LSE_RLINE=92 */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(24[18] 31[12])
    defparam error_10.GSR = "ENABLED";
    LUT4 mux_74_i11_3_lut (.A(n1465), .B(det_q4_28[11]), .C(n13836), .Z(n1834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i11_3_lut.init = 16'hcaca;
    LUT4 mux_74_i12_3_lut (.A(n1464), .B(det_q4_28[12]), .C(n13836), .Z(n1833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i12_3_lut.init = 16'hcaca;
    LUT4 mux_90_i3_3_lut (.A(n1473), .B(det_q4_28[3]), .C(n13829), .Z(n2378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i3_3_lut.init = 16'hcaca;
    LUT4 mux_90_i4_3_lut (.A(n1472), .B(det_q4_28[4]), .C(n13829), .Z(n2377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i4_3_lut.init = 16'hcaca;
    LUT4 mux_90_i5_3_lut (.A(n1471), .B(det_q4_28[5]), .C(n13829), .Z(n2376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i5_3_lut.init = 16'hcaca;
    LUT4 mux_90_i6_3_lut (.A(n1470), .B(det_q4_28[6]), .C(n13829), .Z(n2375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i6_3_lut.init = 16'hcaca;
    LUT4 mux_90_i7_3_lut (.A(n1469), .B(det_q4_28[7]), .C(n13829), .Z(n2374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i7_3_lut.init = 16'hcaca;
    LUT4 mux_90_i8_3_lut (.A(n1468), .B(det_q4_28[8]), .C(n13829), .Z(n2373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i8_3_lut.init = 16'hcaca;
    LUT4 mux_90_i9_3_lut (.A(n1467), .B(det_q4_28[9]), .C(n13829), .Z(n2372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i9_3_lut.init = 16'hcaca;
    LUT4 mux_90_i10_3_lut (.A(n1466), .B(det_q4_28[10]), .C(n13829), .Z(n2371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i10_3_lut.init = 16'hcaca;
    LUT4 mux_90_i11_3_lut (.A(n1465), .B(det_q4_28[11]), .C(n13829), .Z(n2370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i11_3_lut.init = 16'hcaca;
    LUT4 mux_90_i12_3_lut (.A(n1464), .B(det_q4_28[12]), .C(n13829), .Z(n2369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i12_3_lut.init = 16'hcaca;
    LUT4 mux_90_i13_3_lut (.A(n1463), .B(det_q4_28[13]), .C(n13829), .Z(n2368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i13_3_lut.init = 16'hcaca;
    LUT4 mux_90_i14_3_lut (.A(n1462), .B(det_q4_28[14]), .C(n13829), .Z(n2367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i14_3_lut.init = 16'hcaca;
    LUT4 mux_90_i15_3_lut (.A(n1461), .B(det_q4_28[15]), .C(n13829), .Z(n2366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i15_3_lut.init = 16'hcaca;
    LUT4 mux_90_i16_3_lut (.A(n1460), .B(det_q4_28[16]), .C(n13829), .Z(n2365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i16_3_lut.init = 16'hcaca;
    LUT4 mux_90_i17_3_lut (.A(n1459), .B(det_q4_28[17]), .C(n13829), .Z(n2364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i17_3_lut.init = 16'hcaca;
    LUT4 mux_90_i18_3_lut (.A(n1458), .B(det_q4_28[18]), .C(n13829), .Z(n2363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i18_3_lut.init = 16'hcaca;
    LUT4 mux_90_i19_3_lut (.A(n1457), .B(det_q4_28[19]), .C(n13829), .Z(n2362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i19_3_lut.init = 16'hcaca;
    LUT4 mux_90_i20_3_lut (.A(n1456), .B(det_q4_28[20]), .C(n13829), .Z(n2361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i20_3_lut.init = 16'hcaca;
    LUT4 mux_90_i21_3_lut (.A(n1455), .B(det_q4_28[21]), .C(n13829), .Z(n2360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i21_3_lut.init = 16'hcaca;
    LUT4 mux_90_i22_3_lut (.A(n1454), .B(det_q4_28[22]), .C(n13829), .Z(n2359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i22_3_lut.init = 16'hcaca;
    LUT4 mux_90_i23_3_lut (.A(n1453), .B(det_q4_28[23]), .C(n13829), .Z(n2358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i23_3_lut.init = 16'hcaca;
    LUT4 mux_90_i24_3_lut (.A(n1452), .B(det_q4_28[24]), .C(n13829), .Z(n2357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i24_3_lut.init = 16'hcaca;
    LUT4 mux_90_i25_3_lut (.A(n1451), .B(det_q4_28[25]), .C(n13829), .Z(n2356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i25_3_lut.init = 16'hcaca;
    LUT4 mux_90_i26_3_lut (.A(n1450), .B(det_q4_28[26]), .C(n13829), .Z(n2355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i26_3_lut.init = 16'hcaca;
    LUT4 mux_90_i27_3_lut (.A(n1449), .B(det_q4_28[27]), .C(n13829), .Z(n2354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i27_3_lut.init = 16'hcaca;
    LUT4 mux_90_i28_3_lut (.A(n1448), .B(det_q4_28[28]), .C(n13829), .Z(n2353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i28_3_lut.init = 16'hcaca;
    LUT4 mux_90_i29_3_lut (.A(n1447), .B(det_q4_28[29]), .C(n13829), .Z(n2352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i29_3_lut.init = 16'hcaca;
    LUT4 mux_74_i13_3_lut (.A(n1463), .B(det_q4_28[13]), .C(n13836), .Z(n1832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i13_3_lut.init = 16'hcaca;
    LUT4 mux_90_i30_3_lut (.A(n1446), .B(det_q4_28[30]), .C(n13829), .Z(n2351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i30_3_lut.init = 16'hcaca;
    LUT4 mux_90_i31_3_lut (.A(n1445), .B(det_q4_28[31]), .C(n13829), .Z(n2350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i31_3_lut.init = 16'hcaca;
    LUT4 mux_74_i1_3_lut (.A(n1475), .B(det_q4_28[1]), .C(n13836), .Z(n1844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i1_3_lut.init = 16'hcaca;
    LUT4 mux_74_i2_3_lut (.A(n1474), .B(det_q4_28[2]), .C(n13836), .Z(n1843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i2_3_lut.init = 16'hcaca;
    LUT4 mux_74_i3_3_lut (.A(n1473), .B(det_q4_28[3]), .C(n13836), .Z(n1842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i3_3_lut.init = 16'hcaca;
    LUT4 mux_74_i4_3_lut (.A(n1472), .B(det_q4_28[4]), .C(n13836), .Z(n1841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i4_3_lut.init = 16'hcaca;
    LUT4 mux_74_i5_3_lut (.A(n1471), .B(det_q4_28[5]), .C(n13836), .Z(n1840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i5_3_lut.init = 16'hcaca;
    LUT4 mux_74_i6_3_lut (.A(n1470), .B(det_q4_28[6]), .C(n13836), .Z(n1839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i6_3_lut.init = 16'hcaca;
    LUT4 mux_74_i7_3_lut (.A(n1469), .B(det_q4_28[7]), .C(n13836), .Z(n1838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i7_3_lut.init = 16'hcaca;
    LUT4 mux_74_i8_3_lut (.A(n1468), .B(det_q4_28[8]), .C(n13836), .Z(n1837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i8_3_lut.init = 16'hcaca;
    LUT4 mux_74_i9_3_lut (.A(n1467), .B(det_q4_28[9]), .C(n13836), .Z(n1836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i9_3_lut.init = 16'hcaca;
    LUT4 mux_74_i10_3_lut (.A(n1466), .B(det_q4_28[10]), .C(n13836), .Z(n1835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i10_3_lut.init = 16'hcaca;
    LUT4 mux_74_i14_3_lut (.A(n1462), .B(det_q4_28[14]), .C(n13836), .Z(n1831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i14_3_lut.init = 16'hcaca;
    LUT4 mux_74_i15_3_lut (.A(n1461), .B(det_q4_28[15]), .C(n13836), .Z(n1830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i15_3_lut.init = 16'hcaca;
    LUT4 mux_74_i16_3_lut (.A(n1460), .B(det_q4_28[16]), .C(n13836), .Z(n1829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i16_3_lut.init = 16'hcaca;
    LUT4 mux_74_i17_3_lut (.A(n1459), .B(det_q4_28[17]), .C(n13836), .Z(n1828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i17_3_lut.init = 16'hcaca;
    LUT4 mux_74_i18_3_lut (.A(n1458), .B(det_q4_28[18]), .C(n13836), .Z(n1827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i18_3_lut.init = 16'hcaca;
    LUT4 i1540_2_lut (.A(n2382), .B(inv_det_31__N_227), .Z(n46)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1540_2_lut.init = 16'h1111;
    LUT4 i1564_2_lut (.A(n1846), .B(inv_det_31__N_227), .Z(n38)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1564_2_lut.init = 16'h1111;
    LUT4 mux_98_i31_3_lut (.A(n1445), .B(det_q4_28[31]), .C(n2583), .Z(n2616[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i31_3_lut.init = 16'hcaca;
    LUT4 i710_2_lut (.A(n1444), .B(n2583), .Z(n2616[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i710_2_lut.init = 16'h2222;
    LUT4 mux_98_i29_3_lut (.A(n1447), .B(det_q4_28[29]), .C(n2583), .Z(n2616[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i29_3_lut.init = 16'hcaca;
    LUT4 mux_74_i19_3_lut (.A(n1457), .B(det_q4_28[19]), .C(n13836), .Z(n1826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i19_3_lut.init = 16'hcaca;
    LUT4 mux_74_i20_3_lut (.A(n1456), .B(det_q4_28[20]), .C(n13836), .Z(n1825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i20_3_lut.init = 16'hcaca;
    LUT4 mux_74_i21_3_lut (.A(n1455), .B(det_q4_28[21]), .C(n13836), .Z(n1824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i21_3_lut.init = 16'hcaca;
    LUT4 mux_74_i22_3_lut (.A(n1454), .B(det_q4_28[22]), .C(n13836), .Z(n1823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i22_3_lut.init = 16'hcaca;
    LUT4 mux_74_i23_3_lut (.A(n1453), .B(det_q4_28[23]), .C(n13836), .Z(n1822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i23_3_lut.init = 16'hcaca;
    LUT4 mux_74_i24_3_lut (.A(n1452), .B(det_q4_28[24]), .C(n13836), .Z(n1821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i24_3_lut.init = 16'hcaca;
    LUT4 mux_74_i25_3_lut (.A(n1451), .B(det_q4_28[25]), .C(n13836), .Z(n1820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i25_3_lut.init = 16'hcaca;
    LUT4 mux_74_i26_3_lut (.A(n1450), .B(det_q4_28[26]), .C(n13836), .Z(n1819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i26_3_lut.init = 16'hcaca;
    LUT4 mux_74_i27_3_lut (.A(n1449), .B(det_q4_28[27]), .C(n13836), .Z(n1818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i27_3_lut.init = 16'hcaca;
    LUT4 mux_74_i28_3_lut (.A(n1448), .B(det_q4_28[28]), .C(n13836), .Z(n1817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i28_3_lut.init = 16'hcaca;
    LUT4 mux_74_i29_3_lut (.A(n1447), .B(det_q4_28[29]), .C(n13836), .Z(n1816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i29_3_lut.init = 16'hcaca;
    LUT4 mux_74_i30_3_lut (.A(n1446), .B(det_q4_28[30]), .C(n13836), .Z(n1815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i30_3_lut.init = 16'hcaca;
    LUT4 mux_74_i31_3_lut (.A(n1445), .B(det_q4_28[31]), .C(n13836), .Z(n1814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_74_i31_3_lut.init = 16'hcaca;
    LUT4 i1483_4_lut (.A(n68), .B(inv_det_31__N_227), .C(n68_adj_1), .D(n68_adj_2), 
         .Z(n64)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+(C (D))))) */ ;
    defparam i1483_4_lut.init = 16'h0311;
    LUT4 i1489_2_lut (.A(n68_adj_2), .B(inv_det_31__N_227), .Z(n63)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1489_2_lut.init = 16'h1111;
    LUT4 mux_98_i30_3_lut (.A(n1446), .B(det_q4_28[30]), .C(n2583), .Z(n2616[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i30_3_lut.init = 16'hcaca;
    LUT4 mux_98_i27_3_lut (.A(n1449), .B(det_q4_28[27]), .C(n2583), .Z(n2616[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i27_3_lut.init = 16'hcaca;
    LUT4 mux_98_i28_3_lut (.A(n1448), .B(det_q4_28[28]), .C(n2583), .Z(n2616[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i28_3_lut.init = 16'hcaca;
    LUT4 mux_98_i25_3_lut (.A(n1451), .B(det_q4_28[25]), .C(n2583), .Z(n2616[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i25_3_lut.init = 16'hcaca;
    LUT4 mux_98_i26_3_lut (.A(n1450), .B(det_q4_28[26]), .C(n2583), .Z(n2616[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i26_3_lut.init = 16'hcaca;
    LUT4 mux_98_i23_3_lut (.A(n1453), .B(det_q4_28[23]), .C(n2583), .Z(n2616[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i23_3_lut.init = 16'hcaca;
    LUT4 mux_98_i24_3_lut (.A(n1452), .B(det_q4_28[24]), .C(n2583), .Z(n2616[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i24_3_lut.init = 16'hcaca;
    LUT4 mux_98_i21_3_lut (.A(n1455), .B(det_q4_28[21]), .C(n2583), .Z(n2616[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i21_3_lut.init = 16'hcaca;
    LUT4 mux_98_i22_3_lut (.A(n1454), .B(det_q4_28[22]), .C(n2583), .Z(n2616[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i22_3_lut.init = 16'hcaca;
    LUT4 mux_98_i19_3_lut (.A(n1457), .B(det_q4_28[19]), .C(n2583), .Z(n2616[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i19_3_lut.init = 16'hcaca;
    LUT4 mux_98_i20_3_lut (.A(n1456), .B(det_q4_28[20]), .C(n2583), .Z(n2616[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i20_3_lut.init = 16'hcaca;
    LUT4 mux_98_i17_3_lut (.A(n1459), .B(det_q4_28[17]), .C(n2583), .Z(n2616[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i17_3_lut.init = 16'hcaca;
    LUT4 mux_98_i18_3_lut (.A(n1458), .B(det_q4_28[18]), .C(n2583), .Z(n2616[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i18_3_lut.init = 16'hcaca;
    LUT4 mux_98_i15_3_lut (.A(n1461), .B(det_q4_28[15]), .C(n2583), .Z(n2616[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i15_3_lut.init = 16'hcaca;
    LUT4 mux_98_i16_3_lut (.A(n1460), .B(det_q4_28[16]), .C(n2583), .Z(n2616[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i16_3_lut.init = 16'hcaca;
    LUT4 mux_98_i13_3_lut (.A(n1463), .B(det_q4_28[13]), .C(n2583), .Z(n2616[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i13_3_lut.init = 16'hcaca;
    LUT4 mux_98_i14_3_lut (.A(n1462), .B(det_q4_28[14]), .C(n2583), .Z(n2616[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i14_3_lut.init = 16'hcaca;
    LUT4 mux_98_i11_3_lut (.A(n1465), .B(det_q4_28[11]), .C(n2583), .Z(n2616[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i11_3_lut.init = 16'hcaca;
    LUT4 mux_98_i12_3_lut (.A(n1464), .B(det_q4_28[12]), .C(n2583), .Z(n2616[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i12_3_lut.init = 16'hcaca;
    LUT4 mux_98_i9_3_lut (.A(n1467), .B(det_q4_28[9]), .C(n2583), .Z(n2616[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i9_3_lut.init = 16'hcaca;
    LUT4 mux_98_i10_3_lut (.A(n1466), .B(det_q4_28[10]), .C(n2583), .Z(n2616[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i10_3_lut.init = 16'hcaca;
    LUT4 mux_98_i7_3_lut (.A(n1469), .B(det_q4_28[7]), .C(n2583), .Z(n2616[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i7_3_lut.init = 16'hcaca;
    LUT4 mux_98_i8_3_lut (.A(n1468), .B(det_q4_28[8]), .C(n2583), .Z(n2616[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i8_3_lut.init = 16'hcaca;
    LUT4 mux_98_i5_3_lut (.A(n1471), .B(det_q4_28[5]), .C(n2583), .Z(n2616[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i5_3_lut.init = 16'hcaca;
    LUT4 mux_98_i6_3_lut (.A(n1470), .B(det_q4_28[6]), .C(n2583), .Z(n2616[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i6_3_lut.init = 16'hcaca;
    LUT4 mux_98_i3_3_lut (.A(n1473), .B(det_q4_28[3]), .C(n2583), .Z(n2616[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i3_3_lut.init = 16'hcaca;
    LUT4 mux_98_i4_3_lut (.A(n1472), .B(det_q4_28[4]), .C(n2583), .Z(n2616[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i4_3_lut.init = 16'hcaca;
    LUT4 mux_98_i1_3_lut (.A(n1475), .B(det_q4_28[1]), .C(n2583), .Z(n2616[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i1_3_lut.init = 16'hcaca;
    LUT4 mux_98_i2_3_lut (.A(n1474), .B(det_q4_28[2]), .C(n2583), .Z(n2616[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_98_i2_3_lut.init = 16'hcaca;
    LUT4 mux_122_i31_3_lut (.A(n1445), .B(det_q4_28[31]), .C(n13818), 
         .Z(n3422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i31_3_lut.init = 16'hcaca;
    LUT4 mux_122_i29_3_lut (.A(n1447), .B(det_q4_28[29]), .C(n13818), 
         .Z(n3424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i29_3_lut.init = 16'hcaca;
    LUT4 mux_122_i30_3_lut (.A(n1446), .B(det_q4_28[30]), .C(n13818), 
         .Z(n3423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i30_3_lut.init = 16'hcaca;
    LUT4 mux_122_i27_3_lut (.A(n1449), .B(det_q4_28[27]), .C(n13818), 
         .Z(n3426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i27_3_lut.init = 16'hcaca;
    LUT4 mux_122_i28_3_lut (.A(n1448), .B(det_q4_28[28]), .C(n13818), 
         .Z(n3425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i28_3_lut.init = 16'hcaca;
    LUT4 mux_122_i25_3_lut (.A(n1451), .B(det_q4_28[25]), .C(n13818), 
         .Z(n3428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i25_3_lut.init = 16'hcaca;
    LUT4 mux_122_i26_3_lut (.A(n1450), .B(det_q4_28[26]), .C(n13818), 
         .Z(n3427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i26_3_lut.init = 16'hcaca;
    LUT4 mux_122_i23_3_lut (.A(n1453), .B(det_q4_28[23]), .C(n13818), 
         .Z(n3430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i23_3_lut.init = 16'hcaca;
    LUT4 mux_122_i24_3_lut (.A(n1452), .B(det_q4_28[24]), .C(n13818), 
         .Z(n3429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i24_3_lut.init = 16'hcaca;
    LUT4 mux_122_i21_3_lut (.A(n1455), .B(det_q4_28[21]), .C(n13818), 
         .Z(n3432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i21_3_lut.init = 16'hcaca;
    LUT4 mux_122_i22_3_lut (.A(n1454), .B(det_q4_28[22]), .C(n13818), 
         .Z(n3431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i22_3_lut.init = 16'hcaca;
    LUT4 mux_122_i19_3_lut (.A(n1457), .B(det_q4_28[19]), .C(n13818), 
         .Z(n3434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i19_3_lut.init = 16'hcaca;
    LUT4 mux_122_i20_3_lut (.A(n1456), .B(det_q4_28[20]), .C(n13818), 
         .Z(n3433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i20_3_lut.init = 16'hcaca;
    LUT4 mux_122_i17_3_lut (.A(n1459), .B(det_q4_28[17]), .C(n13818), 
         .Z(n3436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i17_3_lut.init = 16'hcaca;
    LUT4 mux_122_i18_3_lut (.A(n1458), .B(det_q4_28[18]), .C(n13818), 
         .Z(n3435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i18_3_lut.init = 16'hcaca;
    LUT4 mux_122_i15_3_lut (.A(n1461), .B(det_q4_28[15]), .C(n13818), 
         .Z(n3438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i15_3_lut.init = 16'hcaca;
    LUT4 mux_122_i16_3_lut (.A(n1460), .B(det_q4_28[16]), .C(n13818), 
         .Z(n3437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i16_3_lut.init = 16'hcaca;
    LUT4 mux_122_i13_3_lut (.A(n1463), .B(det_q4_28[13]), .C(n13818), 
         .Z(n3440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i13_3_lut.init = 16'hcaca;
    LUT4 mux_122_i14_3_lut (.A(n1462), .B(det_q4_28[14]), .C(n13818), 
         .Z(n3439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i14_3_lut.init = 16'hcaca;
    LUT4 mux_122_i11_3_lut (.A(n1465), .B(det_q4_28[11]), .C(n13818), 
         .Z(n3442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i11_3_lut.init = 16'hcaca;
    LUT4 mux_122_i12_3_lut (.A(n1464), .B(det_q4_28[12]), .C(n13818), 
         .Z(n3441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i12_3_lut.init = 16'hcaca;
    LUT4 mux_122_i9_3_lut (.A(n1467), .B(det_q4_28[9]), .C(n13818), .Z(n3444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i9_3_lut.init = 16'hcaca;
    LUT4 mux_122_i10_3_lut (.A(n1466), .B(det_q4_28[10]), .C(n13818), 
         .Z(n3443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i10_3_lut.init = 16'hcaca;
    LUT4 mux_122_i7_3_lut (.A(n1469), .B(det_q4_28[7]), .C(n13818), .Z(n3446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i7_3_lut.init = 16'hcaca;
    LUT4 mux_122_i8_3_lut (.A(n1468), .B(det_q4_28[8]), .C(n13818), .Z(n3445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i8_3_lut.init = 16'hcaca;
    LUT4 mux_122_i5_3_lut (.A(n1471), .B(det_q4_28[5]), .C(n13818), .Z(n3448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i5_3_lut.init = 16'hcaca;
    LUT4 mux_122_i6_3_lut (.A(n1470), .B(det_q4_28[6]), .C(n13818), .Z(n3447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i6_3_lut.init = 16'hcaca;
    LUT4 mux_122_i3_3_lut (.A(n1473), .B(det_q4_28[3]), .C(n13818), .Z(n3450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i3_3_lut.init = 16'hcaca;
    LUT4 mux_122_i4_3_lut (.A(n1472), .B(det_q4_28[4]), .C(n13818), .Z(n3449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i4_3_lut.init = 16'hcaca;
    LUT4 mux_122_i1_3_lut (.A(n1475), .B(det_q4_28[1]), .C(n13818), .Z(n3452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i1_3_lut.init = 16'hcaca;
    LUT4 mux_122_i2_3_lut (.A(n1474), .B(det_q4_28[2]), .C(n13818), .Z(n3451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_122_i2_3_lut.init = 16'hcaca;
    LUT4 mux_124_i31_3_lut (.A(n1445), .B(det_q4_28[31]), .C(n3454), .Z(n3487[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i31_3_lut.init = 16'hcaca;
    LUT4 i769_2_lut (.A(n1444), .B(n3454), .Z(n3487[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i769_2_lut.init = 16'h2222;
    LUT4 mux_124_i29_3_lut (.A(n1447), .B(det_q4_28[29]), .C(n3454), .Z(n3487[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i29_3_lut.init = 16'hcaca;
    LUT4 mux_124_i30_3_lut (.A(n1446), .B(det_q4_28[30]), .C(n3454), .Z(n3487[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i30_3_lut.init = 16'hcaca;
    LUT4 mux_124_i27_3_lut (.A(n1449), .B(det_q4_28[27]), .C(n3454), .Z(n3487[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i27_3_lut.init = 16'hcaca;
    LUT4 mux_124_i28_3_lut (.A(n1448), .B(det_q4_28[28]), .C(n3454), .Z(n3487[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i28_3_lut.init = 16'hcaca;
    LUT4 mux_124_i25_3_lut (.A(n1451), .B(det_q4_28[25]), .C(n3454), .Z(n3487[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i25_3_lut.init = 16'hcaca;
    LUT4 mux_124_i26_3_lut (.A(n1450), .B(det_q4_28[26]), .C(n3454), .Z(n3487[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i26_3_lut.init = 16'hcaca;
    LUT4 mux_124_i23_3_lut (.A(n1453), .B(det_q4_28[23]), .C(n3454), .Z(n3487[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i23_3_lut.init = 16'hcaca;
    LUT4 mux_124_i24_3_lut (.A(n1452), .B(det_q4_28[24]), .C(n3454), .Z(n3487[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i24_3_lut.init = 16'hcaca;
    LUT4 mux_124_i21_3_lut (.A(n1455), .B(det_q4_28[21]), .C(n3454), .Z(n3487[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i21_3_lut.init = 16'hcaca;
    LUT4 mux_124_i22_3_lut (.A(n1454), .B(det_q4_28[22]), .C(n3454), .Z(n3487[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i22_3_lut.init = 16'hcaca;
    LUT4 i1492_2_lut (.A(n3454), .B(inv_det_31__N_227), .Z(n62)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1492_2_lut.init = 16'h1111;
    LUT4 i1528_2_lut (.A(n2650), .B(inv_det_31__N_227), .Z(n50)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1528_2_lut.init = 16'h1111;
    LUT4 i1531_2_lut (.A(n2583), .B(inv_det_31__N_227), .Z(n49)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1531_2_lut.init = 16'h1111;
    LUT4 mux_124_i19_3_lut (.A(n1457), .B(det_q4_28[19]), .C(n3454), .Z(n3487[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i19_3_lut.init = 16'hcaca;
    LUT4 mux_124_i20_3_lut (.A(n1456), .B(det_q4_28[20]), .C(n3454), .Z(n3487[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i20_3_lut.init = 16'hcaca;
    LUT4 mux_124_i17_3_lut (.A(n1459), .B(det_q4_28[17]), .C(n3454), .Z(n3487[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i17_3_lut.init = 16'hcaca;
    LUT4 mux_124_i18_3_lut (.A(n1458), .B(det_q4_28[18]), .C(n3454), .Z(n3487[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i18_3_lut.init = 16'hcaca;
    LUT4 mux_124_i15_3_lut (.A(n1461), .B(det_q4_28[15]), .C(n3454), .Z(n3487[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i15_3_lut.init = 16'hcaca;
    LUT4 mux_124_i16_3_lut (.A(n1460), .B(det_q4_28[16]), .C(n3454), .Z(n3487[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i16_3_lut.init = 16'hcaca;
    LUT4 i1537_2_lut (.A(n2449), .B(inv_det_31__N_227), .Z(n47)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1537_2_lut.init = 16'h1111;
    LUT4 i1534_2_lut (.A(n2516), .B(inv_det_31__N_227), .Z(n48)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1534_2_lut.init = 16'h1111;
    LUT4 mux_124_i13_3_lut (.A(n1463), .B(det_q4_28[13]), .C(n3454), .Z(n3487[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i13_3_lut.init = 16'hcaca;
    LUT4 mux_124_i14_3_lut (.A(n1462), .B(det_q4_28[14]), .C(n3454), .Z(n3487[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i14_3_lut.init = 16'hcaca;
    LUT4 mux_124_i11_3_lut (.A(n1465), .B(det_q4_28[11]), .C(n3454), .Z(n3487[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i11_3_lut.init = 16'hcaca;
    LUT4 mux_124_i12_3_lut (.A(n1464), .B(det_q4_28[12]), .C(n3454), .Z(n3487[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i12_3_lut.init = 16'hcaca;
    LUT4 mux_124_i9_3_lut (.A(n1467), .B(det_q4_28[9]), .C(n3454), .Z(n3487[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i9_3_lut.init = 16'hcaca;
    LUT4 mux_124_i10_3_lut (.A(n1466), .B(det_q4_28[10]), .C(n3454), .Z(n3487[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i10_3_lut.init = 16'hcaca;
    LUT4 mux_124_i7_3_lut (.A(n1469), .B(det_q4_28[7]), .C(n3454), .Z(n3487[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i7_3_lut.init = 16'hcaca;
    LUT4 mux_124_i8_3_lut (.A(n1468), .B(det_q4_28[8]), .C(n3454), .Z(n3487[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i8_3_lut.init = 16'hcaca;
    LUT4 mux_124_i5_3_lut (.A(n1471), .B(det_q4_28[5]), .C(n3454), .Z(n3487[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i5_3_lut.init = 16'hcaca;
    LUT4 mux_124_i6_3_lut (.A(n1470), .B(det_q4_28[6]), .C(n3454), .Z(n3487[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i6_3_lut.init = 16'hcaca;
    LUT4 mux_124_i3_3_lut (.A(n1473), .B(det_q4_28[3]), .C(n3454), .Z(n3487[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i3_3_lut.init = 16'hcaca;
    LUT4 mux_124_i4_3_lut (.A(n1472), .B(det_q4_28[4]), .C(n3454), .Z(n3487[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i4_3_lut.init = 16'hcaca;
    LUT4 mux_124_i1_3_lut (.A(n1475), .B(det_q4_28[1]), .C(n3454), .Z(n3487[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i1_3_lut.init = 16'hcaca;
    CCU2C equal_1414_32 (.A0(det_q4_28[21]), .B0(det_q4_28[16]), .C0(det_q4_28[2]), 
          .D0(det_q4_28[28]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n13634), .S1(inv_det_31__N_227));
    defparam equal_1414_32.INIT0 = 16'h0001;
    defparam equal_1414_32.INIT1 = 16'h0000;
    defparam equal_1414_32.INJECT1_0 = "YES";
    defparam equal_1414_32.INJECT1_1 = "NO";
    CCU2C equal_1414_31 (.A0(det_q4_28[6]), .B0(det_q4_28[22]), .C0(det_q4_28[14]), 
          .D0(det_q4_28[30]), .A1(det_q4_28[4]), .B1(det_q4_28[24]), .C1(det_q4_28[12]), 
          .D1(det_q4_28[26]), .CIN(n13633), .COUT(n13634));
    defparam equal_1414_31.INIT0 = 16'h0001;
    defparam equal_1414_31.INIT1 = 16'h0001;
    defparam equal_1414_31.INJECT1_0 = "YES";
    defparam equal_1414_31.INJECT1_1 = "YES";
    LUT4 mux_124_i2_3_lut (.A(n1474), .B(det_q4_28[2]), .C(n3454), .Z(n3487[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_124_i2_3_lut.init = 16'hcaca;
    CCU2C equal_1414_29 (.A0(det_q4_28[1]), .B0(det_q4_28[9]), .C0(det_q4_28[11]), 
          .D0(det_q4_28[18]), .A1(det_q4_28[31]), .B1(det_q4_28[13]), 
          .C1(det_q4_28[23]), .D1(det_q4_28[20]), .CIN(n13632), .COUT(n13633));
    defparam equal_1414_29.INIT0 = 16'h0001;
    defparam equal_1414_29.INIT1 = 16'h0001;
    defparam equal_1414_29.INJECT1_0 = "YES";
    defparam equal_1414_29.INJECT1_1 = "YES";
    LUT4 mux_90_i1_3_lut (.A(n1475), .B(det_q4_28[1]), .C(n13829), .Z(n2380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_90_i1_3_lut.init = 16'hcaca;
    CCU2C equal_1414_27 (.A0(det_q4_28[29]), .B0(det_q4_28[19]), .C0(det_q4_28[17]), 
          .D0(det_q4_28[8]), .A1(det_q4_28[3]), .B1(det_q4_28[15]), .C1(det_q4_28[5]), 
          .D1(det_q4_28[7]), .CIN(n13631), .COUT(n13632));
    defparam equal_1414_27.INIT0 = 16'h0001;
    defparam equal_1414_27.INIT1 = 16'h0001;
    defparam equal_1414_27.INJECT1_0 = "YES";
    defparam equal_1414_27.INJECT1_1 = "YES";
    CCU2C equal_1414_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(det_q4_28[0]), .B1(det_q4_28[27]), .C1(det_q4_28[10]), .D1(det_q4_28[25]), 
          .COUT(n13631));   // c:/users/luso/documents/rtl_fpga/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam equal_1414_0.INIT0 = 16'h000F;
    defparam equal_1414_0.INIT1 = 16'h0001;
    defparam equal_1414_0.INJECT1_0 = "NO";
    defparam equal_1414_0.INJECT1_1 = "YES";
    
endmodule
