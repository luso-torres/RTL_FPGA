module handshaking(
input GO;
input Function;
input Data_Ready;
input clk;
output EnableA;
output EnableB;
output ResetB;
output Request_Data;
output add_sub);




endmodule