module converter_D(H,G,F,E,D);
input H,G,F,E;
output D;


assign D = H&G;


endmodule
