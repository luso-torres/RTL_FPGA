module meio_subtrator_flux(
input A, B
output D, Bout);




endmodule

