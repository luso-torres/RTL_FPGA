module decoder_4_16 (a_in,a_out);
input [3:0] a_in;
output reg [15:0] a_out;

always@(*) begin
	case (a_in)
		4'b0000: a_out = 16'b0000000000000001;
		4'b0001: a_out = 16'b0000000000000010;
		4'b0010: a_out = 16'b0000000000000100;
		4'b0011: a_out = 16'b0000000000001000;
		4'b0100: a_out = 16'b0000000000010000;
		4'b0101: a_out = 16'b0000000000100000;
		4'b0110: a_out = 16'b0000000001000000;
		4'b0111: a_out = 16'b0000000010000000;
		4'b1000: a_out = 16'b0000000100000000;
		4'b1001: a_out = 16'b0000001000000000;
		4'b1010: a_out = 16'b0000010000000000;
		4'b1011: a_out = 16'b0000100000000000;
		4'b1100: a_out = 16'b0001000000000000;
		4'b1101: a_out = 16'b0010000000000000;
		4'b1110: a_out = 16'b0100000000000000;
		4'b1111: a_out = 16'b1000000000000000;
		default: a_out = 16'b0000000000000000;
	endcase


end


endmodule