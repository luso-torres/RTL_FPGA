// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Thu Aug 14 21:58:43 2025
//
// Verilog Description of module matrix_inv
//

module matrix_inv (clk, reset, start, a, b, c, d, a_inv, b_inv, 
            c_inv, d_inv, error, ready) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(1[8:18])
    input clk;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(2[35:38])
    input reset;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(3[35:40])
    input start;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(4[35:40])
    input [15:0]a;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    input [15:0]b;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    input [15:0]c;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    input [15:0]d;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    output [15:0]a_inv;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    output [15:0]b_inv;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    output [15:0]c_inv;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    output [15:0]d_inv;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    output error;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(7[36:41])
    output ready;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(8[36:41])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(2[35:38])
    
    wire GND_net, VCC_net, reset_c, n6875, a_c_15, a_c_14, a_c_13, 
        a_c_12, a_c_11, a_c_10, a_c_9, a_c_8, a_c_7, a_c_6, a_c_5, 
        a_c_4, a_c_3, a_c_2, a_c_1, a_c_0, b_c_15, b_c_14, b_c_13, 
        b_c_12, b_c_11, b_c_10, b_c_9, b_c_8, b_c_7, b_c_6, b_c_5, 
        b_c_4, b_c_3, b_c_2, b_c_1, b_c_0, c_c_15, c_c_14, c_c_13, 
        c_c_12, c_c_11, c_c_10, c_c_9, c_c_8, c_c_7, c_c_6, c_c_5, 
        c_c_4, c_c_3, c_c_2, c_c_1, c_c_0, d_c_15, d_c_14, d_c_13, 
        d_c_12, d_c_11, d_c_10, d_c_9, d_c_8, d_c_7, d_c_6, d_c_5, 
        d_c_4, d_c_3, d_c_2, d_c_1, d_c_0, a_inv_c_15, a_inv_c_14, 
        a_inv_c_13, a_inv_c_12, a_inv_c_11, a_inv_c_10, a_inv_c_9, 
        a_inv_c_8, a_inv_c_7, a_inv_c_6, a_inv_c_5, a_inv_c_4, a_inv_c_3, 
        a_inv_c_2, a_inv_c_1, a_inv_c_0, b_inv_c_15, b_inv_c_14, b_inv_c_13, 
        b_inv_c_12, b_inv_c_11, b_inv_c_10, b_inv_c_9, b_inv_c_8, 
        b_inv_c_7, b_inv_c_6, b_inv_c_5, b_inv_c_4, b_inv_c_3, b_inv_c_2, 
        b_inv_c_1, b_inv_c_0, c_inv_c_15, c_inv_c_14, c_inv_c_13, 
        c_inv_c_12, c_inv_c_11, c_inv_c_10, c_inv_c_9, c_inv_c_8, 
        c_inv_c_7, c_inv_c_6, c_inv_c_5, c_inv_c_4, c_inv_c_3, c_inv_c_2, 
        c_inv_c_1, c_inv_c_0, d_inv_c_15, d_inv_c_14, d_inv_c_13, 
        d_inv_c_12, d_inv_c_11, d_inv_c_10, d_inv_c_9, d_inv_c_8, 
        d_inv_c_7, d_inv_c_6, d_inv_c_5, d_inv_c_4, d_inv_c_3, d_inv_c_2, 
        d_inv_c_1, d_inv_c_0, n6874, n6873, n6872, n6871, n6870, 
        n6869, n179, n178;
    wire [31:0]det_q4_28;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(24[34:43])
    wire [15:0]a_reg;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(25[34:39])
    wire [15:0]b_reg;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(25[41:46])
    wire [15:0]c_reg;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(25[48:53])
    wire [15:0]d_reg;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(25[55:60])
    
    wire n6868, det_zero_reg, n7184, n7439, n6867, n6373, n6866, 
        n7185, n6865, n7186, n7187, n7188, n7189, n7190, n6864, 
        n6863, n6862, n6861, n6860, n6859, n6858, n6857, n6856, 
        n6855, n6854, n6447, n6446, n6445, n6444, n6443, n6442, 
        n6441, n6440, n6853, n6439, n6852, n6438, n6851, n6437, 
        n6850, n6436, n6435, n6434, n6433, n6432, n6431, n6430, 
        n6429, n6428, n6427, n6426, n6425, n6424, n6423, n6422, 
        n6421, n6420, n6419, n6849, n6848, n6847, n6418, n6846, 
        n6845, n6844, n6417, n6843, n6842, n6841, n6840, n6839, 
        n6838, n6837, n6836, n6835, n6941, n6940, n6939, n6938, 
        n6937, n6936, n6935, n6934, n6933, n6932, n6931, n6930, 
        n6929, n6928, n6927, n6926, n6925, n6924, n6923, n6922, 
        n6921, n53_adj_1114, n60_adj_1115, n6920, n6919, n6918, 
        n6917, n6916, n6915, n6914, n6913, n6912, n6911, n6910, 
        n6909, n6834, n6833, n7223, n7224, n7225, n7226;
    wire [47:0]prod_a;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(34[34:40])
    
    wire n173, n172, n171, n170, n169, n168, n167, n166, n165, 
        n164, n163, n162, n161, n160, n159;
    wire [47:0]prod_b;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(34[42:48])
    
    wire n158, n157, n156, n155, n154, n153, n152, n151, n150, 
        n149, n148, n147, n6832, n6831, n6830;
    wire [47:0]prod_c;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(34[50:56])
    
    wire n6829, n6828, n6827, n6826, n6825, n6824, n6823, n6822, 
        n6821, n6820, n6819, n6818, n6817, n7352, n7415;
    wire [47:0]prod_d;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(34[58:64])
    
    wire n7353, n7414, n7354, n7413, n7355, n7412, n7356, n7411, 
        n7357, n7410, n7358, n7409, n7359, n7408, n7360, n6816, 
        n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
        n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
        n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, 
        n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
        n98, n99, n100, n101;
    wire [31:0]det_q4_28_31__N_551;
    
    wire det_zero_reg_N_907, det_zero_reg_N_905, n6815, n6814, n6813, 
        n6812, n6811, n6810, n6809, n6808, n6807, n6806, n7851, 
        n6805, n6804, n6803, n6802, n6801, n6800, n6799, n6798, 
        n6797, n6796, n6795, n6794, n6793, n6792, n6791, n6790, 
        n6789, n6788, n6787, n6786, n6785, n7419, n6784, n6783, 
        n6782, n6781, n6780, n6779, n6778, n6777, n6776, n6775, 
        n6774, n6773, n6772, n6771, n6770, n6769, n6768, n6767, 
        n6766, n6765, n6764, n6763, n6762, n6761, n6760, n179_adj_1116, 
        n178_adj_1117, n177, n176, n175, n174, n173_adj_1118, n172_adj_1119, 
        n171_adj_1120, n7462, n7440, n6372, n7461, n7441, n6371, 
        n170_adj_1121, n169_adj_1122, n7227, n168_adj_1123, n167_adj_1124, 
        n166_adj_1125, n7228, n165_adj_1126, n164_adj_1127, n163_adj_1128, 
        n162_adj_1129, n161_adj_1130, n160_adj_1131, n159_adj_1132, 
        n158_adj_1133, n157_adj_1134, n156_adj_1135, n155_adj_1136, 
        n154_adj_1137, n153_adj_1138, n152_adj_1139, n151_adj_1140, 
        n150_adj_1141, n149_adj_1142, n148_adj_1143, n147_adj_1144, 
        n6759, n6758, n6757, n6756, n6755, n6754, n6753, n6752, 
        n6751, n6750, n6749, n6748, n6747, n6746, n6745, n6744, 
        n7255, n7229, n7318, n7256, n7317, n7230, n7257, n7316, 
        n7258, n7231, n7315, n7259, n7314, n7232, n7260, n7313, 
        n7261, n7312, n7262, n7311, n7263, n7310, n7264, n7309, 
        n7265, n7308, n7266, n7307, n7267, n7306, n7268, n7305, 
        n7269, n7304, n7270, n7303, n7271, n7302, n7272, n7301, 
        n7273, n7300, n7274, n7299, n7275, n7298, n7276, n7297, 
        n7277, n7296, n7233, n7278, n7295, n7279, n7234, n7294, 
        n7280, n6743, n7235, n6742, n7293, n6741, n7236, n7281, 
        n7292, n7282, n7291, n7283, n7290, n7284, n7289, n7285, 
        n7288, n7286, n7287, n7191, n7192, n7193, n7194, n7195, 
        n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
        n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, 
        n6740, n7212, n6739, n7237, n6738, n7213, n6737, n7238, 
        n6736, n7214, n6735, n7239, n6734, n7215, n6733;
    wire [47:0]a_inv_15__N_487;
    wire [47:0]b_inv_15__N_503;
    wire [47:0]c_inv_15__N_519;
    wire [47:0]d_inv_15__N_535;
    
    wire n7407, n7361, n7406, n7362, n7405, n7363, n7404, n7364, 
        n7403, n7365, n7402, n7366, n7401, n7367, n7400, n7368, 
        n7399, n7369, n7398, n7370, n7397, n7371, n7396, n7372, 
        n7395, n7373, n7394, n7374, n7393, n7375, n7392, n7376, 
        n7391, n7377, n7390, n7378, n7389, n7379, n7388, n7380, 
        n7387, n7381, n7386, n7382, n7385, n7383, n7384, n7159, 
        n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, 
        n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, 
        n177_adj_1145, n176_adj_1146, n175_adj_1147, n174_adj_1148, 
        n173_adj_1149, n172_adj_1150, n171_adj_1151, n170_adj_1152, 
        n169_adj_1153, n168_adj_1154, n167_adj_1155, n166_adj_1156, 
        n165_adj_1157, n164_adj_1158, n163_adj_1159, n162_adj_1160, 
        n161_adj_1161, n160_adj_1162, n159_adj_1163, n158_adj_1164, 
        n157_adj_1165, n156_adj_1166, n155_adj_1167, n154_adj_1168, 
        n153_adj_1169, n152_adj_1170, n151_adj_1171, n150_adj_1172, 
        n149_adj_1173, n148_adj_1174, n147_adj_1175, n6732, n6731, 
        n6730, n6729, n6728, n6727, n6726, n6725, n6724, n6723, 
        n6722, n6721, n6720, n6719, n6718, n6717, n130, n7549, 
        n128, n7548, n126, n7547, n124, n7546, n122, n7545, 
        n120, n7544, n118, n7543, n116, n7542, n114, n7541, 
        n112, n7540, n110, n7539, n108, n7538, n106, n7537, 
        n104, n7536, n102, n7535, n7500, n7534, n7501, n7533, 
        n7502, n7532, n7503, n7531, n7504, n7530, n7505, n7529, 
        n7506, n7528, n7507, n7527, n7508, n7526, n7509, n7525, 
        n7510, n7524, n7511, n7523, n7512, n7522, n7513, n7521, 
        n7514, n7520, n7515, n7519, n68_adj_1176, n7518, n7127, 
        n7499, n7128, n7498, n7129, n7497, n7130, n7496, n7131, 
        n7495, n7132, n7494, n7133, n7493, n7134, n7492, n7135, 
        n7491, n7136, n7490, n7137, n7489, n7138, n7488, n7139, 
        n7487, n7140, n7486, n7141, n7485, n7142, n7484, n7143, 
        n7483, n7144, n7482, n7145, n7481, n7146, n7480, n7147, 
        n7479, n7148, n7478, n7149, n7477, n7150, n7476, n7151, 
        n7475, n7152, n7474, n7153, n7473, n7154, n7472, n7155, 
        n7471, n7156, n7470, n7157, n7469, n7158, n7468, n6716, 
        n6699, n6698, n6697, n6696, n6695, n6694, n6693, n6692, 
        n6691, n6690, n6689, n6688, n6687, n6974, n6973, n6972, 
        n6971, n6970, n6969, n6968, n6967, n6966, n6965, n6964, 
        n6963, n6962, n6961, n6960, n6959, n6958, n6957, n6956, 
        n6955, n6954, n6953, n6952, n6951, n6950, n6949, n6948, 
        n6947, n6946, n6945, n6944, n6943, n6942, n7216, n7217, 
        n7218, n6416, n7219, n7220, n7221, n7222, n6686, n6685, 
        n6684, n6683, n6682, n6681, n6680, n6679, n6678, n6677, 
        n6676, n6675, n6674, n6673, n6672, n6671, n6670, n7853, 
        n4610, n4609, n4608, n4607, n4606, n4605, n4604, n4603, 
        n4602, n4601, n4600, n4599, n4598, n4597, n4596, n4595, 
        n4594, n4593, n4592, n4591, n4590, n7855, n7857, n7859, 
        n7861, n7863, n7865, n7895, n7897, n7899, n7901, n7903, 
        n7905, n7907, n7909, n7911, n7893, n7891, n7889, n7887, 
        n7885, n7883, n7881, n7879, n7877, n7875, n7873, n52_adj_1177, 
        n7871, n7869, n7867, n7240, n6669, n7460, n7176, n7177, 
        n7178, n7179, n7180, n7181, n7182, n7183, n6668, n6667, 
        n6666, n6665, n6664, n6663, n6662, n6661, n6660, n6659, 
        n6658, n6657, n6656, n6655, n6654, n6653, n6652, n6651, 
        n6650, n6649, n6648, n6647, n6646, n6908, n7442, n6907, 
        n6906, n6905, n6904, n6903, n6902, n6901, n6900, n6899, 
        n6898, n6897, n6896, n6895, n6894, n6893, n6892, n6891, 
        n6890, n6889, n6888, n6887, n6886, n6885, n6884, n6883, 
        n6882, n6881, n6880, n6879, n6878, n6877, n6876, n6645, 
        n6644, n6643, n6642, n6641, n6640, n6639, n6638, n6637, 
        n6636, n6635, n6634, n6633, n6632, n6631, n6630, n6629, 
        n6628, n6627, n6626, n6625, n6624, n6623, n6622, n6621, 
        n6620, n6619, n6618, n6617, n6616, n6615, n6614, n6613, 
        n6612, n6611, n6610, n6609, n6608, n6607, n6606, n6605, 
        n6604, n6603, n6602, n6601, n6600, n6599, n179_adj_1178, 
        n178_adj_1179, n177_adj_1180, n176_adj_1181, n175_adj_1182, 
        n174_adj_1183, n173_adj_1184, n172_adj_1185, n171_adj_1186, 
        n170_adj_1187, n169_adj_1188, n168_adj_1189, n167_adj_1190, 
        n166_adj_1191, n165_adj_1192, n164_adj_1193, n163_adj_1194, 
        n162_adj_1195, n161_adj_1196, n160_adj_1197, n159_adj_1198, 
        n158_adj_1199, n157_adj_1200, n7350, n7349, n7348, n7347, 
        n7346, n7345, n7344, n7343, n7342, n7341, n7340, n7339, 
        n7338, n7337, n7336, n7335, n7334, n7333, n7332, n7331, 
        n7330, n7329, n7328, n7327, n7326, n7325, n7324, n7323, 
        n7322, n7321, n7320, n7319, n156_adj_1201, n155_adj_1202, 
        n154_adj_1203, n153_adj_1204, n152_adj_1205, n151_adj_1206, 
        n150_adj_1207, n149_adj_1208, n148_adj_1209, n147_adj_1210, 
        n6598, n6597, n6596, n6595, n6594, n6593, n6592, n6591, 
        n6370, n7459, n7443, n6369, n7458, n7444, n6368, n7457, 
        n7445, n6367, n7456, n7446, n6366, n7455, n7447, n6365, 
        n7454, n7448, n6364, n7453, n7449, n6363, n7452, n7450, 
        n6362, n7451, n6590, n6589, n6588, n7241, n6587, n7242, 
        n6586, n7243, n6585, n7244, n6584, n7245, n6583, n7246, 
        n6582, n7247, n6581, n7248, n6580, n7249, n130_adj_1211, 
        n7250, n7126, n7251, n128_adj_1212, n7252, n7125, n7253, 
        n126_adj_1213, n7254, n7124, n124_adj_1214, n7123, n122_adj_1215, 
        n7122, n120_adj_1216, n7121, n118_adj_1217, n7120, n116_adj_1218, 
        n7119, n114_adj_1219, n7118, n112_adj_1220, n7117, n110_adj_1221, 
        n7116, n108_adj_1222, n7115, n106_adj_1223, n7114, n104_adj_1224, 
        n7113, n102_adj_1225, n7112, n7111, n7110, n7109, n7108, 
        n7107, n5373, n5308, n5307, n5306, n5305, n5304, n5303, 
        n5302, n5301, n5300, n5299, n5298, n5297, n5296, n5295, 
        n5294, n5293, n7106, n7105, n7104, n7103, n7102, n7101, 
        n7100, n7099, n7098, n7097, n7096, n68_adj_1226, n7095, 
        n7059, n7058, n7057, n7056, n7055, n7054, n7053, n7052, 
        n7051, n7050, n7417, n7049, n6579, n7048, n7047, n7046, 
        n6578, n7045, n6577, n7044, n7043, n7042, n7041, n7040, 
        n7039, n7038, n7037, n7036, n7035, n5277, n5212, n5211, 
        n5210, n5209, n5208, n5207, n5206, n5205, n5204, n5203, 
        n5202, n5201, n5200, n5199, n5198, n5197, n7008, n7034, 
        n7033, n7032, n7418, n7031, n7030, n7029, n6576, n7028, 
        n6575, n7027, n6574, n6573, next_state_2__N_68_c_0;
    wire [2:0]next_state_2__N_65;
    
    wire n6572, n6571, n6570, n6569, n6568, n6567, n6566, n6565, 
        n6564, n6563, n6562, n6561, n6560, n6559, n6558, n6557, 
        n179_adj_1227, n178_adj_1228, n50_adj_1229, n6556, n4589, 
        n6555, n4588, n6554, n6553, n6552, n49_adj_1230, n6551, 
        n6550;
    wire [2:0]proximo_estado_2__N_952;
    
    wire n4646, n4587, n4586, n4585, n7916, n6549, n7026;
    wire [32:0]regA;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(27[8:12])
    
    wire n4584, clk_c_enable_410, clk_c_enable_395, n4583, n6548, 
        n48_adj_1231, n177_adj_1232, n176_adj_1233, n175_adj_1234, n174_adj_1235, 
        n6547, n7025, n7024, n7023, n6546, n7022, n7021, n7020, 
        n6545, n7019, n7913, n6544, n7018, n6543, n7017, n6542, 
        n7016, n6541, n7015, n6540, n7014, n6539, n7013, n6538, 
        n7012, n6537, n7011, n6536, n7010, n6535, n7009, n6534, 
        n6533, n6532, n7517, n6531, n7516, n6530, n6529, n6361, 
        n6528, n7467, n6527, n6526;
    wire [31:0]quotient_31__N_908;
    
    wire n6360, n6525, n7466, n6524, n7436, n6523, n6359, n6522, 
        n7465, n6521, n7437, n6520, n6358, n6519, n7464, n6518, 
        n7438, n6517, n6516, n6515, n6514, n6513, n6512, n6511, 
        n6510, n6509, n6508, n6507, n6506, n2820, n6357, n6505, 
        n4582, n2813, clk_c_enable_431, clk_c_enable_145, n2810, n2809, 
        n6504, n2808, clk_c_enable_363, n6503, n6502, n58_adj_1236, 
        n7463, n6501, n6500, n3859, n3860, n3861, n3863, clk_c_enable_239, 
        n4581, n6499, n44_adj_1237, n43_adj_1238, n6498, n6497, 
        n6496, n37_adj_1239, n4580, clk_c_enable_432, n6495, n6494, 
        n6493, n6492, n6491, n6490, n6489, n6488, n6487, n6486, 
        n6485, n6484, n6483, n6482, n6481, n6480, n6479, n6478, 
        n6477, n6476, n4579, n8033, n8032, n4578, n6475, n6474, 
        n6473, n6472, n6471, n6470, n6469, n6468, n6467, n6466, 
        n6465, n6464, n6463, n6462, n6461, n6460, n6459, n6458, 
        n6457, n6456, n6455, n6454, n6453, n6975, n6976, n6977, 
        n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
        n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
        n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
        n7002, n7003, n7004, n7005, n7006, n7007, n6452, n6451, 
        n6450, n6449, n6448, n6415, n6414, n6413, n6412, n6411, 
        n6410, n6409, n6408, n6407, n6406, n6405, n6404, n6403, 
        n6402, n6401, n6400, n6399, n6398, n6397, n6396, n6395, 
        n6394, n6393, n6392, n6391, n7550, n6390, n7551, n7094, 
        n7552, n6389, n7553, n6388, n7554, n6387, n7555, n6386, 
        n7556, n6385, n7557, n6384, n7558, n6383, n7559, n6382, 
        n7560, n6381, n7561, n6380, n7562, n6379, n7563, n6378, 
        n7564, n6377, n7565, n6376, n7566, n6375, n7584, n6356, 
        n7583, n7585, n7582, n7586, n7581, n7587, n7580, n7588, 
        n7579, n7589, n7578, n7590, n7577, n7591, n7576, n7592, 
        n7575, n7593, n7574, n7594, n7573, n7595, n7572, n7596, 
        n7571, n7597, n7570, n7598, n7569, n7599, n7568, n7600, 
        n7567, n7601, n7093, n6374, n7076, n7077, n7078, n7079, 
        n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, 
        n7088, n7089, n7090, n7091, n7092, n7351, n7416, n7602, 
        n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, 
        n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, 
        n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, 
        n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, 
        n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, 
        n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, 
        n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, 
        n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, 
        n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, 
        n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, 
        n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, 
        n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, 
        n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, 
        n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, 
        n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, 
        n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, 
        n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, 
        n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, 
        n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, 
        n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, 
        n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, 
        n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, 
        n7779, n7849, n8266, n8265, n8264, n8263, n38_adj_1240, 
        n41_adj_1241, n44_adj_1242, n47_adj_1243, n50_adj_1244, n53_adj_1245, 
        n56_adj_1246, n59_adj_1247, n62_adj_1248, n65_adj_1249, n68_adj_1250, 
        n71_adj_1251, n74_adj_1252, n77_adj_1253, n80_adj_1254, n83_adj_1255, 
        n86_adj_1256, n8262, n8040, clk_c_enable_348, clk_c_enable_411, 
        n8817, n38_adj_1257, n41_adj_1258, n44_adj_1259, n47_adj_1260, 
        n50_adj_1261, n53_adj_1262, n56_adj_1263, n59_adj_1264, n62_adj_1265, 
        n65_adj_1266, n68_adj_1267, n71_adj_1268, n74_adj_1269, n77_adj_1270, 
        n80_adj_1271, n83_adj_1272, n86_adj_1273, n8725, n8724, n8381, 
        n8380, n8379, n8378, n8377, n8376, n8375, n8374, n8373, 
        n8372, n8371, n8370, n8369, n8368, n8367, n8366, n8365, 
        n8360, n8359, n8358, n8357, n8356, n8355, n8354, n8353, 
        n8352, n8351, n8350, n8349, n8348, n8347, n8346, n8344, 
        n8343, n8342, n8341, n8340, n8339, n8338, n8337, n8336, 
        n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328, 
        n8327, n8326, n8325, n8324, n8323, n8322, n8321, n8320, 
        n8319, n8318, n8317, n8316, n8315, n8314, n8312, n8311, 
        n8310, n8309, n8308, n8307, n8306, n72_adj_1274, n8305, 
        n75_adj_1275, n8304, n78_adj_1276, n8303, n81_adj_1277, n8302, 
        n84_adj_1278, n8301, n87_adj_1279, n8300, n90_adj_1280, n8299, 
        n93_adj_1281, n8298, n96_adj_1282, n99_adj_1283, n102_adj_1284, 
        n105, n108_adj_1285, n8293, n111, n8292, n114_adj_1286, 
        n8291, n117, n8290, n120_adj_1287, n8289, n123, n8288, 
        n126_adj_1288, n8287, n129, n8286, n132, n135, n8284, 
        n138, n8283, n141, n8282, n144, n8281, n147_adj_1289, 
        n8280, n150_adj_1290, n8279, n153_adj_1291, n8278, n156_adj_1292, 
        n8277, n159_adj_1293, n162_adj_1294, n8275, n165_adj_1295, 
        n8274, n168_adj_1296, n8273, n8272, n8267, n8268, n8269, 
        n55_adj_1297, n8270, n8271, n62_adj_1298, n8261;
    
    VHI i2 (.Z(VCC_net));
    LUT4 i30_4_lut (.A(n53_adj_1114), .B(n60_adj_1115), .C(n43_adj_1238), 
         .D(n44_adj_1237), .Z(n62_adj_1298)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i30_4_lut.init = 16'hfffe;
    OB a_inv_pad_15 (.I(a_inv_c_15), .O(a_inv[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    FD1P3AX b_reg_i0_i0 (.D(b_c_0), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i0.GSR = "ENABLED";
    ALU54B lat_alu_9 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n6913), .SIGNEDIB(n6986), .SIGNEDCIN(n7059), .A35(n6912), 
           .A34(n6911), .A33(n6910), .A32(n6909), .A31(n6908), .A30(n6907), 
           .A29(n6906), .A28(n6905), .A27(n6904), .A26(n6903), .A25(n6902), 
           .A24(n6901), .A23(n6900), .A22(n6899), .A21(n6898), .A20(n6897), 
           .A19(n6896), .A18(n6895), .A17(n6894), .A16(n6893), .A15(n6892), 
           .A14(n6891), .A13(n6890), .A12(n6889), .A11(n6888), .A10(n6887), 
           .A9(n6886), .A8(n6885), .A7(n6884), .A6(n6883), .A5(n6882), 
           .A4(n6881), .A3(n6880), .A2(n6879), .A1(n6878), .A0(n6877), 
           .B35(n6985), .B34(n6984), .B33(n6983), .B32(n6982), .B31(n6981), 
           .B30(n6980), .B29(n6979), .B28(n6978), .B27(n6977), .B26(n6976), 
           .B25(n6975), .B24(n6974), .B23(n6973), .B22(n6972), .B21(n6971), 
           .B20(n6970), .B19(n6969), .B18(n6968), .B17(n6967), .B16(n6966), 
           .B15(n6965), .B14(n6964), .B13(n6963), .B12(n6962), .B11(n6961), 
           .B10(n6960), .B9(n6959), .B8(n6958), .B7(n6957), .B6(n6956), 
           .B5(n6955), .B4(n6954), .B3(n6953), .B2(n6952), .B1(n6951), 
           .B0(n6950), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n6949), .MA34(n6948), .MA33(n6947), .MA32(n6946), .MA31(n6945), 
           .MA30(n6944), .MA29(n6943), .MA28(n6942), .MA27(n6941), .MA26(n6940), 
           .MA25(n6939), .MA24(n6938), .MA23(n6937), .MA22(n6936), .MA21(n6935), 
           .MA20(n6934), .MA19(n6933), .MA18(n6932), .MA17(n6931), .MA16(n6930), 
           .MA15(n6929), .MA14(n6928), .MA13(n6927), .MA12(n6926), .MA11(n6925), 
           .MA10(n6924), .MA9(n6923), .MA8(n6922), .MA7(n6921), .MA6(n6920), 
           .MA5(n6919), .MA4(n6918), .MA3(n6917), .MA2(n6916), .MA1(n6915), 
           .MA0(n6914), .MB35(n7022), .MB34(n7021), .MB33(n7020), .MB32(n7019), 
           .MB31(n7018), .MB30(n7017), .MB29(n7016), .MB28(n7015), .MB27(n7014), 
           .MB26(n7013), .MB25(n7012), .MB24(n7011), .MB23(n7010), .MB22(n7009), 
           .MB21(n7008), .MB20(n7007), .MB19(n7006), .MB18(n7005), .MB17(n7004), 
           .MB16(n7003), .MB15(n7002), .MB14(n7001), .MB13(n7000), .MB12(n6999), 
           .MB11(n6998), .MB10(n6997), .MB9(n6996), .MB8(n6995), .MB7(n6994), 
           .MB6(n6993), .MB5(n6992), .MB4(n6991), .MB3(n6990), .MB2(n6989), 
           .MB1(n6988), .MB0(n6987), .CIN53(n7058), .CIN52(n7057), .CIN51(n7056), 
           .CIN50(n7055), .CIN49(n7054), .CIN48(n7053), .CIN47(n7052), 
           .CIN46(n7051), .CIN45(n7050), .CIN44(n7049), .CIN43(n7048), 
           .CIN42(n7047), .CIN41(n7046), .CIN40(n7045), .CIN39(n7044), 
           .CIN38(n7043), .CIN37(n7042), .CIN36(n7041), .CIN35(n7040), 
           .CIN34(n7039), .CIN33(n7038), .CIN32(n7037), .CIN31(n7036), 
           .CIN30(n7035), .CIN29(n7034), .CIN28(n7033), .CIN27(n7032), 
           .CIN26(n7031), .CIN25(n7030), .CIN24(n7029), .CIN23(n7028), 
           .CIN22(n7027), .CIN21(n7026), .CIN20(n7025), .CIN19(n7024), 
           .CIN18(n7023), .CIN17(n177), .CIN16(n178_adj_1117), .CIN15(n179_adj_1116), 
           .CIN14(n6716), .CIN13(n6717), .CIN12(n6718), .CIN11(n6719), 
           .CIN10(n6720), .CIN9(n6721), .CIN8(n6722), .CIN7(n6723), 
           .CIN6(n6724), .CIN5(n6725), .CIN4(n6726), .CIN3(n6727), .CIN2(n6728), 
           .CIN1(n6729), .CIN0(n6730), .OP10(GND_net), .OP9(VCC_net), 
           .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), 
           .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), 
           .OP0(VCC_net), .R29(n147_adj_1144), .R28(n148_adj_1143), .R27(n149_adj_1142), 
           .R26(n150_adj_1141), .R25(n151_adj_1140), .R24(n152_adj_1139), 
           .R23(n153_adj_1138), .R22(n154_adj_1137), .R21(n155_adj_1136), 
           .R20(n156_adj_1135), .R19(n157_adj_1134), .R18(n158_adj_1133), 
           .R17(n159_adj_1132), .R16(n160_adj_1131), .R15(n161_adj_1130), 
           .R14(n162_adj_1129), .R13(n163_adj_1128), .R12(n164_adj_1127), 
           .R11(n165_adj_1126), .R10(n166_adj_1125), .R9(n167_adj_1124), 
           .R8(n168_adj_1123), .R7(n169_adj_1122), .R6(n170_adj_1121), 
           .R5(n171_adj_1120), .R4(n172_adj_1119), .R3(n173_adj_1118), 
           .R2(n174), .R1(n175), .R0(n176));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam lat_alu_9.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_9.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_9.REG_FLAG_CLK = "NONE";
    defparam lat_alu_9.REG_FLAG_CE = "CE0";
    defparam lat_alu_9.REG_FLAG_RST = "RST0";
    defparam lat_alu_9.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASK01 = "0x00000000000000";
    defparam lat_alu_9.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_9.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_9.CLK0_DIV = "ENABLED";
    defparam lat_alu_9.CLK1_DIV = "ENABLED";
    defparam lat_alu_9.CLK2_DIV = "ENABLED";
    defparam lat_alu_9.CLK3_DIV = "ENABLED";
    defparam lat_alu_9.MCPAT = "0x00000000000000";
    defparam lat_alu_9.MASKPAT = "0x00000000000000";
    defparam lat_alu_9.RNDPAT = "0x00000000000000";
    defparam lat_alu_9.GSR = "DISABLED";
    defparam lat_alu_9.RESETMODE = "SYNC";
    defparam lat_alu_9.MULT9_MODE = "DISABLED";
    defparam lat_alu_9.LEGACY = "DISABLED";
    MULT18X18D lat_mult_10 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(GND_net), .B16(n5293), .B15(n5294), 
            .B14(n5295), .B13(n5296), .B12(n5297), .B11(n5298), .B10(n5299), 
            .B9(n5300), .B8(n5301), .B7(n5302), .B6(n5303), .B5(n5304), 
            .B4(n5305), .B3(n5306), .B2(n5307), .B1(n5308), .B0(n5373), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n7181), .ROA16(n7180), 
            .ROA15(n7179), .ROA14(n7178), .ROA13(n7177), .ROA12(n7176), 
            .ROA11(n7175), .ROA10(n7174), .ROA9(n7173), .ROA8(n7172), 
            .ROA7(n7171), .ROA6(n7170), .ROA5(n7169), .ROA4(n7168), 
            .ROA3(n7167), .ROA2(n7166), .ROA1(n7165), .ROA0(n7164), 
            .ROB17(n7199), .ROB16(n7198), .ROB15(n7197), .ROB14(n7196), 
            .ROB13(n7195), .ROB12(n7194), .ROB11(n7193), .ROB10(n7192), 
            .ROB9(n7191), .ROB8(n7190), .ROB7(n7189), .ROB6(n7188), 
            .ROB5(n7187), .ROB4(n7186), .ROB3(n7185), .ROB2(n7184), 
            .ROB1(n7183), .ROB0(n7182), .P35(n7236), .P34(n7235), .P33(n7234), 
            .P32(n7233), .P31(n7232), .P30(n7231), .P29(n7230), .P28(n7229), 
            .P27(n7228), .P26(n7227), .P25(n7226), .P24(n7225), .P23(n7224), 
            .P22(n7223), .P21(n7222), .P20(n7221), .P19(n7220), .P18(n7219), 
            .P17(n7218), .P16(n7217), .P15(n7216), .P14(n7215), .P13(n7214), 
            .P12(n7213), .P11(n7212), .P10(n7211), .P9(n7210), .P8(n7209), 
            .P7(n7208), .P6(n7207), .P5(n7206), .P4(n7205), .P3(n7204), 
            .P2(n7203), .P1(n7202), .P0(n7201), .SIGNEDP(n7200));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam lat_mult_10.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_10.REG_INPUTA_CE = "CE3";
    defparam lat_mult_10.REG_INPUTA_RST = "RST3";
    defparam lat_mult_10.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTB_CE = "CE0";
    defparam lat_mult_10.REG_INPUTB_RST = "RST0";
    defparam lat_mult_10.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTC_CE = "CE0";
    defparam lat_mult_10.REG_INPUTC_RST = "RST0";
    defparam lat_mult_10.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_10.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_10.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_10.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_10.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_10.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_10.CLK0_DIV = "ENABLED";
    defparam lat_mult_10.CLK1_DIV = "ENABLED";
    defparam lat_mult_10.CLK2_DIV = "ENABLED";
    defparam lat_mult_10.CLK3_DIV = "ENABLED";
    defparam lat_mult_10.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_10.GSR = "DISABLED";
    defparam lat_mult_10.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_10.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_10.MULT_BYPASS = "DISABLED";
    defparam lat_mult_10.RESETMODE = "ASYNC";
    LUT4 i26_4_lut (.A(n37_adj_1239), .B(n52_adj_1177), .C(det_q4_28_31__N_551[3]), 
         .D(det_q4_28_31__N_551[31]), .Z(n58_adj_1236)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i26_4_lut.init = 16'hfffe;
    FD1P3AX c_reg_i0_i0 (.D(c_c_0), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i0.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i0 (.D(d_c_0), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i0.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i0 (.D(det_q4_28_31__N_551[0]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i0.GSR = "ENABLED";
    FD1P3AX prod_d__3_res11_e2__i1 (.D(a_reg[0]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n130));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i1.GSR = "DISABLED";
    MULT18X18D lat_mult_7 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(GND_net), .B16(GND_net), 
            .B15(GND_net), .B14(GND_net), .B13(GND_net), .B12(GND_net), 
            .B11(GND_net), .B10(GND_net), .B9(GND_net), .B8(GND_net), 
            .B7(GND_net), .B6(GND_net), .B5(GND_net), .B4(GND_net), 
            .B3(GND_net), .B2(GND_net), .B1(GND_net), .B0(GND_net), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n6967), .ROA16(n6966), 
            .ROA15(n6965), .ROA14(n6964), .ROA13(n6963), .ROA12(n6962), 
            .ROA11(n6961), .ROA10(n6960), .ROA9(n6959), .ROA8(n6958), 
            .ROA7(n6957), .ROA6(n6956), .ROA5(n6955), .ROA4(n6954), 
            .ROA3(n6953), .ROA2(n6952), .ROA1(n6951), .ROA0(n6950), 
            .ROB17(n6985), .ROB16(n6984), .ROB15(n6983), .ROB14(n6982), 
            .ROB13(n6981), .ROB12(n6980), .ROB11(n6979), .ROB10(n6978), 
            .ROB9(n6977), .ROB8(n6976), .ROB7(n6975), .ROB6(n6974), 
            .ROB5(n6973), .ROB4(n6972), .ROB3(n6971), .ROB2(n6970), 
            .ROB1(n6969), .ROB0(n6968), .P35(n7022), .P34(n7021), .P33(n7020), 
            .P32(n7019), .P31(n7018), .P30(n7017), .P29(n7016), .P28(n7015), 
            .P27(n7014), .P26(n7013), .P25(n7012), .P24(n7011), .P23(n7010), 
            .P22(n7009), .P21(n7008), .P20(n7007), .P19(n7006), .P18(n7005), 
            .P17(n7004), .P16(n7003), .P15(n7002), .P14(n7001), .P13(n7000), 
            .P12(n6999), .P11(n6998), .P10(n6997), .P9(n6996), .P8(n6995), 
            .P7(n6994), .P6(n6993), .P5(n6992), .P4(n6991), .P3(n6990), 
            .P2(n6989), .P1(n6988), .P0(n6987), .SIGNEDP(n6986));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam lat_mult_7.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_7.REG_INPUTA_CE = "CE3";
    defparam lat_mult_7.REG_INPUTA_RST = "RST3";
    defparam lat_mult_7.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTB_CE = "CE0";
    defparam lat_mult_7.REG_INPUTB_RST = "RST0";
    defparam lat_mult_7.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTC_CE = "CE0";
    defparam lat_mult_7.REG_INPUTC_RST = "RST0";
    defparam lat_mult_7.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_7.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_7.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_7.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_7.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_7.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_7.CLK0_DIV = "ENABLED";
    defparam lat_mult_7.CLK1_DIV = "ENABLED";
    defparam lat_mult_7.CLK2_DIV = "ENABLED";
    defparam lat_mult_7.CLK3_DIV = "ENABLED";
    defparam lat_mult_7.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_7.GSR = "DISABLED";
    defparam lat_mult_7.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_7.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_7.MULT_BYPASS = "DISABLED";
    defparam lat_mult_7.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_6 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(GND_net), .B16(GND_net), 
            .B15(GND_net), .B14(GND_net), .B13(GND_net), .B12(GND_net), 
            .B11(GND_net), .B10(GND_net), .B9(GND_net), .B8(GND_net), 
            .B7(GND_net), .B6(GND_net), .B5(GND_net), .B4(GND_net), 
            .B3(GND_net), .B2(GND_net), .B1(GND_net), .B0(GND_net), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n6894), .ROA16(n6893), 
            .ROA15(n6892), .ROA14(n6891), .ROA13(n6890), .ROA12(n6889), 
            .ROA11(n6888), .ROA10(n6887), .ROA9(n6886), .ROA8(n6885), 
            .ROA7(n6884), .ROA6(n6883), .ROA5(n6882), .ROA4(n6881), 
            .ROA3(n6880), .ROA2(n6879), .ROA1(n6878), .ROA0(n6877), 
            .ROB17(n6912), .ROB16(n6911), .ROB15(n6910), .ROB14(n6909), 
            .ROB13(n6908), .ROB12(n6907), .ROB11(n6906), .ROB10(n6905), 
            .ROB9(n6904), .ROB8(n6903), .ROB7(n6902), .ROB6(n6901), 
            .ROB5(n6900), .ROB4(n6899), .ROB3(n6898), .ROB2(n6897), 
            .ROB1(n6896), .ROB0(n6895), .P35(n6949), .P34(n6948), .P33(n6947), 
            .P32(n6946), .P31(n6945), .P30(n6944), .P29(n6943), .P28(n6942), 
            .P27(n6941), .P26(n6940), .P25(n6939), .P24(n6938), .P23(n6937), 
            .P22(n6936), .P21(n6935), .P20(n6934), .P19(n6933), .P18(n6932), 
            .P17(n6931), .P16(n6930), .P15(n6929), .P14(n6928), .P13(n6927), 
            .P12(n6926), .P11(n6925), .P10(n6924), .P9(n6923), .P8(n6922), 
            .P7(n6921), .P6(n6920), .P5(n6919), .P4(n6918), .P3(n6917), 
            .P2(n6916), .P1(n6915), .P0(n6914), .SIGNEDP(n6913));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam lat_mult_6.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_6.REG_INPUTA_CE = "CE3";
    defparam lat_mult_6.REG_INPUTA_RST = "RST3";
    defparam lat_mult_6.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTB_CE = "CE0";
    defparam lat_mult_6.REG_INPUTB_RST = "RST0";
    defparam lat_mult_6.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTC_CE = "CE0";
    defparam lat_mult_6.REG_INPUTC_RST = "RST0";
    defparam lat_mult_6.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_6.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_6.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_6.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_6.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_6.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_6.CLK0_DIV = "ENABLED";
    defparam lat_mult_6.CLK1_DIV = "ENABLED";
    defparam lat_mult_6.CLK2_DIV = "ENABLED";
    defparam lat_mult_6.CLK3_DIV = "ENABLED";
    defparam lat_mult_6.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_6.GSR = "DISABLED";
    defparam lat_mult_6.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_6.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_6.MULT_BYPASS = "DISABLED";
    defparam lat_mult_6.RESETMODE = "ASYNC";
    FD1P3AX b_s_res8_e3_e3__i1 (.D(n86_adj_1256), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5277));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i1.GSR = "DISABLED";
    MULT18X18D lat_mult_5 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(GND_net), .B16(n5197), .B15(n5198), 
            .B14(n5199), .B13(n5200), .B12(n5201), .B11(n5202), .B10(n5203), 
            .B9(n5204), .B8(n5205), .B7(n5206), .B6(n5207), .B5(n5208), 
            .B4(n5209), .B3(n5210), .B2(n5211), .B1(n5212), .B0(n5277), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n6821), .ROA16(n6820), 
            .ROA15(n6819), .ROA14(n6818), .ROA13(n6817), .ROA12(n6816), 
            .ROA11(n6815), .ROA10(n6814), .ROA9(n6813), .ROA8(n6812), 
            .ROA7(n6811), .ROA6(n6810), .ROA5(n6809), .ROA4(n6808), 
            .ROA3(n6807), .ROA2(n6806), .ROA1(n6805), .ROA0(n6804), 
            .ROB17(n6839), .ROB16(n6838), .ROB15(n6837), .ROB14(n6836), 
            .ROB13(n6835), .ROB12(n6834), .ROB11(n6833), .ROB10(n6832), 
            .ROB9(n6831), .ROB8(n6830), .ROB7(n6829), .ROB6(n6828), 
            .ROB5(n6827), .ROB4(n6826), .ROB3(n6825), .ROB2(n6824), 
            .ROB1(n6823), .ROB0(n6822), .P35(n6876), .P34(n6875), .P33(n6874), 
            .P32(n6873), .P31(n6872), .P30(n6871), .P29(n6870), .P28(n6869), 
            .P27(n6868), .P26(n6867), .P25(n6866), .P24(n6865), .P23(n6864), 
            .P22(n6863), .P21(n6862), .P20(n6861), .P19(n6860), .P18(n6859), 
            .P17(n6858), .P16(n6857), .P15(n6856), .P14(n6855), .P13(n6854), 
            .P12(n6853), .P11(n6852), .P10(n6851), .P9(n6850), .P8(n6849), 
            .P7(n6848), .P6(n6847), .P5(n6846), .P4(n6845), .P3(n6844), 
            .P2(n6843), .P1(n6842), .P0(n6841), .SIGNEDP(n6840));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam lat_mult_5.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_5.REG_INPUTA_CE = "CE3";
    defparam lat_mult_5.REG_INPUTA_RST = "RST3";
    defparam lat_mult_5.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTB_CE = "CE0";
    defparam lat_mult_5.REG_INPUTB_RST = "RST0";
    defparam lat_mult_5.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTC_CE = "CE0";
    defparam lat_mult_5.REG_INPUTC_RST = "RST0";
    defparam lat_mult_5.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_5.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_5.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_5.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_5.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_5.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_5.CLK0_DIV = "ENABLED";
    defparam lat_mult_5.CLK1_DIV = "ENABLED";
    defparam lat_mult_5.CLK2_DIV = "ENABLED";
    defparam lat_mult_5.CLK3_DIV = "ENABLED";
    defparam lat_mult_5.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_5.GSR = "DISABLED";
    defparam lat_mult_5.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_5.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_5.MULT_BYPASS = "DISABLED";
    defparam lat_mult_5.RESETMODE = "ASYNC";
    MULT18X18D prod_b__1_res7_mult_2 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(GND_net), .B16(n5197), .B15(n5198), 
            .B14(n5199), .B13(n5200), .B12(n5201), .B11(n5202), .B10(n5203), 
            .B9(n5204), .B8(n5205), .B7(n5206), .B6(n5207), .B5(n5208), 
            .B4(n5209), .B3(n5210), .B2(n5211), .B1(n5212), .B0(n5277), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n6748), .ROA16(n6747), 
            .ROA15(n6746), .ROA14(n6745), .ROA13(n6744), .ROA12(n6743), 
            .ROA11(n6742), .ROA10(n6741), .ROA9(n6740), .ROA8(n6739), 
            .ROA7(n6738), .ROA6(n6737), .ROA5(n6736), .ROA4(n6735), 
            .ROA3(n6734), .ROA2(n6733), .ROA1(n6732), .ROA0(n6731), 
            .ROB17(n6766), .ROB16(n6765), .ROB15(n6764), .ROB14(n6763), 
            .ROB13(n6762), .ROB12(n6761), .ROB11(n6760), .ROB10(n6759), 
            .ROB9(n6758), .ROB8(n6757), .ROB7(n6756), .ROB6(n6755), 
            .ROB5(n6754), .ROB4(n6753), .ROB3(n6752), .ROB2(n6751), 
            .ROB1(n6750), .ROB0(n6749), .P35(n6803), .P34(n6802), .P33(n6801), 
            .P32(n6800), .P31(n6799), .P30(n6798), .P29(n6797), .P28(n6796), 
            .P27(n6795), .P26(n6794), .P25(n6793), .P24(n6792), .P23(n6791), 
            .P22(n6790), .P21(n6789), .P20(n6788), .P19(n6787), .P18(n6786), 
            .P17(n6785), .P16(n6784), .P15(n6783), .P14(n6782), .P13(n6781), 
            .P12(n6780), .P11(n6779), .P10(n6778), .P9(n6777), .P8(n6776), 
            .P7(n6775), .P6(n6774), .P5(n6773), .P4(n6772), .P3(n6771), 
            .P2(n6770), .P1(n6769), .P0(n6768), .SIGNEDP(n6767));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam prod_b__1_res7_mult_2.REG_INPUTA_CE = "CE3";
    defparam prod_b__1_res7_mult_2.REG_INPUTA_RST = "RST3";
    defparam prod_b__1_res7_mult_2.REG_INPUTB_CLK = "NONE";
    defparam prod_b__1_res7_mult_2.REG_INPUTB_CE = "CE0";
    defparam prod_b__1_res7_mult_2.REG_INPUTB_RST = "RST0";
    defparam prod_b__1_res7_mult_2.REG_INPUTC_CLK = "NONE";
    defparam prod_b__1_res7_mult_2.REG_INPUTC_CE = "CE0";
    defparam prod_b__1_res7_mult_2.REG_INPUTC_RST = "RST0";
    defparam prod_b__1_res7_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam prod_b__1_res7_mult_2.REG_PIPELINE_CE = "CE0";
    defparam prod_b__1_res7_mult_2.REG_PIPELINE_RST = "RST0";
    defparam prod_b__1_res7_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam prod_b__1_res7_mult_2.REG_OUTPUT_CE = "CE0";
    defparam prod_b__1_res7_mult_2.REG_OUTPUT_RST = "RST0";
    defparam prod_b__1_res7_mult_2.CLK0_DIV = "ENABLED";
    defparam prod_b__1_res7_mult_2.CLK1_DIV = "ENABLED";
    defparam prod_b__1_res7_mult_2.CLK2_DIV = "ENABLED";
    defparam prod_b__1_res7_mult_2.CLK3_DIV = "ENABLED";
    defparam prod_b__1_res7_mult_2.HIGHSPEED_CLK = "NONE";
    defparam prod_b__1_res7_mult_2.GSR = "DISABLED";
    defparam prod_b__1_res7_mult_2.CAS_MATCH_REG = "FALSE";
    defparam prod_b__1_res7_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam prod_b__1_res7_mult_2.MULT_BYPASS = "DISABLED";
    defparam prod_b__1_res7_mult_2.RESETMODE = "ASYNC";
    ALU54B lat_alu_4 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n6553), .SIGNEDIB(n6626), .SIGNEDCIN(n6699), .A35(n6552), 
           .A34(n6551), .A33(n6550), .A32(n6549), .A31(n6548), .A30(n6547), 
           .A29(n6546), .A28(n6545), .A27(n6544), .A26(n6543), .A25(n6542), 
           .A24(n6541), .A23(n6540), .A22(n6539), .A21(n6538), .A20(n6537), 
           .A19(n6536), .A18(n6535), .A17(n6534), .A16(n6533), .A15(n6532), 
           .A14(n6531), .A13(n6530), .A12(n6529), .A11(n6528), .A10(n6527), 
           .A9(n6526), .A8(n6525), .A7(n6524), .A6(n6523), .A5(n6522), 
           .A4(n6521), .A3(n6520), .A2(n6519), .A1(n6518), .A0(n6517), 
           .B35(n6625), .B34(n6624), .B33(n6623), .B32(n6622), .B31(n6621), 
           .B30(n6620), .B29(n6619), .B28(n6618), .B27(n6617), .B26(n6616), 
           .B25(n6615), .B24(n6614), .B23(n6613), .B22(n6612), .B21(n6611), 
           .B20(n6610), .B19(n6609), .B18(n6608), .B17(n6607), .B16(n6606), 
           .B15(n6605), .B14(n6604), .B13(n6603), .B12(n6602), .B11(n6601), 
           .B10(n6600), .B9(n6599), .B8(n6598), .B7(n6597), .B6(n6596), 
           .B5(n6595), .B4(n6594), .B3(n6593), .B2(n6592), .B1(n6591), 
           .B0(n6590), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n6589), .MA34(n6588), .MA33(n6587), .MA32(n6586), .MA31(n6585), 
           .MA30(n6584), .MA29(n6583), .MA28(n6582), .MA27(n6581), .MA26(n6580), 
           .MA25(n6579), .MA24(n6578), .MA23(n6577), .MA22(n6576), .MA21(n6575), 
           .MA20(n6574), .MA19(n6573), .MA18(n6572), .MA17(n6571), .MA16(n6570), 
           .MA15(n6569), .MA14(n6568), .MA13(n6567), .MA12(n6566), .MA11(n6565), 
           .MA10(n6564), .MA9(n6563), .MA8(n6562), .MA7(n6561), .MA6(n6560), 
           .MA5(n6559), .MA4(n6558), .MA3(n6557), .MA2(n6556), .MA1(n6555), 
           .MA0(n6554), .MB35(n6662), .MB34(n6661), .MB33(n6660), .MB32(n6659), 
           .MB31(n6658), .MB30(n6657), .MB29(n6656), .MB28(n6655), .MB27(n6654), 
           .MB26(n6653), .MB25(n6652), .MB24(n6651), .MB23(n6650), .MB22(n6649), 
           .MB21(n6648), .MB20(n6647), .MB19(n6646), .MB18(n6645), .MB17(n6644), 
           .MB16(n6643), .MB15(n6642), .MB14(n6641), .MB13(n6640), .MB12(n6639), 
           .MB11(n6638), .MB10(n6637), .MB9(n6636), .MB8(n6635), .MB7(n6634), 
           .MB6(n6633), .MB5(n6632), .MB4(n6631), .MB3(n6630), .MB2(n6629), 
           .MB1(n6628), .MB0(n6627), .CIN53(n6698), .CIN52(n6697), .CIN51(n6696), 
           .CIN50(n6695), .CIN49(n6694), .CIN48(n6693), .CIN47(n6692), 
           .CIN46(n6691), .CIN45(n6690), .CIN44(n6689), .CIN43(n6688), 
           .CIN42(n6687), .CIN41(n6686), .CIN40(n6685), .CIN39(n6684), 
           .CIN38(n6683), .CIN37(n6682), .CIN36(n6681), .CIN35(n6680), 
           .CIN34(n6679), .CIN33(n6678), .CIN32(n6677), .CIN31(n6676), 
           .CIN30(n6675), .CIN29(n6674), .CIN28(n6673), .CIN27(n6672), 
           .CIN26(n6671), .CIN25(n6670), .CIN24(n6669), .CIN23(n6668), 
           .CIN22(n6667), .CIN21(n6666), .CIN20(n6665), .CIN19(n6664), 
           .CIN18(n6663), .CIN17(n177_adj_1180), .CIN16(n178_adj_1179), 
           .CIN15(n179_adj_1178), .CIN14(n6356), .CIN13(n6357), .CIN12(n6358), 
           .CIN11(n6359), .CIN10(n6360), .CIN9(n6361), .CIN8(n6362), 
           .CIN7(n6363), .CIN6(n6364), .CIN5(n6365), .CIN4(n6366), .CIN3(n6367), 
           .CIN2(n6368), .CIN1(n6369), .CIN0(n6370), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R29(n147_adj_1210), .R28(n148_adj_1209), 
           .R27(n149_adj_1208), .R26(n150_adj_1207), .R25(n151_adj_1206), 
           .R24(n152_adj_1205), .R23(n153_adj_1204), .R22(n154_adj_1203), 
           .R21(n155_adj_1202), .R20(n156_adj_1201), .R19(n157_adj_1200), 
           .R18(n158_adj_1199), .R17(n159_adj_1198), .R16(n160_adj_1197), 
           .R15(n161_adj_1196), .R14(n162_adj_1195), .R13(n163_adj_1194), 
           .R12(n164_adj_1193), .R11(n165_adj_1192), .R10(n166_adj_1191), 
           .R9(n167_adj_1190), .R8(n168_adj_1189), .R7(n169_adj_1188), 
           .R6(n170_adj_1187), .R5(n171_adj_1186), .R4(n172_adj_1185), 
           .R3(n173_adj_1184), .R2(n174_adj_1183), .R1(n175_adj_1182), 
           .R0(n176_adj_1181));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam lat_alu_4.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_4.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_4.REG_FLAG_CLK = "NONE";
    defparam lat_alu_4.REG_FLAG_CE = "CE0";
    defparam lat_alu_4.REG_FLAG_RST = "RST0";
    defparam lat_alu_4.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASK01 = "0x00000000000000";
    defparam lat_alu_4.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_4.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_4.CLK0_DIV = "ENABLED";
    defparam lat_alu_4.CLK1_DIV = "ENABLED";
    defparam lat_alu_4.CLK2_DIV = "ENABLED";
    defparam lat_alu_4.CLK3_DIV = "ENABLED";
    defparam lat_alu_4.MCPAT = "0x00000000000000";
    defparam lat_alu_4.MASKPAT = "0x00000000000000";
    defparam lat_alu_4.RNDPAT = "0x00000000000000";
    defparam lat_alu_4.GSR = "DISABLED";
    defparam lat_alu_4.RESETMODE = "SYNC";
    defparam lat_alu_4.MULT9_MODE = "DISABLED";
    defparam lat_alu_4.LEGACY = "DISABLED";
    ALU54B lat_alu_8 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n6767), .SIGNEDIB(n6840), .SIGNEDCIN(GND_net), .A35(n6766), 
           .A34(n6765), .A33(n6764), .A32(n6763), .A31(n6762), .A30(n6761), 
           .A29(n6760), .A28(n6759), .A27(n6758), .A26(n6757), .A25(n6756), 
           .A24(n6755), .A23(n6754), .A22(n6753), .A21(n6752), .A20(n6751), 
           .A19(n6750), .A18(n6749), .A17(n6748), .A16(n6747), .A15(n6746), 
           .A14(n6745), .A13(n6744), .A12(n6743), .A11(n6742), .A10(n6741), 
           .A9(n6740), .A8(n6739), .A7(n6738), .A6(n6737), .A5(n6736), 
           .A4(n6735), .A3(n6734), .A2(n6733), .A1(n6732), .A0(n6731), 
           .B35(n6839), .B34(n6838), .B33(n6837), .B32(n6836), .B31(n6835), 
           .B30(n6834), .B29(n6833), .B28(n6832), .B27(n6831), .B26(n6830), 
           .B25(n6829), .B24(n6828), .B23(n6827), .B22(n6826), .B21(n6825), 
           .B20(n6824), .B19(n6823), .B18(n6822), .B17(n6821), .B16(n6820), 
           .B15(n6819), .B14(n6818), .B13(n6817), .B12(n6816), .B11(n6815), 
           .B10(n6814), .B9(n6813), .B8(n6812), .B7(n6811), .B6(n6810), 
           .B5(n6809), .B4(n6808), .B3(n6807), .B2(n6806), .B1(n6805), 
           .B0(n6804), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n6803), .MA34(n6802), .MA33(n6801), .MA32(n6800), .MA31(n6799), 
           .MA30(n6798), .MA29(n6797), .MA28(n6796), .MA27(n6795), .MA26(n6794), 
           .MA25(n6793), .MA24(n6792), .MA23(n6791), .MA22(n6790), .MA21(n6789), 
           .MA20(n6788), .MA19(n6787), .MA18(n6786), .MA17(n6785), .MA16(n6784), 
           .MA15(n6783), .MA14(n6782), .MA13(n6781), .MA12(n6780), .MA11(n6779), 
           .MA10(n6778), .MA9(n6777), .MA8(n6776), .MA7(n6775), .MA6(n6774), 
           .MA5(n6773), .MA4(n6772), .MA3(n6771), .MA2(n6770), .MA1(n6769), 
           .MA0(n6768), .MB35(n6876), .MB34(n6875), .MB33(n6874), .MB32(n6873), 
           .MB31(n6872), .MB30(n6871), .MB29(n6870), .MB28(n6869), .MB27(n6868), 
           .MB26(n6867), .MB25(n6866), .MB24(n6865), .MB23(n6864), .MB22(n6863), 
           .MB21(n6862), .MB20(n6861), .MB19(n6860), .MB18(n6859), .MB17(n6858), 
           .MB16(n6857), .MB15(n6856), .MB14(n6855), .MB13(n6854), .MB12(n6853), 
           .MB11(n6852), .MB10(n6851), .MB9(n6850), .MB8(n6849), .MB7(n6848), 
           .MB6(n6847), .MB5(n6846), .MB4(n6845), .MB3(n6844), .MB2(n6843), 
           .MB1(n6842), .MB0(n6841), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n7058), 
           .R52(n7057), .R51(n7056), .R50(n7055), .R49(n7054), .R48(n7053), 
           .R47(n7052), .R46(n7051), .R45(n7050), .R44(n7049), .R43(n7048), 
           .R42(n7047), .R41(n7046), .R40(n7045), .R39(n7044), .R38(n7043), 
           .R37(n7042), .R36(n7041), .R35(n7040), .R34(n7039), .R33(n7038), 
           .R32(n7037), .R31(n7036), .R30(n7035), .R29(n7034), .R28(n7033), 
           .R27(n7032), .R26(n7031), .R25(n7030), .R24(n7029), .R23(n7028), 
           .R22(n7027), .R21(n7026), .R20(n7025), .R19(n7024), .R18(n7023), 
           .R17(n177), .R16(n178_adj_1117), .R15(n179_adj_1116), .R14(n6716), 
           .R13(n6717), .R12(n6718), .R11(n6719), .R10(n6720), .R9(n6721), 
           .R8(n6722), .R7(n6723), .R6(n6724), .R5(n6725), .R4(n6726), 
           .R3(n6727), .R2(n6728), .R1(n6729), .R0(n6730), .SIGNEDR(n7059));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam lat_alu_8.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_8.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_8.REG_FLAG_CLK = "NONE";
    defparam lat_alu_8.REG_FLAG_CE = "CE0";
    defparam lat_alu_8.REG_FLAG_RST = "RST0";
    defparam lat_alu_8.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASK01 = "0x00000000000000";
    defparam lat_alu_8.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_8.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_8.CLK0_DIV = "ENABLED";
    defparam lat_alu_8.CLK1_DIV = "ENABLED";
    defparam lat_alu_8.CLK2_DIV = "ENABLED";
    defparam lat_alu_8.CLK3_DIV = "ENABLED";
    defparam lat_alu_8.MCPAT = "0x00000000000000";
    defparam lat_alu_8.MASKPAT = "0x00000000000000";
    defparam lat_alu_8.RNDPAT = "0x00000000000000";
    defparam lat_alu_8.GSR = "DISABLED";
    defparam lat_alu_8.RESETMODE = "SYNC";
    defparam lat_alu_8.MULT9_MODE = "DISABLED";
    defparam lat_alu_8.LEGACY = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i1 (.D(n179_adj_1227), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_c[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i1.GSR = "DISABLED";
    MULT18X18D mult_3 (.A17(d_c_15), .A16(d_c_15), .A15(d_c_15), .A14(d_c_14), 
            .A13(d_c_13), .A12(d_c_12), .A11(d_c_11), .A10(d_c_10), 
            .A9(d_c_9), .A8(d_c_8), .A7(d_c_7), .A6(d_c_6), .A5(d_c_5), 
            .A4(d_c_4), .A3(d_c_3), .A2(d_c_2), .A1(d_c_1), .A0(d_c_0), 
            .B17(a_c_15), .B16(a_c_15), .B15(a_c_15), .B14(a_c_14), 
            .B13(a_c_13), .B12(a_c_12), .B11(a_c_11), .B10(a_c_10), 
            .B9(a_c_9), .B8(a_c_8), .B7(a_c_7), .B6(a_c_6), .B5(a_c_5), 
            .B4(a_c_4), .B3(a_c_3), .B2(a_c_2), .B1(a_c_1), .B0(a_c_0), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(n8817), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P31(n37), .P30(n38), 
            .P29(n39), .P28(n40), .P27(n41), .P26(n42), .P25(n43), 
            .P24(n44), .P23(n45), .P22(n46), .P21(n47), .P20(n48), 
            .P19(n49), .P18(n50), .P17(n51), .P16(n52), .P15(n53), 
            .P14(n54), .P13(n55), .P12(n56), .P11(n57), .P10(n58), 
            .P9(n59), .P8(n60), .P7(n61), .P6(n62), .P5(n63), .P4(n64), 
            .P3(n65), .P2(n66), .P1(n67), .P0(n68));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:52])
    defparam mult_3.REG_INPUTA_CLK = "CLK3";
    defparam mult_3.REG_INPUTA_CE = "CE3";
    defparam mult_3.REG_INPUTA_RST = "RST3";
    defparam mult_3.REG_INPUTB_CLK = "CLK3";
    defparam mult_3.REG_INPUTB_CE = "CE3";
    defparam mult_3.REG_INPUTB_RST = "RST3";
    defparam mult_3.REG_INPUTC_CLK = "NONE";
    defparam mult_3.REG_INPUTC_CE = "CE0";
    defparam mult_3.REG_INPUTC_RST = "RST0";
    defparam mult_3.REG_PIPELINE_CLK = "NONE";
    defparam mult_3.REG_PIPELINE_CE = "CE0";
    defparam mult_3.REG_PIPELINE_RST = "RST0";
    defparam mult_3.REG_OUTPUT_CLK = "NONE";
    defparam mult_3.REG_OUTPUT_CE = "CE0";
    defparam mult_3.REG_OUTPUT_RST = "RST0";
    defparam mult_3.CLK0_DIV = "ENABLED";
    defparam mult_3.CLK1_DIV = "ENABLED";
    defparam mult_3.CLK2_DIV = "ENABLED";
    defparam mult_3.CLK3_DIV = "ENABLED";
    defparam mult_3.HIGHSPEED_CLK = "NONE";
    defparam mult_3.GSR = "DISABLED";
    defparam mult_3.CAS_MATCH_REG = "FALSE";
    defparam mult_3.SOURCEB_MODE = "B_SHIFT";
    defparam mult_3.MULT_BYPASS = "DISABLED";
    defparam mult_3.RESETMODE = "ASYNC";
    LUT4 i18_4_lut (.A(det_q4_28_31__N_551[19]), .B(det_q4_28_31__N_551[5]), 
         .C(det_q4_28_31__N_551[8]), .D(det_q4_28_31__N_551[6]), .Z(n50_adj_1229)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i18_4_lut.init = 16'hfffe;
    MULT18X18D mult_4 (.A17(c_c_15), .A16(c_c_15), .A15(c_c_15), .A14(c_c_14), 
            .A13(c_c_13), .A12(c_c_12), .A11(c_c_11), .A10(c_c_10), 
            .A9(c_c_9), .A8(c_c_8), .A7(c_c_7), .A6(c_c_6), .A5(c_c_5), 
            .A4(c_c_4), .A3(c_c_3), .A2(c_c_2), .A1(c_c_1), .A0(c_c_0), 
            .B17(b_c_15), .B16(b_c_15), .B15(b_c_15), .B14(b_c_14), 
            .B13(b_c_13), .B12(b_c_12), .B11(b_c_11), .B10(b_c_10), 
            .B9(b_c_9), .B8(b_c_8), .B7(b_c_7), .B6(b_c_6), .B5(b_c_5), 
            .B4(b_c_4), .B3(b_c_3), .B2(b_c_2), .B1(b_c_1), .B0(b_c_0), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(n8817), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P31(n70), .P30(n71), 
            .P29(n72), .P28(n73), .P27(n74), .P26(n75), .P25(n76), 
            .P24(n77), .P23(n78), .P22(n79), .P21(n80), .P20(n81), 
            .P19(n82), .P18(n83), .P17(n84), .P16(n85), .P15(n86), 
            .P14(n87), .P13(n88), .P12(n89), .P11(n90), .P10(n91), 
            .P9(n92), .P8(n93), .P7(n94), .P6(n95), .P5(n96), .P4(n97), 
            .P3(n98), .P2(n99), .P1(n100), .P0(n101));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[55:70])
    defparam mult_4.REG_INPUTA_CLK = "CLK3";
    defparam mult_4.REG_INPUTA_CE = "CE3";
    defparam mult_4.REG_INPUTA_RST = "RST3";
    defparam mult_4.REG_INPUTB_CLK = "CLK3";
    defparam mult_4.REG_INPUTB_CE = "CE3";
    defparam mult_4.REG_INPUTB_RST = "RST3";
    defparam mult_4.REG_INPUTC_CLK = "NONE";
    defparam mult_4.REG_INPUTC_CE = "CE0";
    defparam mult_4.REG_INPUTC_RST = "RST0";
    defparam mult_4.REG_PIPELINE_CLK = "NONE";
    defparam mult_4.REG_PIPELINE_CE = "CE0";
    defparam mult_4.REG_PIPELINE_RST = "RST0";
    defparam mult_4.REG_OUTPUT_CLK = "NONE";
    defparam mult_4.REG_OUTPUT_CE = "CE0";
    defparam mult_4.REG_OUTPUT_RST = "RST0";
    defparam mult_4.CLK0_DIV = "ENABLED";
    defparam mult_4.CLK1_DIV = "ENABLED";
    defparam mult_4.CLK2_DIV = "ENABLED";
    defparam mult_4.CLK3_DIV = "ENABLED";
    defparam mult_4.HIGHSPEED_CLK = "NONE";
    defparam mult_4.GSR = "DISABLED";
    defparam mult_4.CAS_MATCH_REG = "FALSE";
    defparam mult_4.SOURCEB_MODE = "B_SHIFT";
    defparam mult_4.MULT_BYPASS = "DISABLED";
    defparam mult_4.RESETMODE = "ASYNC";
    LUT4 i21_4_lut (.A(det_q4_28_31__N_551[7]), .B(det_q4_28_31__N_551[30]), 
         .C(det_q4_28_31__N_551[14]), .D(det_q4_28_31__N_551[17]), .Z(n53_adj_1114)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i28_4_lut (.A(n55_adj_1297), .B(det_q4_28_31__N_551[18]), .C(n48_adj_1231), 
         .D(det_q4_28_31__N_551[2]), .Z(n60_adj_1115)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(det_q4_28_31__N_551[9]), .B(det_q4_28_31__N_551[26]), 
         .Z(n43_adj_1238)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i11_2_lut.init = 16'heeee;
    FD1P3AX d_inv_reg_res2_i0_i1 (.D(d_inv_15__N_535[32]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i1.GSR = "ENABLED";
    MULT18X18D lat_mult_11 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(GND_net), .B16(GND_net), 
            .B15(GND_net), .B14(GND_net), .B13(GND_net), .B12(GND_net), 
            .B11(GND_net), .B10(GND_net), .B9(GND_net), .B8(GND_net), 
            .B7(GND_net), .B6(GND_net), .B5(GND_net), .B4(GND_net), 
            .B3(GND_net), .B2(GND_net), .B1(GND_net), .B0(GND_net), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n7254), .ROA16(n7253), 
            .ROA15(n7252), .ROA14(n7251), .ROA13(n7250), .ROA12(n7249), 
            .ROA11(n7248), .ROA10(n7247), .ROA9(n7246), .ROA8(n7245), 
            .ROA7(n7244), .ROA6(n7243), .ROA5(n7242), .ROA4(n7241), 
            .ROA3(n7240), .ROA2(n7239), .ROA1(n7238), .ROA0(n7237), 
            .ROB17(n7272), .ROB16(n7271), .ROB15(n7270), .ROB14(n7269), 
            .ROB13(n7268), .ROB12(n7267), .ROB11(n7266), .ROB10(n7265), 
            .ROB9(n7264), .ROB8(n7263), .ROB7(n7262), .ROB6(n7261), 
            .ROB5(n7260), .ROB4(n7259), .ROB3(n7258), .ROB2(n7257), 
            .ROB1(n7256), .ROB0(n7255), .P35(n7309), .P34(n7308), .P33(n7307), 
            .P32(n7306), .P31(n7305), .P30(n7304), .P29(n7303), .P28(n7302), 
            .P27(n7301), .P26(n7300), .P25(n7299), .P24(n7298), .P23(n7297), 
            .P22(n7296), .P21(n7295), .P20(n7294), .P19(n7293), .P18(n7292), 
            .P17(n7291), .P16(n7290), .P15(n7289), .P14(n7288), .P13(n7287), 
            .P12(n7286), .P11(n7285), .P10(n7284), .P9(n7283), .P8(n7282), 
            .P7(n7281), .P6(n7280), .P5(n7279), .P4(n7278), .P3(n7277), 
            .P2(n7276), .P1(n7275), .P0(n7274), .SIGNEDP(n7273));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam lat_mult_11.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_11.REG_INPUTA_CE = "CE3";
    defparam lat_mult_11.REG_INPUTA_RST = "RST3";
    defparam lat_mult_11.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTB_CE = "CE0";
    defparam lat_mult_11.REG_INPUTB_RST = "RST0";
    defparam lat_mult_11.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTC_CE = "CE0";
    defparam lat_mult_11.REG_INPUTC_RST = "RST0";
    defparam lat_mult_11.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_11.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_11.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_11.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_11.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_11.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_11.CLK0_DIV = "ENABLED";
    defparam lat_mult_11.CLK1_DIV = "ENABLED";
    defparam lat_mult_11.CLK2_DIV = "ENABLED";
    defparam lat_mult_11.CLK3_DIV = "ENABLED";
    defparam lat_mult_11.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_11.GSR = "DISABLED";
    defparam lat_mult_11.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_11.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_11.MULT_BYPASS = "DISABLED";
    defparam lat_mult_11.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_12 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(GND_net), .B16(GND_net), 
            .B15(GND_net), .B14(GND_net), .B13(GND_net), .B12(GND_net), 
            .B11(GND_net), .B10(GND_net), .B9(GND_net), .B8(GND_net), 
            .B7(GND_net), .B6(GND_net), .B5(GND_net), .B4(GND_net), 
            .B3(GND_net), .B2(GND_net), .B1(GND_net), .B0(GND_net), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n7327), .ROA16(n7326), 
            .ROA15(n7325), .ROA14(n7324), .ROA13(n7323), .ROA12(n7322), 
            .ROA11(n7321), .ROA10(n7320), .ROA9(n7319), .ROA8(n7318), 
            .ROA7(n7317), .ROA6(n7316), .ROA5(n7315), .ROA4(n7314), 
            .ROA3(n7313), .ROA2(n7312), .ROA1(n7311), .ROA0(n7310), 
            .ROB17(n7345), .ROB16(n7344), .ROB15(n7343), .ROB14(n7342), 
            .ROB13(n7341), .ROB12(n7340), .ROB11(n7339), .ROB10(n7338), 
            .ROB9(n7337), .ROB8(n7336), .ROB7(n7335), .ROB6(n7334), 
            .ROB5(n7333), .ROB4(n7332), .ROB3(n7331), .ROB2(n7330), 
            .ROB1(n7329), .ROB0(n7328), .P35(n7382), .P34(n7381), .P33(n7380), 
            .P32(n7379), .P31(n7378), .P30(n7377), .P29(n7376), .P28(n7375), 
            .P27(n7374), .P26(n7373), .P25(n7372), .P24(n7371), .P23(n7370), 
            .P22(n7369), .P21(n7368), .P20(n7367), .P19(n7366), .P18(n7365), 
            .P17(n7364), .P16(n7363), .P15(n7362), .P14(n7361), .P13(n7360), 
            .P12(n7359), .P11(n7358), .P10(n7357), .P9(n7356), .P8(n7355), 
            .P7(n7354), .P6(n7353), .P5(n7352), .P4(n7351), .P3(n7350), 
            .P2(n7349), .P1(n7348), .P0(n7347), .SIGNEDP(n7346));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam lat_mult_12.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_12.REG_INPUTA_CE = "CE3";
    defparam lat_mult_12.REG_INPUTA_RST = "RST3";
    defparam lat_mult_12.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTB_CE = "CE0";
    defparam lat_mult_12.REG_INPUTB_RST = "RST0";
    defparam lat_mult_12.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTC_CE = "CE0";
    defparam lat_mult_12.REG_INPUTC_RST = "RST0";
    defparam lat_mult_12.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_12.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_12.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_12.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_12.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_12.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_12.CLK0_DIV = "ENABLED";
    defparam lat_mult_12.CLK1_DIV = "ENABLED";
    defparam lat_mult_12.CLK2_DIV = "ENABLED";
    defparam lat_mult_12.CLK3_DIV = "ENABLED";
    defparam lat_mult_12.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_12.GSR = "DISABLED";
    defparam lat_mult_12.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_12.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_12.MULT_BYPASS = "DISABLED";
    defparam lat_mult_12.RESETMODE = "ASYNC";
    FD1P3AX prod_d__3_res11_e3__i33 (.D(n147_adj_1175), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i33.GSR = "DISABLED";
    FD1P3AX b_inv_reg_res4_i0_i1 (.D(b_inv_15__N_503[32]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i1.GSR = "ENABLED";
    LUT4 i12_2_lut (.A(det_q4_28_31__N_551[1]), .B(det_q4_28_31__N_551[4]), 
         .Z(n44_adj_1237)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i12_2_lut.init = 16'heeee;
    ALU54B lat_alu_13 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n7127), .SIGNEDIB(n7200), .SIGNEDCIN(GND_net), .A35(n7126), 
           .A34(n7125), .A33(n7124), .A32(n7123), .A31(n7122), .A30(n7121), 
           .A29(n7120), .A28(n7119), .A27(n7118), .A26(n7117), .A25(n7116), 
           .A24(n7115), .A23(n7114), .A22(n7113), .A21(n7112), .A20(n7111), 
           .A19(n7110), .A18(n7109), .A17(n7108), .A16(n7107), .A15(n7106), 
           .A14(n7105), .A13(n7104), .A12(n7103), .A11(n7102), .A10(n7101), 
           .A9(n7100), .A8(n7099), .A7(n7098), .A6(n7097), .A5(n7096), 
           .A4(n7095), .A3(n7094), .A2(n7093), .A1(n7092), .A0(n7091), 
           .B35(n7199), .B34(n7198), .B33(n7197), .B32(n7196), .B31(n7195), 
           .B30(n7194), .B29(n7193), .B28(n7192), .B27(n7191), .B26(n7190), 
           .B25(n7189), .B24(n7188), .B23(n7187), .B22(n7186), .B21(n7185), 
           .B20(n7184), .B19(n7183), .B18(n7182), .B17(n7181), .B16(n7180), 
           .B15(n7179), .B14(n7178), .B13(n7177), .B12(n7176), .B11(n7175), 
           .B10(n7174), .B9(n7173), .B8(n7172), .B7(n7171), .B6(n7170), 
           .B5(n7169), .B4(n7168), .B3(n7167), .B2(n7166), .B1(n7165), 
           .B0(n7164), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n7163), .MA34(n7162), .MA33(n7161), .MA32(n7160), .MA31(n7159), 
           .MA30(n7158), .MA29(n7157), .MA28(n7156), .MA27(n7155), .MA26(n7154), 
           .MA25(n7153), .MA24(n7152), .MA23(n7151), .MA22(n7150), .MA21(n7149), 
           .MA20(n7148), .MA19(n7147), .MA18(n7146), .MA17(n7145), .MA16(n7144), 
           .MA15(n7143), .MA14(n7142), .MA13(n7141), .MA12(n7140), .MA11(n7139), 
           .MA10(n7138), .MA9(n7137), .MA8(n7136), .MA7(n7135), .MA6(n7134), 
           .MA5(n7133), .MA4(n7132), .MA3(n7131), .MA2(n7130), .MA1(n7129), 
           .MA0(n7128), .MB35(n7236), .MB34(n7235), .MB33(n7234), .MB32(n7233), 
           .MB31(n7232), .MB30(n7231), .MB29(n7230), .MB28(n7229), .MB27(n7228), 
           .MB26(n7227), .MB25(n7226), .MB24(n7225), .MB23(n7224), .MB22(n7223), 
           .MB21(n7222), .MB20(n7221), .MB19(n7220), .MB18(n7219), .MB17(n7218), 
           .MB16(n7217), .MB15(n7216), .MB14(n7215), .MB13(n7214), .MB12(n7213), 
           .MB11(n7212), .MB10(n7211), .MB9(n7210), .MB8(n7209), .MB7(n7208), 
           .MB6(n7207), .MB5(n7206), .MB4(n7205), .MB3(n7204), .MB2(n7203), 
           .MB1(n7202), .MB0(n7201), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n7418), 
           .R52(n7417), .R51(n7416), .R50(n7415), .R49(n7414), .R48(n7413), 
           .R47(n7412), .R46(n7411), .R45(n7410), .R44(n7409), .R43(n7408), 
           .R42(n7407), .R41(n7406), .R40(n7405), .R39(n7404), .R38(n7403), 
           .R37(n7402), .R36(n7401), .R35(n7400), .R34(n7399), .R33(n7398), 
           .R32(n7397), .R31(n7396), .R30(n7395), .R29(n7394), .R28(n7393), 
           .R27(n7392), .R26(n7391), .R25(n7390), .R24(n7389), .R23(n7388), 
           .R22(n7387), .R21(n7386), .R20(n7385), .R19(n7384), .R18(n7383), 
           .R17(n177_adj_1232), .R16(n178_adj_1228), .R15(n179_adj_1227), 
           .R14(n7076), .R13(n7077), .R12(n7078), .R11(n7079), .R10(n7080), 
           .R9(n7081), .R8(n7082), .R7(n7083), .R6(n7084), .R5(n7085), 
           .R4(n7086), .R3(n7087), .R2(n7088), .R1(n7089), .R0(n7090), 
           .SIGNEDR(n7419));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam lat_alu_13.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_13.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_13.REG_FLAG_CLK = "NONE";
    defparam lat_alu_13.REG_FLAG_CE = "CE0";
    defparam lat_alu_13.REG_FLAG_RST = "RST0";
    defparam lat_alu_13.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASK01 = "0x00000000000000";
    defparam lat_alu_13.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_13.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_13.CLK0_DIV = "ENABLED";
    defparam lat_alu_13.CLK1_DIV = "ENABLED";
    defparam lat_alu_13.CLK2_DIV = "ENABLED";
    defparam lat_alu_13.CLK3_DIV = "ENABLED";
    defparam lat_alu_13.MCPAT = "0x00000000000000";
    defparam lat_alu_13.MASKPAT = "0x00000000000000";
    defparam lat_alu_13.RNDPAT = "0x00000000000000";
    defparam lat_alu_13.GSR = "DISABLED";
    defparam lat_alu_13.RESETMODE = "SYNC";
    defparam lat_alu_13.MULT9_MODE = "DISABLED";
    defparam lat_alu_13.LEGACY = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i1 (.D(n179_adj_1116), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i1.GSR = "DISABLED";
    ALU54B lat_alu_14 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n7273), .SIGNEDIB(n7346), .SIGNEDCIN(n7419), .A35(n7272), 
           .A34(n7271), .A33(n7270), .A32(n7269), .A31(n7268), .A30(n7267), 
           .A29(n7266), .A28(n7265), .A27(n7264), .A26(n7263), .A25(n7262), 
           .A24(n7261), .A23(n7260), .A22(n7259), .A21(n7258), .A20(n7257), 
           .A19(n7256), .A18(n7255), .A17(n7254), .A16(n7253), .A15(n7252), 
           .A14(n7251), .A13(n7250), .A12(n7249), .A11(n7248), .A10(n7247), 
           .A9(n7246), .A8(n7245), .A7(n7244), .A6(n7243), .A5(n7242), 
           .A4(n7241), .A3(n7240), .A2(n7239), .A1(n7238), .A0(n7237), 
           .B35(n7345), .B34(n7344), .B33(n7343), .B32(n7342), .B31(n7341), 
           .B30(n7340), .B29(n7339), .B28(n7338), .B27(n7337), .B26(n7336), 
           .B25(n7335), .B24(n7334), .B23(n7333), .B22(n7332), .B21(n7331), 
           .B20(n7330), .B19(n7329), .B18(n7328), .B17(n7327), .B16(n7326), 
           .B15(n7325), .B14(n7324), .B13(n7323), .B12(n7322), .B11(n7321), 
           .B10(n7320), .B9(n7319), .B8(n7318), .B7(n7317), .B6(n7316), 
           .B5(n7315), .B4(n7314), .B3(n7313), .B2(n7312), .B1(n7311), 
           .B0(n7310), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n7309), .MA34(n7308), .MA33(n7307), .MA32(n7306), .MA31(n7305), 
           .MA30(n7304), .MA29(n7303), .MA28(n7302), .MA27(n7301), .MA26(n7300), 
           .MA25(n7299), .MA24(n7298), .MA23(n7297), .MA22(n7296), .MA21(n7295), 
           .MA20(n7294), .MA19(n7293), .MA18(n7292), .MA17(n7291), .MA16(n7290), 
           .MA15(n7289), .MA14(n7288), .MA13(n7287), .MA12(n7286), .MA11(n7285), 
           .MA10(n7284), .MA9(n7283), .MA8(n7282), .MA7(n7281), .MA6(n7280), 
           .MA5(n7279), .MA4(n7278), .MA3(n7277), .MA2(n7276), .MA1(n7275), 
           .MA0(n7274), .MB35(n7382), .MB34(n7381), .MB33(n7380), .MB32(n7379), 
           .MB31(n7378), .MB30(n7377), .MB29(n7376), .MB28(n7375), .MB27(n7374), 
           .MB26(n7373), .MB25(n7372), .MB24(n7371), .MB23(n7370), .MB22(n7369), 
           .MB21(n7368), .MB20(n7367), .MB19(n7366), .MB18(n7365), .MB17(n7364), 
           .MB16(n7363), .MB15(n7362), .MB14(n7361), .MB13(n7360), .MB12(n7359), 
           .MB11(n7358), .MB10(n7357), .MB9(n7356), .MB8(n7355), .MB7(n7354), 
           .MB6(n7353), .MB5(n7352), .MB4(n7351), .MB3(n7350), .MB2(n7349), 
           .MB1(n7348), .MB0(n7347), .CIN53(n7418), .CIN52(n7417), .CIN51(n7416), 
           .CIN50(n7415), .CIN49(n7414), .CIN48(n7413), .CIN47(n7412), 
           .CIN46(n7411), .CIN45(n7410), .CIN44(n7409), .CIN43(n7408), 
           .CIN42(n7407), .CIN41(n7406), .CIN40(n7405), .CIN39(n7404), 
           .CIN38(n7403), .CIN37(n7402), .CIN36(n7401), .CIN35(n7400), 
           .CIN34(n7399), .CIN33(n7398), .CIN32(n7397), .CIN31(n7396), 
           .CIN30(n7395), .CIN29(n7394), .CIN28(n7393), .CIN27(n7392), 
           .CIN26(n7391), .CIN25(n7390), .CIN24(n7389), .CIN23(n7388), 
           .CIN22(n7387), .CIN21(n7386), .CIN20(n7385), .CIN19(n7384), 
           .CIN18(n7383), .CIN17(n177_adj_1232), .CIN16(n178_adj_1228), 
           .CIN15(n179_adj_1227), .CIN14(n7076), .CIN13(n7077), .CIN12(n7078), 
           .CIN11(n7079), .CIN10(n7080), .CIN9(n7081), .CIN8(n7082), 
           .CIN7(n7083), .CIN6(n7084), .CIN5(n7085), .CIN4(n7086), .CIN3(n7087), 
           .CIN2(n7088), .CIN1(n7089), .CIN0(n7090), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R29(n147), .R28(n148), .R27(n149), 
           .R26(n150), .R25(n151), .R24(n152), .R23(n153), .R22(n154), 
           .R21(n155), .R20(n156), .R19(n157), .R18(n158), .R17(n159), 
           .R16(n160), .R15(n161), .R14(n162), .R13(n163), .R12(n164), 
           .R11(n165), .R10(n166), .R9(n167), .R8(n168), .R7(n169), 
           .R6(n170), .R5(n171), .R4(n172), .R3(n173), .R2(n174_adj_1235), 
           .R1(n175_adj_1234), .R0(n176_adj_1233));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam lat_alu_14.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_14.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_14.REG_FLAG_CLK = "NONE";
    defparam lat_alu_14.REG_FLAG_CE = "CE0";
    defparam lat_alu_14.REG_FLAG_RST = "RST0";
    defparam lat_alu_14.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASK01 = "0x00000000000000";
    defparam lat_alu_14.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_14.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_14.CLK0_DIV = "ENABLED";
    defparam lat_alu_14.CLK1_DIV = "ENABLED";
    defparam lat_alu_14.CLK2_DIV = "ENABLED";
    defparam lat_alu_14.CLK3_DIV = "ENABLED";
    defparam lat_alu_14.MCPAT = "0x00000000000000";
    defparam lat_alu_14.MASKPAT = "0x00000000000000";
    defparam lat_alu_14.RNDPAT = "0x00000000000000";
    defparam lat_alu_14.GSR = "DISABLED";
    defparam lat_alu_14.RESETMODE = "SYNC";
    defparam lat_alu_14.MULT9_MODE = "DISABLED";
    defparam lat_alu_14.LEGACY = "DISABLED";
    MULT18X18D prod_d__3_res11_mult_2 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(n68_adj_1176), .B16(n68_adj_1176), 
            .B15(n68_adj_1176), .B14(n102), .B13(n104), .B12(n106), 
            .B11(n108), .B10(n110), .B9(n112), .B8(n114), .B7(n116), 
            .B6(n118), .B5(n120), .B4(n122), .B3(n124), .B2(n126), 
            .B1(n128), .B0(n130), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n7468), 
            .ROA16(n7467), .ROA15(n7466), .ROA14(n7465), .ROA13(n7464), 
            .ROA12(n7463), .ROA11(n7462), .ROA10(n7461), .ROA9(n7460), 
            .ROA8(n7459), .ROA7(n7458), .ROA6(n7457), .ROA5(n7456), 
            .ROA4(n7455), .ROA3(n7454), .ROA2(n7453), .ROA1(n7452), 
            .ROA0(n7451), .ROB17(n7486), .ROB16(n7485), .ROB15(n7484), 
            .ROB14(n7483), .ROB13(n7482), .ROB12(n7481), .ROB11(n7480), 
            .ROB10(n7479), .ROB9(n7478), .ROB8(n7477), .ROB7(n7476), 
            .ROB6(n7475), .ROB5(n7474), .ROB4(n7473), .ROB3(n7472), 
            .ROB2(n7471), .ROB1(n7470), .ROB0(n7469), .P35(n7523), .P34(n7522), 
            .P33(n7521), .P32(n7520), .P31(n7519), .P30(n7518), .P29(n7517), 
            .P28(n7516), .P27(n7515), .P26(n7514), .P25(n7513), .P24(n7512), 
            .P23(n7511), .P22(n7510), .P21(n7509), .P20(n7508), .P19(n7507), 
            .P18(n7506), .P17(n7505), .P16(n7504), .P15(n7503), .P14(n7502), 
            .P13(n7501), .P12(n7500), .P11(n7499), .P10(n7498), .P9(n7497), 
            .P8(n7496), .P7(n7495), .P6(n7494), .P5(n7493), .P4(n7492), 
            .P3(n7491), .P2(n7490), .P1(n7489), .P0(n7488), .SIGNEDP(n7487));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam prod_d__3_res11_mult_2.REG_INPUTA_CE = "CE3";
    defparam prod_d__3_res11_mult_2.REG_INPUTA_RST = "RST3";
    defparam prod_d__3_res11_mult_2.REG_INPUTB_CLK = "NONE";
    defparam prod_d__3_res11_mult_2.REG_INPUTB_CE = "CE0";
    defparam prod_d__3_res11_mult_2.REG_INPUTB_RST = "RST0";
    defparam prod_d__3_res11_mult_2.REG_INPUTC_CLK = "NONE";
    defparam prod_d__3_res11_mult_2.REG_INPUTC_CE = "CE0";
    defparam prod_d__3_res11_mult_2.REG_INPUTC_RST = "RST0";
    defparam prod_d__3_res11_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam prod_d__3_res11_mult_2.REG_PIPELINE_CE = "CE0";
    defparam prod_d__3_res11_mult_2.REG_PIPELINE_RST = "RST0";
    defparam prod_d__3_res11_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam prod_d__3_res11_mult_2.REG_OUTPUT_CE = "CE0";
    defparam prod_d__3_res11_mult_2.REG_OUTPUT_RST = "RST0";
    defparam prod_d__3_res11_mult_2.CLK0_DIV = "ENABLED";
    defparam prod_d__3_res11_mult_2.CLK1_DIV = "ENABLED";
    defparam prod_d__3_res11_mult_2.CLK2_DIV = "ENABLED";
    defparam prod_d__3_res11_mult_2.CLK3_DIV = "ENABLED";
    defparam prod_d__3_res11_mult_2.HIGHSPEED_CLK = "NONE";
    defparam prod_d__3_res11_mult_2.GSR = "DISABLED";
    defparam prod_d__3_res11_mult_2.CAS_MATCH_REG = "FALSE";
    defparam prod_d__3_res11_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam prod_d__3_res11_mult_2.MULT_BYPASS = "DISABLED";
    defparam prod_d__3_res11_mult_2.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_15 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(n68_adj_1176), .B16(n68_adj_1176), 
            .B15(n68_adj_1176), .B14(n102), .B13(n104), .B12(n106), 
            .B11(n108), .B10(n110), .B9(n112), .B8(n114), .B7(n116), 
            .B6(n118), .B5(n120), .B4(n122), .B3(n124), .B2(n126), 
            .B1(n128), .B0(n130), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n7541), 
            .ROA16(n7540), .ROA15(n7539), .ROA14(n7538), .ROA13(n7537), 
            .ROA12(n7536), .ROA11(n7535), .ROA10(n7534), .ROA9(n7533), 
            .ROA8(n7532), .ROA7(n7531), .ROA6(n7530), .ROA5(n7529), 
            .ROA4(n7528), .ROA3(n7527), .ROA2(n7526), .ROA1(n7525), 
            .ROA0(n7524), .ROB17(n7559), .ROB16(n7558), .ROB15(n7557), 
            .ROB14(n7556), .ROB13(n7555), .ROB12(n7554), .ROB11(n7553), 
            .ROB10(n7552), .ROB9(n7551), .ROB8(n7550), .ROB7(n7549), 
            .ROB6(n7548), .ROB5(n7547), .ROB4(n7546), .ROB3(n7545), 
            .ROB2(n7544), .ROB1(n7543), .ROB0(n7542), .P35(n7596), .P34(n7595), 
            .P33(n7594), .P32(n7593), .P31(n7592), .P30(n7591), .P29(n7590), 
            .P28(n7589), .P27(n7588), .P26(n7587), .P25(n7586), .P24(n7585), 
            .P23(n7584), .P22(n7583), .P21(n7582), .P20(n7581), .P19(n7580), 
            .P18(n7579), .P17(n7578), .P16(n7577), .P15(n7576), .P14(n7575), 
            .P13(n7574), .P12(n7573), .P11(n7572), .P10(n7571), .P9(n7570), 
            .P8(n7569), .P7(n7568), .P6(n7567), .P5(n7566), .P4(n7565), 
            .P3(n7564), .P2(n7563), .P1(n7562), .P0(n7561), .SIGNEDP(n7560));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam lat_mult_15.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_15.REG_INPUTA_CE = "CE3";
    defparam lat_mult_15.REG_INPUTA_RST = "RST3";
    defparam lat_mult_15.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTB_CE = "CE0";
    defparam lat_mult_15.REG_INPUTB_RST = "RST0";
    defparam lat_mult_15.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTC_CE = "CE0";
    defparam lat_mult_15.REG_INPUTC_RST = "RST0";
    defparam lat_mult_15.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_15.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_15.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_15.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_15.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_15.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_15.CLK0_DIV = "ENABLED";
    defparam lat_mult_15.CLK1_DIV = "ENABLED";
    defparam lat_mult_15.CLK2_DIV = "ENABLED";
    defparam lat_mult_15.CLK3_DIV = "ENABLED";
    defparam lat_mult_15.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_15.GSR = "DISABLED";
    defparam lat_mult_15.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_15.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_15.MULT_BYPASS = "DISABLED";
    defparam lat_mult_15.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_16 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(n68_adj_1176), .B16(n68_adj_1176), 
            .B15(n68_adj_1176), .B14(n68_adj_1176), .B13(n68_adj_1176), 
            .B12(n68_adj_1176), .B11(n68_adj_1176), .B10(n68_adj_1176), 
            .B9(n68_adj_1176), .B8(n68_adj_1176), .B7(n68_adj_1176), .B6(n68_adj_1176), 
            .B5(n68_adj_1176), .B4(n68_adj_1176), .B3(n68_adj_1176), .B2(n68_adj_1176), 
            .B1(n68_adj_1176), .B0(n68_adj_1176), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n7614), .ROA16(n7613), .ROA15(n7612), .ROA14(n7611), 
            .ROA13(n7610), .ROA12(n7609), .ROA11(n7608), .ROA10(n7607), 
            .ROA9(n7606), .ROA8(n7605), .ROA7(n7604), .ROA6(n7603), 
            .ROA5(n7602), .ROA4(n7601), .ROA3(n7600), .ROA2(n7599), 
            .ROA1(n7598), .ROA0(n7597), .ROB17(n7632), .ROB16(n7631), 
            .ROB15(n7630), .ROB14(n7629), .ROB13(n7628), .ROB12(n7627), 
            .ROB11(n7626), .ROB10(n7625), .ROB9(n7624), .ROB8(n7623), 
            .ROB7(n7622), .ROB6(n7621), .ROB5(n7620), .ROB4(n7619), 
            .ROB3(n7618), .ROB2(n7617), .ROB1(n7616), .ROB0(n7615), 
            .P35(n7669), .P34(n7668), .P33(n7667), .P32(n7666), .P31(n7665), 
            .P30(n7664), .P29(n7663), .P28(n7662), .P27(n7661), .P26(n7660), 
            .P25(n7659), .P24(n7658), .P23(n7657), .P22(n7656), .P21(n7655), 
            .P20(n7654), .P19(n7653), .P18(n7652), .P17(n7651), .P16(n7650), 
            .P15(n7649), .P14(n7648), .P13(n7647), .P12(n7646), .P11(n7645), 
            .P10(n7644), .P9(n7643), .P8(n7642), .P7(n7641), .P6(n7640), 
            .P5(n7639), .P4(n7638), .P3(n7637), .P2(n7636), .P1(n7635), 
            .P0(n7634), .SIGNEDP(n7633));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam lat_mult_16.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_16.REG_INPUTA_CE = "CE3";
    defparam lat_mult_16.REG_INPUTA_RST = "RST3";
    defparam lat_mult_16.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTB_CE = "CE0";
    defparam lat_mult_16.REG_INPUTB_RST = "RST0";
    defparam lat_mult_16.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTC_CE = "CE0";
    defparam lat_mult_16.REG_INPUTC_RST = "RST0";
    defparam lat_mult_16.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_16.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_16.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_16.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_16.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_16.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_16.CLK0_DIV = "ENABLED";
    defparam lat_mult_16.CLK1_DIV = "ENABLED";
    defparam lat_mult_16.CLK2_DIV = "ENABLED";
    defparam lat_mult_16.CLK3_DIV = "ENABLED";
    defparam lat_mult_16.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_16.GSR = "DISABLED";
    defparam lat_mult_16.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_16.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_16.MULT_BYPASS = "DISABLED";
    defparam lat_mult_16.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_17 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(n68_adj_1176), .B16(n68_adj_1176), 
            .B15(n68_adj_1176), .B14(n68_adj_1176), .B13(n68_adj_1176), 
            .B12(n68_adj_1176), .B11(n68_adj_1176), .B10(n68_adj_1176), 
            .B9(n68_adj_1176), .B8(n68_adj_1176), .B7(n68_adj_1176), .B6(n68_adj_1176), 
            .B5(n68_adj_1176), .B4(n68_adj_1176), .B3(n68_adj_1176), .B2(n68_adj_1176), 
            .B1(n68_adj_1176), .B0(n68_adj_1176), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n7687), .ROA16(n7686), .ROA15(n7685), .ROA14(n7684), 
            .ROA13(n7683), .ROA12(n7682), .ROA11(n7681), .ROA10(n7680), 
            .ROA9(n7679), .ROA8(n7678), .ROA7(n7677), .ROA6(n7676), 
            .ROA5(n7675), .ROA4(n7674), .ROA3(n7673), .ROA2(n7672), 
            .ROA1(n7671), .ROA0(n7670), .ROB17(n7705), .ROB16(n7704), 
            .ROB15(n7703), .ROB14(n7702), .ROB13(n7701), .ROB12(n7700), 
            .ROB11(n7699), .ROB10(n7698), .ROB9(n7697), .ROB8(n7696), 
            .ROB7(n7695), .ROB6(n7694), .ROB5(n7693), .ROB4(n7692), 
            .ROB3(n7691), .ROB2(n7690), .ROB1(n7689), .ROB0(n7688), 
            .P35(n7742), .P34(n7741), .P33(n7740), .P32(n7739), .P31(n7738), 
            .P30(n7737), .P29(n7736), .P28(n7735), .P27(n7734), .P26(n7733), 
            .P25(n7732), .P24(n7731), .P23(n7730), .P22(n7729), .P21(n7728), 
            .P20(n7727), .P19(n7726), .P18(n7725), .P17(n7724), .P16(n7723), 
            .P15(n7722), .P14(n7721), .P13(n7720), .P12(n7719), .P11(n7718), 
            .P10(n7717), .P9(n7716), .P8(n7715), .P7(n7714), .P6(n7713), 
            .P5(n7712), .P4(n7711), .P3(n7710), .P2(n7709), .P1(n7708), 
            .P0(n7707), .SIGNEDP(n7706));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam lat_mult_17.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_17.REG_INPUTA_CE = "CE3";
    defparam lat_mult_17.REG_INPUTA_RST = "RST3";
    defparam lat_mult_17.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTB_CE = "CE0";
    defparam lat_mult_17.REG_INPUTB_RST = "RST0";
    defparam lat_mult_17.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTC_CE = "CE0";
    defparam lat_mult_17.REG_INPUTC_RST = "RST0";
    defparam lat_mult_17.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_17.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_17.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_17.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_17.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_17.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_17.CLK0_DIV = "ENABLED";
    defparam lat_mult_17.CLK1_DIV = "ENABLED";
    defparam lat_mult_17.CLK2_DIV = "ENABLED";
    defparam lat_mult_17.CLK3_DIV = "ENABLED";
    defparam lat_mult_17.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_17.GSR = "DISABLED";
    defparam lat_mult_17.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_17.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_17.MULT_BYPASS = "DISABLED";
    defparam lat_mult_17.RESETMODE = "ASYNC";
    ALU54B lat_alu_18 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n7487), .SIGNEDIB(n7560), .SIGNEDCIN(GND_net), .A35(n7486), 
           .A34(n7485), .A33(n7484), .A32(n7483), .A31(n7482), .A30(n7481), 
           .A29(n7480), .A28(n7479), .A27(n7478), .A26(n7477), .A25(n7476), 
           .A24(n7475), .A23(n7474), .A22(n7473), .A21(n7472), .A20(n7471), 
           .A19(n7470), .A18(n7469), .A17(n7468), .A16(n7467), .A15(n7466), 
           .A14(n7465), .A13(n7464), .A12(n7463), .A11(n7462), .A10(n7461), 
           .A9(n7460), .A8(n7459), .A7(n7458), .A6(n7457), .A5(n7456), 
           .A4(n7455), .A3(n7454), .A2(n7453), .A1(n7452), .A0(n7451), 
           .B35(n7559), .B34(n7558), .B33(n7557), .B32(n7556), .B31(n7555), 
           .B30(n7554), .B29(n7553), .B28(n7552), .B27(n7551), .B26(n7550), 
           .B25(n7549), .B24(n7548), .B23(n7547), .B22(n7546), .B21(n7545), 
           .B20(n7544), .B19(n7543), .B18(n7542), .B17(n7541), .B16(n7540), 
           .B15(n7539), .B14(n7538), .B13(n7537), .B12(n7536), .B11(n7535), 
           .B10(n7534), .B9(n7533), .B8(n7532), .B7(n7531), .B6(n7530), 
           .B5(n7529), .B4(n7528), .B3(n7527), .B2(n7526), .B1(n7525), 
           .B0(n7524), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n7523), .MA34(n7522), .MA33(n7521), .MA32(n7520), .MA31(n7519), 
           .MA30(n7518), .MA29(n7517), .MA28(n7516), .MA27(n7515), .MA26(n7514), 
           .MA25(n7513), .MA24(n7512), .MA23(n7511), .MA22(n7510), .MA21(n7509), 
           .MA20(n7508), .MA19(n7507), .MA18(n7506), .MA17(n7505), .MA16(n7504), 
           .MA15(n7503), .MA14(n7502), .MA13(n7501), .MA12(n7500), .MA11(n7499), 
           .MA10(n7498), .MA9(n7497), .MA8(n7496), .MA7(n7495), .MA6(n7494), 
           .MA5(n7493), .MA4(n7492), .MA3(n7491), .MA2(n7490), .MA1(n7489), 
           .MA0(n7488), .MB35(n7596), .MB34(n7595), .MB33(n7594), .MB32(n7593), 
           .MB31(n7592), .MB30(n7591), .MB29(n7590), .MB28(n7589), .MB27(n7588), 
           .MB26(n7587), .MB25(n7586), .MB24(n7585), .MB23(n7584), .MB22(n7583), 
           .MB21(n7582), .MB20(n7581), .MB19(n7580), .MB18(n7579), .MB17(n7578), 
           .MB16(n7577), .MB15(n7576), .MB14(n7575), .MB13(n7574), .MB12(n7573), 
           .MB11(n7572), .MB10(n7571), .MB9(n7570), .MB8(n7569), .MB7(n7568), 
           .MB6(n7567), .MB5(n7566), .MB4(n7565), .MB3(n7564), .MB2(n7563), 
           .MB1(n7562), .MB0(n7561), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n7778), 
           .R52(n7777), .R51(n7776), .R50(n7775), .R49(n7774), .R48(n7773), 
           .R47(n7772), .R46(n7771), .R45(n7770), .R44(n7769), .R43(n7768), 
           .R42(n7767), .R41(n7766), .R40(n7765), .R39(n7764), .R38(n7763), 
           .R37(n7762), .R36(n7761), .R35(n7760), .R34(n7759), .R33(n7758), 
           .R32(n7757), .R31(n7756), .R30(n7755), .R29(n7754), .R28(n7753), 
           .R27(n7752), .R26(n7751), .R25(n7750), .R24(n7749), .R23(n7748), 
           .R22(n7747), .R21(n7746), .R20(n7745), .R19(n7744), .R18(n7743), 
           .R17(n177_adj_1145), .R16(n178), .R15(n179), .R14(n7436), 
           .R13(n7437), .R12(n7438), .R11(n7439), .R10(n7440), .R9(n7441), 
           .R8(n7442), .R7(n7443), .R6(n7444), .R5(n7445), .R4(n7446), 
           .R3(n7447), .R2(n7448), .R1(n7449), .R0(n7450), .SIGNEDR(n7779));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam lat_alu_18.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_18.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_18.REG_FLAG_CLK = "NONE";
    defparam lat_alu_18.REG_FLAG_CE = "CE0";
    defparam lat_alu_18.REG_FLAG_RST = "RST0";
    defparam lat_alu_18.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASK01 = "0x00000000000000";
    defparam lat_alu_18.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_18.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_18.CLK0_DIV = "ENABLED";
    defparam lat_alu_18.CLK1_DIV = "ENABLED";
    defparam lat_alu_18.CLK2_DIV = "ENABLED";
    defparam lat_alu_18.CLK3_DIV = "ENABLED";
    defparam lat_alu_18.MCPAT = "0x00000000000000";
    defparam lat_alu_18.MASKPAT = "0x00000000000000";
    defparam lat_alu_18.RNDPAT = "0x00000000000000";
    defparam lat_alu_18.GSR = "DISABLED";
    defparam lat_alu_18.RESETMODE = "SYNC";
    defparam lat_alu_18.MULT9_MODE = "DISABLED";
    defparam lat_alu_18.LEGACY = "DISABLED";
    ALU54B lat_alu_19 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n7633), .SIGNEDIB(n7706), .SIGNEDCIN(n7779), .A35(n7632), 
           .A34(n7631), .A33(n7630), .A32(n7629), .A31(n7628), .A30(n7627), 
           .A29(n7626), .A28(n7625), .A27(n7624), .A26(n7623), .A25(n7622), 
           .A24(n7621), .A23(n7620), .A22(n7619), .A21(n7618), .A20(n7617), 
           .A19(n7616), .A18(n7615), .A17(n7614), .A16(n7613), .A15(n7612), 
           .A14(n7611), .A13(n7610), .A12(n7609), .A11(n7608), .A10(n7607), 
           .A9(n7606), .A8(n7605), .A7(n7604), .A6(n7603), .A5(n7602), 
           .A4(n7601), .A3(n7600), .A2(n7599), .A1(n7598), .A0(n7597), 
           .B35(n7705), .B34(n7704), .B33(n7703), .B32(n7702), .B31(n7701), 
           .B30(n7700), .B29(n7699), .B28(n7698), .B27(n7697), .B26(n7696), 
           .B25(n7695), .B24(n7694), .B23(n7693), .B22(n7692), .B21(n7691), 
           .B20(n7690), .B19(n7689), .B18(n7688), .B17(n7687), .B16(n7686), 
           .B15(n7685), .B14(n7684), .B13(n7683), .B12(n7682), .B11(n7681), 
           .B10(n7680), .B9(n7679), .B8(n7678), .B7(n7677), .B6(n7676), 
           .B5(n7675), .B4(n7674), .B3(n7673), .B2(n7672), .B1(n7671), 
           .B0(n7670), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n7669), .MA34(n7668), .MA33(n7667), .MA32(n7666), .MA31(n7665), 
           .MA30(n7664), .MA29(n7663), .MA28(n7662), .MA27(n7661), .MA26(n7660), 
           .MA25(n7659), .MA24(n7658), .MA23(n7657), .MA22(n7656), .MA21(n7655), 
           .MA20(n7654), .MA19(n7653), .MA18(n7652), .MA17(n7651), .MA16(n7650), 
           .MA15(n7649), .MA14(n7648), .MA13(n7647), .MA12(n7646), .MA11(n7645), 
           .MA10(n7644), .MA9(n7643), .MA8(n7642), .MA7(n7641), .MA6(n7640), 
           .MA5(n7639), .MA4(n7638), .MA3(n7637), .MA2(n7636), .MA1(n7635), 
           .MA0(n7634), .MB35(n7742), .MB34(n7741), .MB33(n7740), .MB32(n7739), 
           .MB31(n7738), .MB30(n7737), .MB29(n7736), .MB28(n7735), .MB27(n7734), 
           .MB26(n7733), .MB25(n7732), .MB24(n7731), .MB23(n7730), .MB22(n7729), 
           .MB21(n7728), .MB20(n7727), .MB19(n7726), .MB18(n7725), .MB17(n7724), 
           .MB16(n7723), .MB15(n7722), .MB14(n7721), .MB13(n7720), .MB12(n7719), 
           .MB11(n7718), .MB10(n7717), .MB9(n7716), .MB8(n7715), .MB7(n7714), 
           .MB6(n7713), .MB5(n7712), .MB4(n7711), .MB3(n7710), .MB2(n7709), 
           .MB1(n7708), .MB0(n7707), .CIN53(n7778), .CIN52(n7777), .CIN51(n7776), 
           .CIN50(n7775), .CIN49(n7774), .CIN48(n7773), .CIN47(n7772), 
           .CIN46(n7771), .CIN45(n7770), .CIN44(n7769), .CIN43(n7768), 
           .CIN42(n7767), .CIN41(n7766), .CIN40(n7765), .CIN39(n7764), 
           .CIN38(n7763), .CIN37(n7762), .CIN36(n7761), .CIN35(n7760), 
           .CIN34(n7759), .CIN33(n7758), .CIN32(n7757), .CIN31(n7756), 
           .CIN30(n7755), .CIN29(n7754), .CIN28(n7753), .CIN27(n7752), 
           .CIN26(n7751), .CIN25(n7750), .CIN24(n7749), .CIN23(n7748), 
           .CIN22(n7747), .CIN21(n7746), .CIN20(n7745), .CIN19(n7744), 
           .CIN18(n7743), .CIN17(n177_adj_1145), .CIN16(n178), .CIN15(n179), 
           .CIN14(n7436), .CIN13(n7437), .CIN12(n7438), .CIN11(n7439), 
           .CIN10(n7440), .CIN9(n7441), .CIN8(n7442), .CIN7(n7443), 
           .CIN6(n7444), .CIN5(n7445), .CIN4(n7446), .CIN3(n7447), .CIN2(n7448), 
           .CIN1(n7449), .CIN0(n7450), .OP10(GND_net), .OP9(VCC_net), 
           .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), 
           .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), 
           .OP0(VCC_net), .R29(n147_adj_1175), .R28(n148_adj_1174), .R27(n149_adj_1173), 
           .R26(n150_adj_1172), .R25(n151_adj_1171), .R24(n152_adj_1170), 
           .R23(n153_adj_1169), .R22(n154_adj_1168), .R21(n155_adj_1167), 
           .R20(n156_adj_1166), .R19(n157_adj_1165), .R18(n158_adj_1164), 
           .R17(n159_adj_1163), .R16(n160_adj_1162), .R15(n161_adj_1161), 
           .R14(n162_adj_1160), .R13(n163_adj_1159), .R12(n164_adj_1158), 
           .R11(n165_adj_1157), .R10(n166_adj_1156), .R9(n167_adj_1155), 
           .R8(n168_adj_1154), .R7(n169_adj_1153), .R6(n170_adj_1152), 
           .R5(n171_adj_1151), .R4(n172_adj_1150), .R3(n173_adj_1149), 
           .R2(n174_adj_1148), .R1(n175_adj_1147), .R0(n176_adj_1146));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam lat_alu_19.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_19.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_19.REG_FLAG_CLK = "NONE";
    defparam lat_alu_19.REG_FLAG_CE = "CE0";
    defparam lat_alu_19.REG_FLAG_RST = "RST0";
    defparam lat_alu_19.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASK01 = "0x00000000000000";
    defparam lat_alu_19.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_19.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_19.CLK0_DIV = "ENABLED";
    defparam lat_alu_19.CLK1_DIV = "ENABLED";
    defparam lat_alu_19.CLK2_DIV = "ENABLED";
    defparam lat_alu_19.CLK3_DIV = "ENABLED";
    defparam lat_alu_19.MCPAT = "0x00000000000000";
    defparam lat_alu_19.MASKPAT = "0x00000000000000";
    defparam lat_alu_19.RNDPAT = "0x00000000000000";
    defparam lat_alu_19.GSR = "DISABLED";
    defparam lat_alu_19.RESETMODE = "SYNC";
    defparam lat_alu_19.MULT9_MODE = "DISABLED";
    defparam lat_alu_19.LEGACY = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i32 (.D(n148_adj_1174), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[46]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i32.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i31 (.D(n149_adj_1173), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i31.GSR = "DISABLED";
    FD1P3AX a_inv_reg_res1_i0_i1 (.D(a_inv_15__N_487[32]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i1.GSR = "ENABLED";
    FD1P3AX prod_d__3_res11_e3__i30 (.D(n150_adj_1172), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[44]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i30.GSR = "DISABLED";
    LUT4 i23_4_lut (.A(det_q4_28_31__N_551[24]), .B(det_q4_28_31__N_551[21]), 
         .C(det_q4_28_31__N_551[11]), .D(det_q4_28_31__N_551[16]), .Z(n55_adj_1297)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i23_4_lut.init = 16'hfffe;
    FD1P3AX prod_d__3_res11_e3__i29 (.D(n151_adj_1171), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i29.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i28 (.D(n152_adj_1170), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[42]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i28.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i27 (.D(n153_adj_1169), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i27.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i26 (.D(n154_adj_1168), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[40]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i26.GSR = "DISABLED";
    FD1P3AX c_inv_reg_res3_i0_i1 (.D(c_inv_15__N_519[32]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(c_inv_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i1.GSR = "ENABLED";
    FD1P3AX det_zero_reg_83 (.D(det_zero_reg_N_907), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_zero_reg));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_zero_reg_83.GSR = "ENABLED";
    LUT4 i16_2_lut (.A(det_q4_28_31__N_551[28]), .B(det_q4_28_31__N_551[12]), 
         .Z(n48_adj_1231)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i16_2_lut.init = 16'heeee;
    FD1S3JX state_FSM_i1 (.D(n7913), .CK(clk_c), .PD(clk_c_enable_348), 
            .Q(n2813));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(det_q4_28_31__N_551[22]), .B(det_q4_28_31__N_551[29]), 
         .Z(n37_adj_1239)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(det_q4_28_31__N_551[13]), .B(det_q4_28_31__N_551[23]), 
         .C(det_q4_28_31__N_551[15]), .D(det_q4_28_31__N_551[20]), .Z(n52_adj_1177)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i20_4_lut.init = 16'hfffe;
    FD1P3AX prod_d__3_res11_e3__i25 (.D(n155_adj_1167), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i25.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i24 (.D(n156_adj_1166), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[38]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i24.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i23 (.D(n157_adj_1165), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i23.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i22 (.D(n158_adj_1164), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[36]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i22.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i21 (.D(n159_adj_1163), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i21.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i20 (.D(n160_adj_1162), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[34]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i20.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i19 (.D(n161_adj_1161), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i19.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i18 (.D(n162_adj_1160), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[32]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i18.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i1 (.D(n179_adj_1178), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i1.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i17 (.D(n163_adj_1159), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[31]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i17.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i1 (.D(d_reg[0]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n130_adj_1211));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i1.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i16 (.D(n164_adj_1158), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[30]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i16.GSR = "DISABLED";
    CCU2C b_s_res8_e3_add_4_17 (.A0(b_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8293), .S0(n41_adj_1241), .S1(n38_adj_1240));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_17.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_17.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_17.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_17.INJECT1_1 = "NO";
    ALU54B lat_alu_3 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n6407), .SIGNEDIB(n6480), .SIGNEDCIN(GND_net), .A35(n6406), 
           .A34(n6405), .A33(n6404), .A32(n6403), .A31(n6402), .A30(n6401), 
           .A29(n6400), .A28(n6399), .A27(n6398), .A26(n6397), .A25(n6396), 
           .A24(n6395), .A23(n6394), .A22(n6393), .A21(n6392), .A20(n6391), 
           .A19(n6390), .A18(n6389), .A17(n6388), .A16(n6387), .A15(n6386), 
           .A14(n6385), .A13(n6384), .A12(n6383), .A11(n6382), .A10(n6381), 
           .A9(n6380), .A8(n6379), .A7(n6378), .A6(n6377), .A5(n6376), 
           .A4(n6375), .A3(n6374), .A2(n6373), .A1(n6372), .A0(n6371), 
           .B35(n6479), .B34(n6478), .B33(n6477), .B32(n6476), .B31(n6475), 
           .B30(n6474), .B29(n6473), .B28(n6472), .B27(n6471), .B26(n6470), 
           .B25(n6469), .B24(n6468), .B23(n6467), .B22(n6466), .B21(n6465), 
           .B20(n6464), .B19(n6463), .B18(n6462), .B17(n6461), .B16(n6460), 
           .B15(n6459), .B14(n6458), .B13(n6457), .B12(n6456), .B11(n6455), 
           .B10(n6454), .B9(n6453), .B8(n6452), .B7(n6451), .B6(n6450), 
           .B5(n6449), .B4(n6448), .B3(n6447), .B2(n6446), .B1(n6445), 
           .B0(n6444), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n6443), .MA34(n6442), .MA33(n6441), .MA32(n6440), .MA31(n6439), 
           .MA30(n6438), .MA29(n6437), .MA28(n6436), .MA27(n6435), .MA26(n6434), 
           .MA25(n6433), .MA24(n6432), .MA23(n6431), .MA22(n6430), .MA21(n6429), 
           .MA20(n6428), .MA19(n6427), .MA18(n6426), .MA17(n6425), .MA16(n6424), 
           .MA15(n6423), .MA14(n6422), .MA13(n6421), .MA12(n6420), .MA11(n6419), 
           .MA10(n6418), .MA9(n6417), .MA8(n6416), .MA7(n6415), .MA6(n6414), 
           .MA5(n6413), .MA4(n6412), .MA3(n6411), .MA2(n6410), .MA1(n6409), 
           .MA0(n6408), .MB35(n6516), .MB34(n6515), .MB33(n6514), .MB32(n6513), 
           .MB31(n6512), .MB30(n6511), .MB29(n6510), .MB28(n6509), .MB27(n6508), 
           .MB26(n6507), .MB25(n6506), .MB24(n6505), .MB23(n6504), .MB22(n6503), 
           .MB21(n6502), .MB20(n6501), .MB19(n6500), .MB18(n6499), .MB17(n6498), 
           .MB16(n6497), .MB15(n6496), .MB14(n6495), .MB13(n6494), .MB12(n6493), 
           .MB11(n6492), .MB10(n6491), .MB9(n6490), .MB8(n6489), .MB7(n6488), 
           .MB6(n6487), .MB5(n6486), .MB4(n6485), .MB3(n6484), .MB2(n6483), 
           .MB1(n6482), .MB0(n6481), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n6698), 
           .R52(n6697), .R51(n6696), .R50(n6695), .R49(n6694), .R48(n6693), 
           .R47(n6692), .R46(n6691), .R45(n6690), .R44(n6689), .R43(n6688), 
           .R42(n6687), .R41(n6686), .R40(n6685), .R39(n6684), .R38(n6683), 
           .R37(n6682), .R36(n6681), .R35(n6680), .R34(n6679), .R33(n6678), 
           .R32(n6677), .R31(n6676), .R30(n6675), .R29(n6674), .R28(n6673), 
           .R27(n6672), .R26(n6671), .R25(n6670), .R24(n6669), .R23(n6668), 
           .R22(n6667), .R21(n6666), .R20(n6665), .R19(n6664), .R18(n6663), 
           .R17(n177_adj_1180), .R16(n178_adj_1179), .R15(n179_adj_1178), 
           .R14(n6356), .R13(n6357), .R12(n6358), .R11(n6359), .R10(n6360), 
           .R9(n6361), .R8(n6362), .R7(n6363), .R6(n6364), .R5(n6365), 
           .R4(n6366), .R3(n6367), .R2(n6368), .R1(n6369), .R0(n6370), 
           .SIGNEDR(n6699));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam lat_alu_3.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_3.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_3.REG_FLAG_CLK = "NONE";
    defparam lat_alu_3.REG_FLAG_CE = "CE0";
    defparam lat_alu_3.REG_FLAG_RST = "RST0";
    defparam lat_alu_3.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASK01 = "0x00000000000000";
    defparam lat_alu_3.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_3.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_3.CLK0_DIV = "ENABLED";
    defparam lat_alu_3.CLK1_DIV = "ENABLED";
    defparam lat_alu_3.CLK2_DIV = "ENABLED";
    defparam lat_alu_3.CLK3_DIV = "ENABLED";
    defparam lat_alu_3.MCPAT = "0x00000000000000";
    defparam lat_alu_3.MASKPAT = "0x00000000000000";
    defparam lat_alu_3.RNDPAT = "0x00000000000000";
    defparam lat_alu_3.GSR = "DISABLED";
    defparam lat_alu_3.RESETMODE = "SYNC";
    defparam lat_alu_3.MULT9_MODE = "DISABLED";
    defparam lat_alu_3.LEGACY = "DISABLED";
    MULT18X18D lat_mult_2 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(n68_adj_1226), .B16(n68_adj_1226), 
            .B15(n68_adj_1226), .B14(n68_adj_1226), .B13(n68_adj_1226), 
            .B12(n68_adj_1226), .B11(n68_adj_1226), .B10(n68_adj_1226), 
            .B9(n68_adj_1226), .B8(n68_adj_1226), .B7(n68_adj_1226), .B6(n68_adj_1226), 
            .B5(n68_adj_1226), .B4(n68_adj_1226), .B3(n68_adj_1226), .B2(n68_adj_1226), 
            .B1(n68_adj_1226), .B0(n68_adj_1226), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n6607), .ROA16(n6606), .ROA15(n6605), .ROA14(n6604), 
            .ROA13(n6603), .ROA12(n6602), .ROA11(n6601), .ROA10(n6600), 
            .ROA9(n6599), .ROA8(n6598), .ROA7(n6597), .ROA6(n6596), 
            .ROA5(n6595), .ROA4(n6594), .ROA3(n6593), .ROA2(n6592), 
            .ROA1(n6591), .ROA0(n6590), .ROB17(n6625), .ROB16(n6624), 
            .ROB15(n6623), .ROB14(n6622), .ROB13(n6621), .ROB12(n6620), 
            .ROB11(n6619), .ROB10(n6618), .ROB9(n6617), .ROB8(n6616), 
            .ROB7(n6615), .ROB6(n6614), .ROB5(n6613), .ROB4(n6612), 
            .ROB3(n6611), .ROB2(n6610), .ROB1(n6609), .ROB0(n6608), 
            .P35(n6662), .P34(n6661), .P33(n6660), .P32(n6659), .P31(n6658), 
            .P30(n6657), .P29(n6656), .P28(n6655), .P27(n6654), .P26(n6653), 
            .P25(n6652), .P24(n6651), .P23(n6650), .P22(n6649), .P21(n6648), 
            .P20(n6647), .P19(n6646), .P18(n6645), .P17(n6644), .P16(n6643), 
            .P15(n6642), .P14(n6641), .P13(n6640), .P12(n6639), .P11(n6638), 
            .P10(n6637), .P9(n6636), .P8(n6635), .P7(n6634), .P6(n6633), 
            .P5(n6632), .P4(n6631), .P3(n6630), .P2(n6629), .P1(n6628), 
            .P0(n6627), .SIGNEDP(n6626));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam lat_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_2.REG_INPUTA_CE = "CE3";
    defparam lat_mult_2.REG_INPUTA_RST = "RST3";
    defparam lat_mult_2.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTB_CE = "CE0";
    defparam lat_mult_2.REG_INPUTB_RST = "RST0";
    defparam lat_mult_2.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTC_CE = "CE0";
    defparam lat_mult_2.REG_INPUTC_RST = "RST0";
    defparam lat_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_2.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_2.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_2.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_2.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_2.CLK0_DIV = "ENABLED";
    defparam lat_mult_2.CLK1_DIV = "ENABLED";
    defparam lat_mult_2.CLK2_DIV = "ENABLED";
    defparam lat_mult_2.CLK3_DIV = "ENABLED";
    defparam lat_mult_2.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_2.GSR = "DISABLED";
    defparam lat_mult_2.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_2.MULT_BYPASS = "DISABLED";
    defparam lat_mult_2.RESETMODE = "ASYNC";
    MULT18X18D prod_c__2_res9_mult_2 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(GND_net), .B16(n5293), .B15(n5294), 
            .B14(n5295), .B13(n5296), .B12(n5297), .B11(n5298), .B10(n5299), 
            .B9(n5300), .B8(n5301), .B7(n5302), .B6(n5303), .B5(n5304), 
            .B4(n5305), .B3(n5306), .B2(n5307), .B1(n5308), .B0(n5373), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n7108), .ROA16(n7107), 
            .ROA15(n7106), .ROA14(n7105), .ROA13(n7104), .ROA12(n7103), 
            .ROA11(n7102), .ROA10(n7101), .ROA9(n7100), .ROA8(n7099), 
            .ROA7(n7098), .ROA6(n7097), .ROA5(n7096), .ROA4(n7095), 
            .ROA3(n7094), .ROA2(n7093), .ROA1(n7092), .ROA0(n7091), 
            .ROB17(n7126), .ROB16(n7125), .ROB15(n7124), .ROB14(n7123), 
            .ROB13(n7122), .ROB12(n7121), .ROB11(n7120), .ROB10(n7119), 
            .ROB9(n7118), .ROB8(n7117), .ROB7(n7116), .ROB6(n7115), 
            .ROB5(n7114), .ROB4(n7113), .ROB3(n7112), .ROB2(n7111), 
            .ROB1(n7110), .ROB0(n7109), .P35(n7163), .P34(n7162), .P33(n7161), 
            .P32(n7160), .P31(n7159), .P30(n7158), .P29(n7157), .P28(n7156), 
            .P27(n7155), .P26(n7154), .P25(n7153), .P24(n7152), .P23(n7151), 
            .P22(n7150), .P21(n7149), .P20(n7148), .P19(n7147), .P18(n7146), 
            .P17(n7145), .P16(n7144), .P15(n7143), .P14(n7142), .P13(n7141), 
            .P12(n7140), .P11(n7139), .P10(n7138), .P9(n7137), .P8(n7136), 
            .P7(n7135), .P6(n7134), .P5(n7133), .P4(n7132), .P3(n7131), 
            .P2(n7130), .P1(n7129), .P0(n7128), .SIGNEDP(n7127));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam prod_c__2_res9_mult_2.REG_INPUTA_CE = "CE3";
    defparam prod_c__2_res9_mult_2.REG_INPUTA_RST = "RST3";
    defparam prod_c__2_res9_mult_2.REG_INPUTB_CLK = "NONE";
    defparam prod_c__2_res9_mult_2.REG_INPUTB_CE = "CE0";
    defparam prod_c__2_res9_mult_2.REG_INPUTB_RST = "RST0";
    defparam prod_c__2_res9_mult_2.REG_INPUTC_CLK = "NONE";
    defparam prod_c__2_res9_mult_2.REG_INPUTC_CE = "CE0";
    defparam prod_c__2_res9_mult_2.REG_INPUTC_RST = "RST0";
    defparam prod_c__2_res9_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam prod_c__2_res9_mult_2.REG_PIPELINE_CE = "CE0";
    defparam prod_c__2_res9_mult_2.REG_PIPELINE_RST = "RST0";
    defparam prod_c__2_res9_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam prod_c__2_res9_mult_2.REG_OUTPUT_CE = "CE0";
    defparam prod_c__2_res9_mult_2.REG_OUTPUT_RST = "RST0";
    defparam prod_c__2_res9_mult_2.CLK0_DIV = "ENABLED";
    defparam prod_c__2_res9_mult_2.CLK1_DIV = "ENABLED";
    defparam prod_c__2_res9_mult_2.CLK2_DIV = "ENABLED";
    defparam prod_c__2_res9_mult_2.CLK3_DIV = "ENABLED";
    defparam prod_c__2_res9_mult_2.HIGHSPEED_CLK = "NONE";
    defparam prod_c__2_res9_mult_2.GSR = "DISABLED";
    defparam prod_c__2_res9_mult_2.CAS_MATCH_REG = "FALSE";
    defparam prod_c__2_res9_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam prod_c__2_res9_mult_2.MULT_BYPASS = "DISABLED";
    defparam prod_c__2_res9_mult_2.RESETMODE = "ASYNC";
    FD1P3AX prod_d__3_res11_e3__i15 (.D(n165_adj_1157), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[29]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i15.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i14 (.D(n166_adj_1156), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[28]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i14.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i13 (.D(n167_adj_1155), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[27]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i13.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i12 (.D(n168_adj_1154), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[26]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i12.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i11 (.D(n169_adj_1153), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[25]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i11.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i10 (.D(n170_adj_1152), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[24]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i10.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i9 (.D(n171_adj_1151), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[23]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i9.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i8 (.D(n172_adj_1150), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[22]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i8.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i7 (.D(n173_adj_1149), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[21]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i7.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i6 (.D(n174_adj_1148), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[20]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i6.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i5 (.D(n175_adj_1147), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[19]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i5.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i4 (.D(n176_adj_1146), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[18]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i4.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i3 (.D(n177_adj_1145), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_d[17]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i3.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i2 (.D(n178), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_d[16]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i2.GSR = "DISABLED";
    LUT4 i272_1_lut_rep_19 (.A(reset_c), .Z(n8725)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(3[35:40])
    defparam i272_1_lut_rep_19.init = 16'h5555;
    LUT4 i574_2_lut (.A(n2813), .B(next_state_2__N_68_c_0), .Z(n7913)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam i574_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_3_lut (.A(reset_c), .B(n3861), .C(clk_c_enable_239), 
         .Z(clk_c_enable_432)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(3[35:40])
    defparam i1_3_lut_3_lut.init = 16'h5454;
    FD1P3AX a_reg_i0_i0 (.D(a_c_0), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(a_reg[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i0.GSR = "ENABLED";
    MULT18X18D lat_mult_1 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(n68_adj_1226), .B16(n68_adj_1226), 
            .B15(n68_adj_1226), .B14(n68_adj_1226), .B13(n68_adj_1226), 
            .B12(n68_adj_1226), .B11(n68_adj_1226), .B10(n68_adj_1226), 
            .B9(n68_adj_1226), .B8(n68_adj_1226), .B7(n68_adj_1226), .B6(n68_adj_1226), 
            .B5(n68_adj_1226), .B4(n68_adj_1226), .B3(n68_adj_1226), .B2(n68_adj_1226), 
            .B1(n68_adj_1226), .B0(n68_adj_1226), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n6534), .ROA16(n6533), .ROA15(n6532), .ROA14(n6531), 
            .ROA13(n6530), .ROA12(n6529), .ROA11(n6528), .ROA10(n6527), 
            .ROA9(n6526), .ROA8(n6525), .ROA7(n6524), .ROA6(n6523), 
            .ROA5(n6522), .ROA4(n6521), .ROA3(n6520), .ROA2(n6519), 
            .ROA1(n6518), .ROA0(n6517), .ROB17(n6552), .ROB16(n6551), 
            .ROB15(n6550), .ROB14(n6549), .ROB13(n6548), .ROB12(n6547), 
            .ROB11(n6546), .ROB10(n6545), .ROB9(n6544), .ROB8(n6543), 
            .ROB7(n6542), .ROB6(n6541), .ROB5(n6540), .ROB4(n6539), 
            .ROB3(n6538), .ROB2(n6537), .ROB1(n6536), .ROB0(n6535), 
            .P35(n6589), .P34(n6588), .P33(n6587), .P32(n6586), .P31(n6585), 
            .P30(n6584), .P29(n6583), .P28(n6582), .P27(n6581), .P26(n6580), 
            .P25(n6579), .P24(n6578), .P23(n6577), .P22(n6576), .P21(n6575), 
            .P20(n6574), .P19(n6573), .P18(n6572), .P17(n6571), .P16(n6570), 
            .P15(n6569), .P14(n6568), .P13(n6567), .P12(n6566), .P11(n6565), 
            .P10(n6564), .P9(n6563), .P8(n6562), .P7(n6561), .P6(n6560), 
            .P5(n6559), .P4(n6558), .P3(n6557), .P2(n6556), .P1(n6555), 
            .P0(n6554), .SIGNEDP(n6553));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam lat_mult_1.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_1.REG_INPUTA_CE = "CE3";
    defparam lat_mult_1.REG_INPUTA_RST = "RST3";
    defparam lat_mult_1.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTB_CE = "CE0";
    defparam lat_mult_1.REG_INPUTB_RST = "RST0";
    defparam lat_mult_1.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTC_CE = "CE0";
    defparam lat_mult_1.REG_INPUTC_RST = "RST0";
    defparam lat_mult_1.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_1.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_1.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_1.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_1.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_1.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_1.CLK0_DIV = "ENABLED";
    defparam lat_mult_1.CLK1_DIV = "ENABLED";
    defparam lat_mult_1.CLK2_DIV = "ENABLED";
    defparam lat_mult_1.CLK3_DIV = "ENABLED";
    defparam lat_mult_1.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_1.GSR = "DISABLED";
    defparam lat_mult_1.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_1.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_1.MULT_BYPASS = "DISABLED";
    defparam lat_mult_1.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_0 (.A17(quotient_31__N_908[31]), .A16(quotient_31__N_908[31]), 
            .A15(quotient_31__N_908[31]), .A14(quotient_31__N_908[31]), 
            .A13(quotient_31__N_908[31]), .A12(quotient_31__N_908[30]), 
            .A11(quotient_31__N_908[29]), .A10(quotient_31__N_908[28]), 
            .A9(quotient_31__N_908[27]), .A8(quotient_31__N_908[26]), .A7(quotient_31__N_908[25]), 
            .A6(quotient_31__N_908[24]), .A5(quotient_31__N_908[23]), .A4(quotient_31__N_908[22]), 
            .A3(quotient_31__N_908[21]), .A2(quotient_31__N_908[20]), .A1(quotient_31__N_908[19]), 
            .A0(quotient_31__N_908[18]), .B17(n68_adj_1226), .B16(n68_adj_1226), 
            .B15(n68_adj_1226), .B14(n102_adj_1225), .B13(n104_adj_1224), 
            .B12(n106_adj_1223), .B11(n108_adj_1222), .B10(n110_adj_1221), 
            .B9(n112_adj_1220), .B8(n114_adj_1219), .B7(n116_adj_1218), 
            .B6(n118_adj_1217), .B5(n120_adj_1216), .B4(n122_adj_1215), 
            .B3(n124_adj_1214), .B2(n126_adj_1213), .B1(n128_adj_1212), 
            .B0(n130_adj_1211), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n6461), 
            .ROA16(n6460), .ROA15(n6459), .ROA14(n6458), .ROA13(n6457), 
            .ROA12(n6456), .ROA11(n6455), .ROA10(n6454), .ROA9(n6453), 
            .ROA8(n6452), .ROA7(n6451), .ROA6(n6450), .ROA5(n6449), 
            .ROA4(n6448), .ROA3(n6447), .ROA2(n6446), .ROA1(n6445), 
            .ROA0(n6444), .ROB17(n6479), .ROB16(n6478), .ROB15(n6477), 
            .ROB14(n6476), .ROB13(n6475), .ROB12(n6474), .ROB11(n6473), 
            .ROB10(n6472), .ROB9(n6471), .ROB8(n6470), .ROB7(n6469), 
            .ROB6(n6468), .ROB5(n6467), .ROB4(n6466), .ROB3(n6465), 
            .ROB2(n6464), .ROB1(n6463), .ROB0(n6462), .P35(n6516), .P34(n6515), 
            .P33(n6514), .P32(n6513), .P31(n6512), .P30(n6511), .P29(n6510), 
            .P28(n6509), .P27(n6508), .P26(n6507), .P25(n6506), .P24(n6505), 
            .P23(n6504), .P22(n6503), .P21(n6502), .P20(n6501), .P19(n6500), 
            .P18(n6499), .P17(n6498), .P16(n6497), .P15(n6496), .P14(n6495), 
            .P13(n6494), .P12(n6493), .P11(n6492), .P10(n6491), .P9(n6490), 
            .P8(n6489), .P7(n6488), .P6(n6487), .P5(n6486), .P4(n6485), 
            .P3(n6484), .P2(n6483), .P1(n6482), .P0(n6481), .SIGNEDP(n6480));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam lat_mult_0.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_0.REG_INPUTA_CE = "CE3";
    defparam lat_mult_0.REG_INPUTA_RST = "RST3";
    defparam lat_mult_0.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTB_CE = "CE0";
    defparam lat_mult_0.REG_INPUTB_RST = "RST0";
    defparam lat_mult_0.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTC_CE = "CE0";
    defparam lat_mult_0.REG_INPUTC_RST = "RST0";
    defparam lat_mult_0.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_0.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_0.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_0.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_0.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_0.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_0.CLK0_DIV = "ENABLED";
    defparam lat_mult_0.CLK1_DIV = "ENABLED";
    defparam lat_mult_0.CLK2_DIV = "ENABLED";
    defparam lat_mult_0.CLK3_DIV = "ENABLED";
    defparam lat_mult_0.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_0.GSR = "DISABLED";
    defparam lat_mult_0.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_0.MULT_BYPASS = "DISABLED";
    defparam lat_mult_0.RESETMODE = "ASYNC";
    MULT18X18D prod_a__0_res5_mult_2 (.A17(quotient_31__N_908[17]), .A16(quotient_31__N_908[16]), 
            .A15(quotient_31__N_908[15]), .A14(quotient_31__N_908[14]), 
            .A13(quotient_31__N_908[13]), .A12(quotient_31__N_908[12]), 
            .A11(quotient_31__N_908[11]), .A10(quotient_31__N_908[10]), 
            .A9(quotient_31__N_908[9]), .A8(quotient_31__N_908[8]), .A7(quotient_31__N_908[7]), 
            .A6(quotient_31__N_908[6]), .A5(quotient_31__N_908[5]), .A4(quotient_31__N_908[4]), 
            .A3(quotient_31__N_908[3]), .A2(quotient_31__N_908[2]), .A1(quotient_31__N_908[1]), 
            .A0(quotient_31__N_908[0]), .B17(n68_adj_1226), .B16(n68_adj_1226), 
            .B15(n68_adj_1226), .B14(n102_adj_1225), .B13(n104_adj_1224), 
            .B12(n106_adj_1223), .B11(n108_adj_1222), .B10(n110_adj_1221), 
            .B9(n112_adj_1220), .B8(n114_adj_1219), .B7(n116_adj_1218), 
            .B6(n118_adj_1217), .B5(n120_adj_1216), .B4(n122_adj_1215), 
            .B3(n124_adj_1214), .B2(n126_adj_1213), .B1(n128_adj_1212), 
            .B0(n130_adj_1211), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n6388), 
            .ROA16(n6387), .ROA15(n6386), .ROA14(n6385), .ROA13(n6384), 
            .ROA12(n6383), .ROA11(n6382), .ROA10(n6381), .ROA9(n6380), 
            .ROA8(n6379), .ROA7(n6378), .ROA6(n6377), .ROA5(n6376), 
            .ROA4(n6375), .ROA3(n6374), .ROA2(n6373), .ROA1(n6372), 
            .ROA0(n6371), .ROB17(n6406), .ROB16(n6405), .ROB15(n6404), 
            .ROB14(n6403), .ROB13(n6402), .ROB12(n6401), .ROB11(n6400), 
            .ROB10(n6399), .ROB9(n6398), .ROB8(n6397), .ROB7(n6396), 
            .ROB6(n6395), .ROB5(n6394), .ROB4(n6393), .ROB3(n6392), 
            .ROB2(n6391), .ROB1(n6390), .ROB0(n6389), .P35(n6443), .P34(n6442), 
            .P33(n6441), .P32(n6440), .P31(n6439), .P30(n6438), .P29(n6437), 
            .P28(n6436), .P27(n6435), .P26(n6434), .P25(n6433), .P24(n6432), 
            .P23(n6431), .P22(n6430), .P21(n6429), .P20(n6428), .P19(n6427), 
            .P18(n6426), .P17(n6425), .P16(n6424), .P15(n6423), .P14(n6422), 
            .P13(n6421), .P12(n6420), .P11(n6419), .P10(n6418), .P9(n6417), 
            .P8(n6416), .P7(n6415), .P6(n6414), .P5(n6413), .P4(n6412), 
            .P3(n6411), .P2(n6410), .P1(n6409), .P0(n6408), .SIGNEDP(n6407));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam prod_a__0_res5_mult_2.REG_INPUTA_CE = "CE3";
    defparam prod_a__0_res5_mult_2.REG_INPUTA_RST = "RST3";
    defparam prod_a__0_res5_mult_2.REG_INPUTB_CLK = "NONE";
    defparam prod_a__0_res5_mult_2.REG_INPUTB_CE = "CE0";
    defparam prod_a__0_res5_mult_2.REG_INPUTB_RST = "RST0";
    defparam prod_a__0_res5_mult_2.REG_INPUTC_CLK = "NONE";
    defparam prod_a__0_res5_mult_2.REG_INPUTC_CE = "CE0";
    defparam prod_a__0_res5_mult_2.REG_INPUTC_RST = "RST0";
    defparam prod_a__0_res5_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam prod_a__0_res5_mult_2.REG_PIPELINE_CE = "CE0";
    defparam prod_a__0_res5_mult_2.REG_PIPELINE_RST = "RST0";
    defparam prod_a__0_res5_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam prod_a__0_res5_mult_2.REG_OUTPUT_CE = "CE0";
    defparam prod_a__0_res5_mult_2.REG_OUTPUT_RST = "RST0";
    defparam prod_a__0_res5_mult_2.CLK0_DIV = "ENABLED";
    defparam prod_a__0_res5_mult_2.CLK1_DIV = "ENABLED";
    defparam prod_a__0_res5_mult_2.CLK2_DIV = "ENABLED";
    defparam prod_a__0_res5_mult_2.CLK3_DIV = "ENABLED";
    defparam prod_a__0_res5_mult_2.HIGHSPEED_CLK = "NONE";
    defparam prod_a__0_res5_mult_2.GSR = "DISABLED";
    defparam prod_a__0_res5_mult_2.CAS_MATCH_REG = "FALSE";
    defparam prod_a__0_res5_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam prod_a__0_res5_mult_2.MULT_BYPASS = "DISABLED";
    defparam prod_a__0_res5_mult_2.RESETMODE = "ASYNC";
    FD1P3AX c_s_res10_e3_e3__i1 (.D(n86_adj_1273), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5373));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i1.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n8725));
    CCU2C b_s_res8_e3_add_4_15 (.A0(b_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8292), .COUT(n8293), .S0(n47_adj_1243), 
          .S1(n44_adj_1242));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_15.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_15.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_15.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_15.INJECT1_1 = "NO";
    FD1P3AX c_s_res10_e3_e3__i17 (.D(n38_adj_1257), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5293));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i17.GSR = "DISABLED";
    OB a_inv_pad_14 (.I(a_inv_c_14), .O(a_inv[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    FD1P3AX c_s_res10_e3_e3__i16 (.D(n41_adj_1258), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5294));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i16.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i15 (.D(n44_adj_1259), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5295));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i15.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i14 (.D(n47_adj_1260), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5296));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i14.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i13 (.D(n50_adj_1261), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5297));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i13.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i12 (.D(n53_adj_1262), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5298));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i12.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i11 (.D(n56_adj_1263), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5299));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i11.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i10 (.D(n59_adj_1264), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5300));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i10.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i9 (.D(n62_adj_1265), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5301));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i9.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i8 (.D(n65_adj_1266), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5302));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i8.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i7 (.D(n68_adj_1267), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5303));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i7.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i6 (.D(n71_adj_1268), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5304));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i6.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i5 (.D(n74_adj_1269), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5305));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i5.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i4 (.D(n77_adj_1270), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5306));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i4.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i3 (.D(n80_adj_1271), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5307));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i3.GSR = "DISABLED";
    FD1P3AX c_s_res10_e3_e3__i2 (.D(n83_adj_1272), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5308));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_e3__i2.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e3__i1 (.D(n179), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_d[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e3__i1.GSR = "DISABLED";
    FD1P3AX b_reg_i0_i1 (.D(b_c_1), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i1.GSR = "ENABLED";
    LUT4 i145_2_lut (.A(next_state_2__N_68_c_0), .B(n2813), .Z(n2820)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam i145_2_lut.init = 16'h8888;
    OB a_inv_pad_13 (.I(a_inv_c_13), .O(a_inv[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_12 (.I(a_inv_c_12), .O(a_inv[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_11 (.I(a_inv_c_11), .O(a_inv[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_10 (.I(a_inv_c_10), .O(a_inv[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_9 (.I(a_inv_c_9), .O(a_inv[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_8 (.I(a_inv_c_8), .O(a_inv[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_7 (.I(a_inv_c_7), .O(a_inv[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_6 (.I(a_inv_c_6), .O(a_inv[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_5 (.I(a_inv_c_5), .O(a_inv[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_4 (.I(a_inv_c_4), .O(a_inv[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_3 (.I(a_inv_c_3), .O(a_inv[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_2 (.I(a_inv_c_2), .O(a_inv[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_1 (.I(a_inv_c_1), .O(a_inv[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB a_inv_pad_0 (.I(a_inv_c_0), .O(a_inv[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[36:41])
    OB b_inv_pad_15 (.I(b_inv_c_15), .O(b_inv[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_14 (.I(b_inv_c_14), .O(b_inv[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_13 (.I(b_inv_c_13), .O(b_inv[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_12 (.I(b_inv_c_12), .O(b_inv[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_11 (.I(b_inv_c_11), .O(b_inv[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_10 (.I(b_inv_c_10), .O(b_inv[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_9 (.I(b_inv_c_9), .O(b_inv[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_8 (.I(b_inv_c_8), .O(b_inv[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_7 (.I(b_inv_c_7), .O(b_inv[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_6 (.I(b_inv_c_6), .O(b_inv[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_5 (.I(b_inv_c_5), .O(b_inv[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_4 (.I(b_inv_c_4), .O(b_inv[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_3 (.I(b_inv_c_3), .O(b_inv[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_2 (.I(b_inv_c_2), .O(b_inv[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_1 (.I(b_inv_c_1), .O(b_inv[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB b_inv_pad_0 (.I(b_inv_c_0), .O(b_inv[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[43:48])
    OB c_inv_pad_15 (.I(c_inv_c_15), .O(c_inv[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_14 (.I(c_inv_c_14), .O(c_inv[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_13 (.I(c_inv_c_13), .O(c_inv[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_12 (.I(c_inv_c_12), .O(c_inv[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_11 (.I(c_inv_c_11), .O(c_inv[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_10 (.I(c_inv_c_10), .O(c_inv[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_9 (.I(c_inv_c_9), .O(c_inv[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_8 (.I(c_inv_c_8), .O(c_inv[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_7 (.I(c_inv_c_7), .O(c_inv[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_6 (.I(c_inv_c_6), .O(c_inv[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_5 (.I(c_inv_c_5), .O(c_inv[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_4 (.I(c_inv_c_4), .O(c_inv[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_3 (.I(c_inv_c_3), .O(c_inv[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_2 (.I(c_inv_c_2), .O(c_inv[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_1 (.I(c_inv_c_1), .O(c_inv[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB c_inv_pad_0 (.I(c_inv_c_0), .O(c_inv[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[50:55])
    OB d_inv_pad_15 (.I(d_inv_c_15), .O(d_inv[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_14 (.I(d_inv_c_14), .O(d_inv[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_13 (.I(d_inv_c_13), .O(d_inv[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_12 (.I(d_inv_c_12), .O(d_inv[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_11 (.I(d_inv_c_11), .O(d_inv[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_10 (.I(d_inv_c_10), .O(d_inv[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_9 (.I(d_inv_c_9), .O(d_inv[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_8 (.I(d_inv_c_8), .O(d_inv[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_7 (.I(d_inv_c_7), .O(d_inv[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_6 (.I(d_inv_c_6), .O(d_inv[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_5 (.I(d_inv_c_5), .O(d_inv[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_4 (.I(d_inv_c_4), .O(d_inv[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_3 (.I(d_inv_c_3), .O(d_inv[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_2 (.I(d_inv_c_2), .O(d_inv[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_1 (.I(d_inv_c_1), .O(d_inv[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB d_inv_pad_0 (.I(d_inv_c_0), .O(d_inv[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(6[57:62])
    OB error_pad (.I(GND_net), .O(error));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(7[36:41])
    OB ready_pad (.I(GND_net), .O(ready));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(8[36:41])
    IB clk_pad (.I(clk), .O(clk_c));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(2[35:38])
    IB reset_pad (.I(reset), .O(reset_c));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(3[35:40])
    IB next_state_2__N_68_pad_0 (.I(start), .O(next_state_2__N_68_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(4[35:40])
    IB a_pad_15 (.I(a[15]), .O(a_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_14 (.I(a[14]), .O(a_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_13 (.I(a[13]), .O(a_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_12 (.I(a[12]), .O(a_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_11 (.I(a[11]), .O(a_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_10 (.I(a[10]), .O(a_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_9 (.I(a[9]), .O(a_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_8 (.I(a[8]), .O(a_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_7 (.I(a[7]), .O(a_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_6 (.I(a[6]), .O(a_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_5 (.I(a[5]), .O(a_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_4 (.I(a[4]), .O(a_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_3 (.I(a[3]), .O(a_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_2 (.I(a[2]), .O(a_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_1 (.I(a[1]), .O(a_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB a_pad_0 (.I(a[0]), .O(a_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[36:37])
    IB b_pad_15 (.I(b[15]), .O(b_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_14 (.I(b[14]), .O(b_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_13 (.I(b[13]), .O(b_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_12 (.I(b[12]), .O(b_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_11 (.I(b[11]), .O(b_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_10 (.I(b[10]), .O(b_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_9 (.I(b[9]), .O(b_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_8 (.I(b[8]), .O(b_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_7 (.I(b[7]), .O(b_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_6 (.I(b[6]), .O(b_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_5 (.I(b[5]), .O(b_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_4 (.I(b[4]), .O(b_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_3 (.I(b[3]), .O(b_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_2 (.I(b[2]), .O(b_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_1 (.I(b[1]), .O(b_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB b_pad_0 (.I(b[0]), .O(b_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[39:40])
    IB c_pad_15 (.I(c[15]), .O(c_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_14 (.I(c[14]), .O(c_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_13 (.I(c[13]), .O(c_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_12 (.I(c[12]), .O(c_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_11 (.I(c[11]), .O(c_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_10 (.I(c[10]), .O(c_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_9 (.I(c[9]), .O(c_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_8 (.I(c[8]), .O(c_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_7 (.I(c[7]), .O(c_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_6 (.I(c[6]), .O(c_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_5 (.I(c[5]), .O(c_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_4 (.I(c[4]), .O(c_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_3 (.I(c[3]), .O(c_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_2 (.I(c[2]), .O(c_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_1 (.I(c[1]), .O(c_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB c_pad_0 (.I(c[0]), .O(c_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[42:43])
    IB d_pad_15 (.I(d[15]), .O(d_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_14 (.I(d[14]), .O(d_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_13 (.I(d[13]), .O(d_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_12 (.I(d[12]), .O(d_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_11 (.I(d[11]), .O(d_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_10 (.I(d[10]), .O(d_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_9 (.I(d[9]), .O(d_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_8 (.I(d[8]), .O(d_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_7 (.I(d[7]), .O(d_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_6 (.I(d[6]), .O(d_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_5 (.I(d[5]), .O(d_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_4 (.I(d[4]), .O(d_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_3 (.I(d[3]), .O(d_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_2 (.I(d[2]), .O(d_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_1 (.I(d[1]), .O(d_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    IB d_pad_0 (.I(d[0]), .O(d_c_0));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(5[45:46])
    LUT4 i577_3_lut (.A(n2810), .B(clk_c_enable_145), .C(next_state_2__N_65[2]), 
         .Z(n7916)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam i577_3_lut.init = 16'hcece;
    LUT4 i693_1_lut (.A(n2810), .Z(n8032)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam i693_1_lut.init = 16'h5555;
    FD1P3AX b_reg_i0_i2 (.D(b_c_2), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i3 (.D(b_c_3), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i3.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i4 (.D(b_c_4), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i4.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i5 (.D(b_c_5), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i5.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i6 (.D(b_c_6), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i6.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i7 (.D(b_c_7), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i7.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i8 (.D(b_c_8), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i8.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i9 (.D(b_c_9), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i9.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i10 (.D(b_c_10), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i10.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i11 (.D(b_c_11), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i11.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i12 (.D(b_c_12), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i12.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i13 (.D(b_c_13), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i13.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i14 (.D(b_c_14), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i14.GSR = "ENABLED";
    FD1P3AX b_reg_i0_i15 (.D(b_c_15), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(b_reg[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_reg_i0_i15.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i1 (.D(c_c_1), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i1.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i2 (.D(c_c_2), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i3 (.D(c_c_3), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i3.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i4 (.D(c_c_4), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i4.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i5 (.D(c_c_5), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i5.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i6 (.D(c_c_6), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i6.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i7 (.D(c_c_7), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i7.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i8 (.D(c_c_8), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i8.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i9 (.D(c_c_9), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i9.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i10 (.D(c_c_10), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i10.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i11 (.D(c_c_11), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i11.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i12 (.D(c_c_12), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i12.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i13 (.D(c_c_13), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i13.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i14 (.D(c_c_14), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i14.GSR = "ENABLED";
    FD1P3AX c_reg_i0_i15 (.D(c_c_15), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(c_reg[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_reg_i0_i15.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i1 (.D(d_c_1), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i1.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i2 (.D(d_c_2), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i3 (.D(d_c_3), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i3.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i4 (.D(d_c_4), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i4.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i5 (.D(d_c_5), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i5.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i6 (.D(d_c_6), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i6.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i7 (.D(d_c_7), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i7.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i8 (.D(d_c_8), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i8.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i9 (.D(d_c_9), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i9.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i10 (.D(d_c_10), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i10.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i11 (.D(d_c_11), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i11.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i12 (.D(d_c_12), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i12.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i13 (.D(d_c_13), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i13.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i14 (.D(d_c_14), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i14.GSR = "ENABLED";
    FD1P3AX d_reg_i0_i15 (.D(d_c_15), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(d_reg[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_reg_i0_i15.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i1 (.D(det_q4_28_31__N_551[1]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i1.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i2 (.D(det_q4_28_31__N_551[2]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i2.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i3 (.D(det_q4_28_31__N_551[3]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i3.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i4 (.D(det_q4_28_31__N_551[4]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i4.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i5 (.D(det_q4_28_31__N_551[5]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i5.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i6 (.D(det_q4_28_31__N_551[6]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i6.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i7 (.D(det_q4_28_31__N_551[7]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i7.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i8 (.D(det_q4_28_31__N_551[8]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i8.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i9 (.D(det_q4_28_31__N_551[9]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i9.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i10 (.D(det_q4_28_31__N_551[10]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i10.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i11 (.D(det_q4_28_31__N_551[11]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i11.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i12 (.D(det_q4_28_31__N_551[12]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i12.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i13 (.D(det_q4_28_31__N_551[13]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i13.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i14 (.D(det_q4_28_31__N_551[14]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i14.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i15 (.D(det_q4_28_31__N_551[15]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i15.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i16 (.D(det_q4_28_31__N_551[16]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[16]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i16.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i17 (.D(det_q4_28_31__N_551[17]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[17]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i17.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i18 (.D(det_q4_28_31__N_551[18]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[18]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i18.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i19 (.D(det_q4_28_31__N_551[19]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[19]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i19.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i20 (.D(det_q4_28_31__N_551[20]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[20]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i20.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i21 (.D(det_q4_28_31__N_551[21]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[21]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i21.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i22 (.D(det_q4_28_31__N_551[22]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[22]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i22.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i23 (.D(det_q4_28_31__N_551[23]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[23]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i23.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i24 (.D(det_q4_28_31__N_551[24]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[24]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i24.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i25 (.D(det_q4_28_31__N_551[25]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[25]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i25.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i26 (.D(det_q4_28_31__N_551[26]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[26]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i26.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i27 (.D(det_q4_28_31__N_551[27]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[27]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i27.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i28 (.D(det_q4_28_31__N_551[28]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[28]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i28.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i29 (.D(det_q4_28_31__N_551[29]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[29]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i29.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i30 (.D(det_q4_28_31__N_551[30]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[30]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i30.GSR = "ENABLED";
    FD1P3AX det_q4_28_i0_i31 (.D(det_q4_28_31__N_551[31]), .SP(clk_c_enable_145), 
            .CK(clk_c), .Q(det_q4_28[31]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam det_q4_28_i0_i31.GSR = "ENABLED";
    FD1P3AX prod_d__3_res11_e2__i2 (.D(a_reg[1]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n128));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i2.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i3 (.D(a_reg[2]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n126));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i3.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i4 (.D(a_reg[3]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n124));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i4.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i5 (.D(a_reg[4]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n122));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i5.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i6 (.D(a_reg[5]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n120));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i6.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i7 (.D(a_reg[6]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n118));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i7.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i8 (.D(a_reg[7]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n116));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i8.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i9 (.D(a_reg[8]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n114));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i9.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i10 (.D(a_reg[9]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n112));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i10.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i11 (.D(a_reg[10]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n110));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i11.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i12 (.D(a_reg[11]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n108));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i12.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i13 (.D(a_reg[12]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n106));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i13.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i14 (.D(a_reg[13]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n104));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i14.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i15 (.D(a_reg[14]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n102));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i15.GSR = "DISABLED";
    FD1P3AX prod_d__3_res11_e2__i16 (.D(a_reg[15]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n68_adj_1176));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(106[31:44])
    defparam prod_d__3_res11_e2__i16.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i2 (.D(n83_adj_1255), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5212));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i2.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i3 (.D(n80_adj_1254), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5211));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i3.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i4 (.D(n77_adj_1253), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5210));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i4.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i5 (.D(n74_adj_1252), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5209));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i5.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i6 (.D(n71_adj_1251), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5208));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i6.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i7 (.D(n68_adj_1250), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5207));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i7.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i8 (.D(n65_adj_1249), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5206));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i8.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i9 (.D(n62_adj_1248), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5205));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i9.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i10 (.D(n59_adj_1247), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5204));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i10.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i11 (.D(n56_adj_1246), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5203));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i11.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i12 (.D(n53_adj_1245), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5202));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i12.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i13 (.D(n50_adj_1244), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5201));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i13.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i14 (.D(n47_adj_1243), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5200));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i14.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i15 (.D(n44_adj_1242), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5199));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i15.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i16 (.D(n41_adj_1241), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5198));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i16.GSR = "DISABLED";
    FD1P3AX b_s_res8_e3_e3__i17 (.D(n38_adj_1240), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n5197));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_e3__i17.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i2 (.D(n178_adj_1228), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_c[16]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i2.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i3 (.D(n177_adj_1232), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_c[17]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i3.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i4 (.D(n176_adj_1233), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_c[18]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i4.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i5 (.D(n175_adj_1234), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_c[19]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i5.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i6 (.D(n174_adj_1235), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_c[20]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i6.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i7 (.D(n173), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[21]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i7.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i8 (.D(n172), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[22]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i8.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i9 (.D(n171), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[23]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i9.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i10 (.D(n170), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[24]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i10.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i11 (.D(n169), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[25]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i11.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i12 (.D(n168), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[26]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i12.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i13 (.D(n167), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[27]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i13.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i14 (.D(n166), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[28]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i14.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i15 (.D(n165), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[29]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i15.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i16 (.D(n164), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[30]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i16.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i17 (.D(n163), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[31]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i17.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i18 (.D(n162), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[32]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i18.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i19 (.D(n161), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i19.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i20 (.D(n160), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[34]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i20.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i21 (.D(n159), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i21.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i22 (.D(n158), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[36]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i22.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i23 (.D(n157), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i23.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i24 (.D(n156), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[38]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i24.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i25 (.D(n155), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i25.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i26 (.D(n154), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[40]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i26.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i27 (.D(n153), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i27.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i28 (.D(n152), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[42]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i28.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i29 (.D(n151), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i29.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i30 (.D(n150), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[44]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i30.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i31 (.D(n149), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i31.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i32 (.D(n148), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[46]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i32.GSR = "DISABLED";
    FD1P3AX prod_c__2_res9_e3__i33 (.D(n147), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_c[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(105[31:44])
    defparam prod_c__2_res9_e3__i33.GSR = "DISABLED";
    FD1P3AX d_inv_reg_res2_i0_i2 (.D(d_inv_15__N_535[33]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i2.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i3 (.D(d_inv_15__N_535[34]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i3.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i4 (.D(d_inv_15__N_535[35]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i4.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i5 (.D(d_inv_15__N_535[36]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i5.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i6 (.D(d_inv_15__N_535[37]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i6.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i7 (.D(d_inv_15__N_535[38]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i7.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i8 (.D(d_inv_15__N_535[39]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i8.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i9 (.D(d_inv_15__N_535[40]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i9.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i10 (.D(d_inv_15__N_535[41]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i10.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i11 (.D(d_inv_15__N_535[42]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i11.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i12 (.D(d_inv_15__N_535[43]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i12.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i13 (.D(d_inv_15__N_535[44]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i13.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i14 (.D(d_inv_15__N_535[45]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i14.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i15 (.D(d_inv_15__N_535[46]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i15.GSR = "ENABLED";
    FD1P3AX d_inv_reg_res2_i0_i16 (.D(d_inv_15__N_535[47]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(d_inv_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam d_inv_reg_res2_i0_i16.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i2 (.D(b_inv_15__N_503[33]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i2.GSR = "ENABLED";
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    divNRDA_FSM u_recip (.regA({regA}), .n4577({n4578, n4579, n4580, 
            n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, 
            n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
            n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, 
            n4605, n4606, n4607, n4608, n4609, n4610}), .clk_c(clk_c), 
            .n168(n168_adj_1296), .clk_c_enable_239(clk_c_enable_239), .det_q4_28({det_q4_28}), 
            .quotient_31__N_908({quotient_31__N_908}), .n3859(n3859), .n3860(n3860), 
            .n7851(n7851), .\next_state_2__N_65[2] (next_state_2__N_65[2]), 
            .n7891(n7891), .n7885(n7885), .n7887(n7887), .n7865(n7865), 
            .n7867(n7867), .n3861(n3861), .n7883(n7883), .n7877(n7877), 
            .n7873(n7873), .n7879(n7879), .n7875(n7875), .n8724(n8724), 
            .n3863(n3863), .n4646(n4646), .n7899(n7899), .n7897(n7897), 
            .n7909(n7909), .n7911(n7911), .n165(n165_adj_1295), .n162(n162_adj_1294), 
            .n159(n159_adj_1293), .n156(n156_adj_1292), .n153(n153_adj_1291), 
            .n150(n150_adj_1290), .n147(n147_adj_1289), .n144(n144), .n141(n141), 
            .n138(n138), .n135(n135), .n132(n132), .n129(n129), .n126(n126_adj_1288), 
            .n123(n123), .n120(n120_adj_1287), .n117(n117), .n114(n114_adj_1286), 
            .n111(n111), .n108(n108_adj_1285), .n105(n105), .n102(n102_adj_1284), 
            .n99(n99_adj_1283), .n96(n96_adj_1282), .n93(n93_adj_1281), 
            .n90(n90_adj_1280), .n87(n87_adj_1279), .n84(n84_adj_1278), 
            .n81(n81_adj_1277), .n78(n78_adj_1276), .n75(n75_adj_1275), 
            .n72(n72_adj_1274), .n7881(n7881), .\proximo_estado_2__N_952[0] (proximo_estado_2__N_952[0]), 
            .n7889(n7889), .n8033(n8033), .GND_net(GND_net), .VCC_net(VCC_net), 
            .n7905(n7905), .n7869(n7869), .n7871(n7871), .n7893(n7893), 
            .n7895(n7895), .n7907(n7907), .n7861(n7861), .n8040(n8040), 
            .clk_c_enable_432(clk_c_enable_432), .n7863(n7863), .n7857(n7857), 
            .n7859(n7859), .n7901(n7901), .n7853(n7853), .n7855(n7855), 
            .n7903(n7903), .n7849(n7849));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(56[17] 64[6])
    FD1S3AX state_FSM_i7_rep_25 (.D(n2808), .CK(clk_c), .Q(clk_c_enable_348));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i7_rep_25.GSR = "ENABLED";
    FD1S3AX state_FSM_i2_rep_22 (.D(n2820), .CK(clk_c), .Q(n8817));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i2_rep_22.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i3 (.D(b_inv_15__N_503[34]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i3.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i4 (.D(b_inv_15__N_503[35]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i4.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i5 (.D(b_inv_15__N_503[36]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i5.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i6 (.D(b_inv_15__N_503[37]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i6.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i7 (.D(b_inv_15__N_503[38]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i7.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i8 (.D(b_inv_15__N_503[39]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i8.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i9 (.D(b_inv_15__N_503[40]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i9.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i10 (.D(b_inv_15__N_503[41]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i10.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i11 (.D(b_inv_15__N_503[42]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i11.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i12 (.D(b_inv_15__N_503[43]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i12.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i13 (.D(b_inv_15__N_503[44]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i13.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i14 (.D(b_inv_15__N_503[45]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i14.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i15 (.D(b_inv_15__N_503[46]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i15.GSR = "ENABLED";
    FD1P3AX b_inv_reg_res4_i0_i16 (.D(b_inv_15__N_503[47]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(b_inv_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam b_inv_reg_res4_i0_i16.GSR = "ENABLED";
    FD1P3AX prod_b__1_res7_e3__i2 (.D(n178_adj_1117), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[16]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i2.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i3 (.D(n177), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_b[17]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i3.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i4 (.D(n176), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_b[18]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i4.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i5 (.D(n175), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_b[19]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i5.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i6 (.D(n174), .SP(clk_c_enable_395), .CK(clk_c), 
            .Q(prod_b[20]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i6.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i7 (.D(n173_adj_1118), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[21]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i7.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i8 (.D(n172_adj_1119), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[22]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i8.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i9 (.D(n171_adj_1120), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[23]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i9.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i10 (.D(n170_adj_1121), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[24]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i10.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i11 (.D(n169_adj_1122), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[25]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i11.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i12 (.D(n168_adj_1123), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[26]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i12.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i13 (.D(n167_adj_1124), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[27]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i13.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i14 (.D(n166_adj_1125), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[28]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i14.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i15 (.D(n165_adj_1126), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[29]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i15.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i16 (.D(n164_adj_1127), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[30]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i16.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i17 (.D(n163_adj_1128), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[31]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i17.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i18 (.D(n162_adj_1129), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[32]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i18.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i19 (.D(n161_adj_1130), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i19.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i20 (.D(n160_adj_1131), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[34]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i20.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i21 (.D(n159_adj_1132), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i21.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i22 (.D(n158_adj_1133), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[36]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i22.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i23 (.D(n157_adj_1134), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i23.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i24 (.D(n156_adj_1135), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[38]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i24.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i25 (.D(n155_adj_1136), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i25.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i26 (.D(n154_adj_1137), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[40]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i26.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i27 (.D(n153_adj_1138), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i27.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i28 (.D(n152_adj_1139), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[42]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i28.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i29 (.D(n151_adj_1140), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i29.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i30 (.D(n150_adj_1141), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[44]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i30.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i31 (.D(n149_adj_1142), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i31.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i32 (.D(n148_adj_1143), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[46]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i32.GSR = "DISABLED";
    FD1P3AX prod_b__1_res7_e3__i33 (.D(n147_adj_1144), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_b[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(104[31:44])
    defparam prod_b__1_res7_e3__i33.GSR = "DISABLED";
    FD1P3AX a_inv_reg_res1_i0_i2 (.D(a_inv_15__N_487[33]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i2.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i3 (.D(a_inv_15__N_487[34]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i3.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i4 (.D(a_inv_15__N_487[35]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i4.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i5 (.D(a_inv_15__N_487[36]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i5.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i6 (.D(a_inv_15__N_487[37]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i6.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i7 (.D(a_inv_15__N_487[38]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i7.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i8 (.D(a_inv_15__N_487[39]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i8.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i9 (.D(a_inv_15__N_487[40]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i9.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i10 (.D(a_inv_15__N_487[41]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i10.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i11 (.D(a_inv_15__N_487[42]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i11.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i12 (.D(a_inv_15__N_487[43]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i12.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i13 (.D(a_inv_15__N_487[44]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i13.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i14 (.D(a_inv_15__N_487[45]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i14.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i15 (.D(a_inv_15__N_487[46]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i15.GSR = "ENABLED";
    FD1P3AX a_inv_reg_res1_i0_i16 (.D(a_inv_15__N_487[47]), .SP(clk_c_enable_348), 
            .CK(clk_c), .Q(a_inv_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_inv_reg_res1_i0_i16.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i2 (.D(c_inv_15__N_519[33]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_1));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i2.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i3 (.D(c_inv_15__N_519[34]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_2));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i3.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i4 (.D(c_inv_15__N_519[35]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_3));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i4.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i5 (.D(c_inv_15__N_519[36]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_4));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i5.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i6 (.D(c_inv_15__N_519[37]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_5));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i6.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i7 (.D(c_inv_15__N_519[38]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_6));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i7.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i8 (.D(c_inv_15__N_519[39]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_7));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i8.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i9 (.D(c_inv_15__N_519[40]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_8));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i9.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i10 (.D(c_inv_15__N_519[41]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_9));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i10.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i11 (.D(c_inv_15__N_519[42]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_10));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i11.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i12 (.D(c_inv_15__N_519[43]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_11));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i12.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i13 (.D(c_inv_15__N_519[44]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_12));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i13.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i14 (.D(c_inv_15__N_519[45]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_13));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i14.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i15 (.D(c_inv_15__N_519[46]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_14));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i15.GSR = "ENABLED";
    FD1P3AX c_inv_reg_res3_i0_i16 (.D(c_inv_15__N_519[47]), .SP(clk_c_enable_363), 
            .CK(clk_c), .Q(c_inv_c_15));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam c_inv_reg_res3_i0_i16.GSR = "ENABLED";
    FD1S3AX state_FSM_i2 (.D(n2820), .CK(clk_c), .Q(clk_c_enable_431));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1S3AX state_FSM_i3 (.D(clk_c_enable_431), .CK(clk_c), .Q(clk_c_enable_145));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3AX state_FSM_i4 (.D(n7916), .CK(clk_c), .Q(n2810));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(next_state_2__N_65[2]), .CK(clk_c), .CD(n8032), 
            .Q(n2809));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3AX state_FSM_i6 (.D(n2809), .CK(clk_c), .Q(n2808));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3AX state_FSM_i7 (.D(n2808), .CK(clk_c), .Q(clk_c_enable_363));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1P3AX prod_a__0_res5_e3__i2 (.D(n178_adj_1179), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[16]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i2.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i3 (.D(n177_adj_1180), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[17]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i3.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i4 (.D(n176_adj_1181), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[18]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i4.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i5 (.D(n175_adj_1182), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[19]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i5.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i6 (.D(n174_adj_1183), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[20]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i6.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i7 (.D(n173_adj_1184), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[21]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i7.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i8 (.D(n172_adj_1185), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[22]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i8.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i9 (.D(n171_adj_1186), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[23]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i9.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i10 (.D(n170_adj_1187), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[24]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i10.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i11 (.D(n169_adj_1188), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[25]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i11.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i12 (.D(n168_adj_1189), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[26]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i12.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i13 (.D(n167_adj_1190), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[27]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i13.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i14 (.D(n166_adj_1191), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[28]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i14.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i15 (.D(n165_adj_1192), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[29]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i15.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i16 (.D(n164_adj_1193), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[30]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i16.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i17 (.D(n163_adj_1194), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[31]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i17.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i18 (.D(n162_adj_1195), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[32]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i18.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i19 (.D(n161_adj_1196), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i19.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i20 (.D(n160_adj_1197), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[34]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i20.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i21 (.D(n159_adj_1198), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i21.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i22 (.D(n158_adj_1199), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[36]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i22.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i23 (.D(n157_adj_1200), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i23.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i24 (.D(n156_adj_1201), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[38]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i24.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i25 (.D(n155_adj_1202), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i25.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i26 (.D(n154_adj_1203), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[40]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i26.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i27 (.D(n153_adj_1204), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i27.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i28 (.D(n152_adj_1205), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[42]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i28.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i29 (.D(n151_adj_1206), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i29.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i30 (.D(n150_adj_1207), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[44]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i30.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i31 (.D(n149_adj_1208), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i31.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i32 (.D(n148_adj_1209), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[46]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i32.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e3__i33 (.D(n147_adj_1210), .SP(clk_c_enable_395), 
            .CK(clk_c), .Q(prod_a[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e3__i33.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i2 (.D(d_reg[1]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n128_adj_1212));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i2.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i3 (.D(d_reg[2]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n126_adj_1213));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i3.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i4 (.D(d_reg[3]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n124_adj_1214));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i4.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i5 (.D(d_reg[4]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n122_adj_1215));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i5.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i6 (.D(d_reg[5]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n120_adj_1216));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i6.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i7 (.D(d_reg[6]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n118_adj_1217));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i7.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i8 (.D(d_reg[7]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n116_adj_1218));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i8.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i9 (.D(d_reg[8]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n114_adj_1219));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i9.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i10 (.D(d_reg[9]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n112_adj_1220));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i10.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i11 (.D(d_reg[10]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n110_adj_1221));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i11.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i12 (.D(d_reg[11]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n108_adj_1222));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i12.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i13 (.D(d_reg[12]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n106_adj_1223));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i13.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i14 (.D(d_reg[13]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n104_adj_1224));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i14.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i15 (.D(d_reg[14]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n102_adj_1225));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i15.GSR = "DISABLED";
    FD1P3AX prod_a__0_res5_e2__i16 (.D(d_reg[15]), .SP(clk_c_enable_410), 
            .CK(clk_c), .Q(n68_adj_1226));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(103[31:44])
    defparam prod_a__0_res5_e2__i16.GSR = "DISABLED";
    CCU2C add_852_35 (.A0(regA[32]), .B0(n4646), .C0(n4578), .D0(n8724), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n8381), 
          .S0(n72_adj_1274));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_35.INIT0 = 16'h74b8;
    defparam add_852_35.INIT1 = 16'h0000;
    defparam add_852_35.INJECT1_0 = "NO";
    defparam add_852_35.INJECT1_1 = "NO";
    CCU2C add_852_33 (.A0(regA[30]), .B0(n4646), .C0(n4580), .D0(n7909), 
          .A1(regA[31]), .B1(n4646), .C1(n4579), .D1(n7911), .CIN(n8380), 
          .COUT(n8381), .S0(n78_adj_1276), .S1(n75_adj_1275));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_33.INIT0 = 16'h74b8;
    defparam add_852_33.INIT1 = 16'h74b8;
    defparam add_852_33.INJECT1_0 = "NO";
    defparam add_852_33.INJECT1_1 = "NO";
    CCU2C add_852_31 (.A0(regA[28]), .B0(n4646), .C0(n4582), .D0(n7905), 
          .A1(regA[29]), .B1(n4646), .C1(n4581), .D1(n7907), .CIN(n8379), 
          .COUT(n8380), .S0(n84_adj_1278), .S1(n81_adj_1277));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_31.INIT0 = 16'h74b8;
    defparam add_852_31.INIT1 = 16'h74b8;
    defparam add_852_31.INJECT1_0 = "NO";
    defparam add_852_31.INJECT1_1 = "NO";
    CCU2C add_852_29 (.A0(regA[26]), .B0(n4646), .C0(n4584), .D0(n7901), 
          .A1(regA[27]), .B1(n4646), .C1(n4583), .D1(n7903), .CIN(n8378), 
          .COUT(n8379), .S0(n90_adj_1280), .S1(n87_adj_1279));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_29.INIT0 = 16'h74b8;
    defparam add_852_29.INIT1 = 16'h74b8;
    defparam add_852_29.INJECT1_0 = "NO";
    defparam add_852_29.INJECT1_1 = "NO";
    CCU2C add_852_27 (.A0(regA[24]), .B0(n4646), .C0(n4586), .D0(n7897), 
          .A1(regA[25]), .B1(n4646), .C1(n4585), .D1(n7899), .CIN(n8377), 
          .COUT(n8378), .S0(n96_adj_1282), .S1(n93_adj_1281));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_27.INIT0 = 16'h74b8;
    defparam add_852_27.INIT1 = 16'h74b8;
    defparam add_852_27.INJECT1_0 = "NO";
    defparam add_852_27.INJECT1_1 = "NO";
    CCU2C add_852_25 (.A0(regA[22]), .B0(n4646), .C0(n4588), .D0(n7893), 
          .A1(regA[23]), .B1(n4646), .C1(n4587), .D1(n7895), .CIN(n8376), 
          .COUT(n8377), .S0(n102_adj_1284), .S1(n99_adj_1283));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_25.INIT0 = 16'h74b8;
    defparam add_852_25.INIT1 = 16'h74b8;
    defparam add_852_25.INJECT1_0 = "NO";
    defparam add_852_25.INJECT1_1 = "NO";
    CCU2C add_852_23 (.A0(regA[20]), .B0(n4646), .C0(n4590), .D0(n7861), 
          .A1(regA[21]), .B1(n4646), .C1(n4589), .D1(n7863), .CIN(n8375), 
          .COUT(n8376), .S0(n108_adj_1285), .S1(n105));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_23.INIT0 = 16'h74b8;
    defparam add_852_23.INIT1 = 16'h74b8;
    defparam add_852_23.INJECT1_0 = "NO";
    defparam add_852_23.INJECT1_1 = "NO";
    CCU2C add_852_21 (.A0(regA[18]), .B0(n4646), .C0(n4592), .D0(n7857), 
          .A1(regA[19]), .B1(n4646), .C1(n4591), .D1(n7859), .CIN(n8374), 
          .COUT(n8375), .S0(n114_adj_1286), .S1(n111));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_21.INIT0 = 16'h74b8;
    defparam add_852_21.INIT1 = 16'h74b8;
    defparam add_852_21.INJECT1_0 = "NO";
    defparam add_852_21.INJECT1_1 = "NO";
    CCU2C add_852_19 (.A0(regA[16]), .B0(n4646), .C0(n4594), .D0(n7853), 
          .A1(regA[17]), .B1(n4646), .C1(n4593), .D1(n7855), .CIN(n8373), 
          .COUT(n8374), .S0(n120_adj_1287), .S1(n117));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_19.INIT0 = 16'h74b8;
    defparam add_852_19.INIT1 = 16'h74b8;
    defparam add_852_19.INJECT1_0 = "NO";
    defparam add_852_19.INJECT1_1 = "NO";
    CCU2C add_852_17 (.A0(regA[14]), .B0(n4646), .C0(n4596), .D0(n7849), 
          .A1(regA[15]), .B1(n4646), .C1(n4595), .D1(n7851), .CIN(n8372), 
          .COUT(n8373), .S0(n126_adj_1288), .S1(n123));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_17.INIT0 = 16'h74b8;
    defparam add_852_17.INIT1 = 16'h74b8;
    defparam add_852_17.INJECT1_0 = "NO";
    defparam add_852_17.INJECT1_1 = "NO";
    CCU2C add_852_15 (.A0(regA[12]), .B0(n4646), .C0(n4598), .D0(n7889), 
          .A1(regA[13]), .B1(n4646), .C1(n4597), .D1(n7891), .CIN(n8371), 
          .COUT(n8372), .S0(n132), .S1(n129));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_15.INIT0 = 16'h74b8;
    defparam add_852_15.INIT1 = 16'h74b8;
    defparam add_852_15.INJECT1_0 = "NO";
    defparam add_852_15.INJECT1_1 = "NO";
    CCU2C add_852_13 (.A0(regA[10]), .B0(n4646), .C0(n4600), .D0(n7885), 
          .A1(regA[11]), .B1(n4646), .C1(n4599), .D1(n7887), .CIN(n8370), 
          .COUT(n8371), .S0(n138), .S1(n135));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_13.INIT0 = 16'h74b8;
    defparam add_852_13.INIT1 = 16'h74b8;
    defparam add_852_13.INJECT1_0 = "NO";
    defparam add_852_13.INJECT1_1 = "NO";
    CCU2C add_852_11 (.A0(regA[8]), .B0(n4646), .C0(n4602), .D0(n7881), 
          .A1(regA[9]), .B1(n4646), .C1(n4601), .D1(n7883), .CIN(n8369), 
          .COUT(n8370), .S0(n144), .S1(n141));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_11.INIT0 = 16'h74b8;
    defparam add_852_11.INIT1 = 16'h74b8;
    defparam add_852_11.INJECT1_0 = "NO";
    defparam add_852_11.INJECT1_1 = "NO";
    CCU2C add_852_9 (.A0(regA[6]), .B0(n4646), .C0(n4604), .D0(n7877), 
          .A1(regA[7]), .B1(n4646), .C1(n4603), .D1(n7879), .CIN(n8368), 
          .COUT(n8369), .S0(n150_adj_1290), .S1(n147_adj_1289));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_9.INIT0 = 16'h74b8;
    defparam add_852_9.INIT1 = 16'h74b8;
    defparam add_852_9.INJECT1_0 = "NO";
    defparam add_852_9.INJECT1_1 = "NO";
    CCU2C add_852_7 (.A0(regA[4]), .B0(n4646), .C0(n4606), .D0(n7873), 
          .A1(regA[5]), .B1(n4646), .C1(n4605), .D1(n7875), .CIN(n8367), 
          .COUT(n8368), .S0(n156_adj_1292), .S1(n153_adj_1291));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_7.INIT0 = 16'h74b8;
    defparam add_852_7.INIT1 = 16'h74b8;
    defparam add_852_7.INJECT1_0 = "NO";
    defparam add_852_7.INJECT1_1 = "NO";
    CCU2C add_852_5 (.A0(regA[2]), .B0(n4646), .C0(n4608), .D0(n7869), 
          .A1(regA[3]), .B1(n4646), .C1(n4607), .D1(n7871), .CIN(n8366), 
          .COUT(n8367), .S0(n162_adj_1294), .S1(n159_adj_1293));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_5.INIT0 = 16'h74b8;
    defparam add_852_5.INIT1 = 16'h74b8;
    defparam add_852_5.INJECT1_0 = "NO";
    defparam add_852_5.INJECT1_1 = "NO";
    CCU2C add_852_3 (.A0(regA[0]), .B0(n4646), .C0(n4610), .D0(n7865), 
          .A1(regA[1]), .B1(n4646), .C1(n4609), .D1(n7867), .CIN(n8365), 
          .COUT(n8366), .S0(n168_adj_1296), .S1(n165_adj_1295));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_3.INIT0 = 16'h74b8;
    defparam add_852_3.INIT1 = 16'h74b8;
    defparam add_852_3.INJECT1_0 = "NO";
    defparam add_852_3.INJECT1_1 = "NO";
    CCU2C add_852_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n3860), .B1(n3859), .C1(n3863), .D1(n8724), .COUT(n8365));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam add_852_1.INIT0 = 16'h0000;
    defparam add_852_1.INIT1 = 16'h01ff;
    defparam add_852_1.INJECT1_0 = "NO";
    defparam add_852_1.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_32 (.A0(prod_d[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8360), .S0(d_inv_15__N_535[46]), .S1(d_inv_15__N_535[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_30 (.A0(prod_d[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8359), .COUT(n8360), .S0(d_inv_15__N_535[44]), 
          .S1(d_inv_15__N_535[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_28 (.A0(prod_d[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8358), .COUT(n8359), .S0(d_inv_15__N_535[42]), 
          .S1(d_inv_15__N_535[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_26 (.A0(prod_d[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8357), .COUT(n8358), .S0(d_inv_15__N_535[40]), 
          .S1(d_inv_15__N_535[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_24 (.A0(prod_d[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8356), .COUT(n8357), .S0(d_inv_15__N_535[38]), 
          .S1(d_inv_15__N_535[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_22 (.A0(prod_d[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8355), .COUT(n8356), .S0(d_inv_15__N_535[36]), 
          .S1(d_inv_15__N_535[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_20 (.A0(prod_d[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8354), .COUT(n8355), .S0(d_inv_15__N_535[34]), 
          .S1(d_inv_15__N_535[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_18 (.A0(prod_d[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8353), .COUT(n8354), .S0(d_inv_15__N_535[32]), 
          .S1(d_inv_15__N_535[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_16 (.A0(prod_d[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8352), .COUT(n8353));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_14 (.A0(prod_d[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8351), .COUT(n8352));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_12 (.A0(prod_d[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8350), .COUT(n8351));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_10 (.A0(prod_d[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8349), .COUT(n8350));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_8 (.A0(prod_d[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8348), .COUT(n8349));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_6 (.A0(prod_d[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8347), .COUT(n8348));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_4 (.A0(prod_d[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8346), .COUT(n8347));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_440_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_440_add_4_2 (.A0(prod_d[15]), .B0(prod_d[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_d[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n8346));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_440_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_440_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_440_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_440_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_32 (.A0(prod_c[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8344), .S0(c_inv_15__N_519[46]), .S1(c_inv_15__N_519[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_30 (.A0(prod_c[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8343), .COUT(n8344), .S0(c_inv_15__N_519[44]), 
          .S1(c_inv_15__N_519[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_28 (.A0(prod_c[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8342), .COUT(n8343), .S0(c_inv_15__N_519[42]), 
          .S1(c_inv_15__N_519[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_26 (.A0(prod_c[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8341), .COUT(n8342), .S0(c_inv_15__N_519[40]), 
          .S1(c_inv_15__N_519[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_24 (.A0(prod_c[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8340), .COUT(n8341), .S0(c_inv_15__N_519[38]), 
          .S1(c_inv_15__N_519[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_24.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_13 (.A0(b_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8291), .COUT(n8292), .S0(n53_adj_1245), 
          .S1(n50_adj_1244));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_13.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_13.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_13.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_13.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_11 (.A0(b_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8290), .COUT(n8291), .S0(n59_adj_1247), 
          .S1(n56_adj_1246));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_11.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_11.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_11.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_11.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_9 (.A0(b_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8289), .COUT(n8290), .S0(n65_adj_1249), .S1(n62_adj_1248));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_9.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_9.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_9.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_9.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_7 (.A0(b_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8288), .COUT(n8289), .S0(n71_adj_1251), .S1(n68_adj_1250));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_7.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_7.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_7.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_7.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_5 (.A0(b_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8287), .COUT(n8288), .S0(n77_adj_1253), .S1(n74_adj_1252));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_5.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_5.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_5.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_5.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_3 (.A0(b_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8286), .COUT(n8287), .S0(n83_adj_1255), .S1(n80_adj_1254));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_3.INIT0 = 16'h5555;
    defparam b_s_res8_e3_add_4_3.INIT1 = 16'h5555;
    defparam b_s_res8_e3_add_4_3.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_3.INJECT1_1 = "NO";
    CCU2C b_s_res8_e3_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n8286), .S1(n86_adj_1256));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(98[28:55])
    defparam b_s_res8_e3_add_4_1.INIT0 = 16'h0000;
    defparam b_s_res8_e3_add_4_1.INIT1 = 16'haaa5;
    defparam b_s_res8_e3_add_4_1.INJECT1_0 = "NO";
    defparam b_s_res8_e3_add_4_1.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_17 (.A0(c_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8284), .S0(n41_adj_1258), .S1(n38_adj_1257));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_17.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_17.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_17.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_17.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_15 (.A0(c_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8283), .COUT(n8284), .S0(n47_adj_1260), 
          .S1(n44_adj_1259));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_15.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_15.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_15.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_15.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_13 (.A0(c_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8282), .COUT(n8283), .S0(n53_adj_1262), 
          .S1(n50_adj_1261));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_13.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_13.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_13.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_13.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_11 (.A0(c_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8281), .COUT(n8282), .S0(n59_adj_1264), 
          .S1(n56_adj_1263));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_11.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_11.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_11.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_11.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_9 (.A0(c_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8280), .COUT(n8281), .S0(n65_adj_1266), .S1(n62_adj_1265));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_9.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_9.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_9.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_9.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_7 (.A0(c_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8279), .COUT(n8280), .S0(n71_adj_1268), .S1(n68_adj_1267));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_7.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_7.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_7.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_7.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_5 (.A0(c_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8278), .COUT(n8279), .S0(n77_adj_1270), .S1(n74_adj_1269));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_5.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_5.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_5.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_5.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_3 (.A0(c_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n8277), .COUT(n8278), .S0(n83_adj_1272), .S1(n80_adj_1271));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_3.INIT0 = 16'h5555;
    defparam c_s_res10_e3_add_4_3.INIT1 = 16'h5555;
    defparam c_s_res10_e3_add_4_3.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_3.INJECT1_1 = "NO";
    CCU2C c_s_res10_e3_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n8277), .S1(n86_adj_1273));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(99[28:55])
    defparam c_s_res10_e3_add_4_1.INIT0 = 16'h0000;
    defparam c_s_res10_e3_add_4_1.INIT1 = 16'haaa5;
    defparam c_s_res10_e3_add_4_1.INJECT1_0 = "NO";
    defparam c_s_res10_e3_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_32 (.A0(prod_a[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8275), .S0(a_inv_15__N_487[46]), .S1(a_inv_15__N_487[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_30 (.A0(prod_a[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8274), .COUT(n8275), .S0(a_inv_15__N_487[44]), 
          .S1(a_inv_15__N_487[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_28 (.A0(prod_a[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8273), .COUT(n8274), .S0(a_inv_15__N_487[42]), 
          .S1(a_inv_15__N_487[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_26 (.A0(prod_a[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8272), .COUT(n8273), .S0(a_inv_15__N_487[40]), 
          .S1(a_inv_15__N_487[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_24 (.A0(prod_a[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8271), .COUT(n8272), .S0(a_inv_15__N_487[38]), 
          .S1(a_inv_15__N_487[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_22 (.A0(prod_a[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8270), .COUT(n8271), .S0(a_inv_15__N_487[36]), 
          .S1(a_inv_15__N_487[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_20 (.A0(prod_a[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8269), .COUT(n8270), .S0(a_inv_15__N_487[34]), 
          .S1(a_inv_15__N_487[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_18 (.A0(prod_a[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8268), .COUT(n8269), .S0(a_inv_15__N_487[32]), 
          .S1(a_inv_15__N_487[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_16 (.A0(prod_a[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8267), .COUT(n8268));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_14 (.A0(prod_a[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8266), .COUT(n8267));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_12 (.A0(prod_a[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8265), .COUT(n8266));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_10 (.A0(prod_a[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8264), .COUT(n8265));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_8 (.A0(prod_a[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8263), .COUT(n8264));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_6 (.A0(prod_a[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8262), .COUT(n8263));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_4 (.A0(prod_a[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8261), .COUT(n8262));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_437_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_437_add_4_2 (.A0(prod_a[15]), .B0(prod_a[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_a[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n8261));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_437_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_437_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_437_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_437_add_4_2.INJECT1_1 = "NO";
    FD1P3AX a_reg_i0_i1 (.D(a_c_1), .SP(clk_c_enable_411), .CK(clk_c), 
            .Q(a_reg[1]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_452_add_4_22 (.A0(prod_c[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8339), .COUT(n8340), .S0(c_inv_15__N_519[36]), 
          .S1(c_inv_15__N_519[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_20 (.A0(prod_c[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8338), .COUT(n8339), .S0(c_inv_15__N_519[34]), 
          .S1(c_inv_15__N_519[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_18 (.A0(prod_c[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8337), .COUT(n8338), .S0(c_inv_15__N_519[32]), 
          .S1(c_inv_15__N_519[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_16 (.A0(prod_c[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8336), .COUT(n8337));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_14 (.A0(prod_c[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8335), .COUT(n8336));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_12 (.A0(prod_c[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8334), .COUT(n8335));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_10 (.A0(prod_c[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8333), .COUT(n8334));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_8 (.A0(prod_c[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8332), .COUT(n8333));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_6 (.A0(prod_c[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8331), .COUT(n8332));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_4 (.A0(prod_c[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8330), .COUT(n8331));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_452_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_452_add_4_2 (.A0(prod_c[15]), .B0(prod_c[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_c[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n8330));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_452_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_452_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_452_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_452_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_34 (.A0(n70), .B0(n37), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n8329), 
          .S0(det_q4_28_31__N_551[31]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_34.INIT1 = 16'h0000;
    defparam _add_1_455_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_32 (.A0(n72), .B0(n39), .C0(GND_net), .D0(VCC_net), 
          .A1(n71), .B1(n38), .C1(GND_net), .D1(VCC_net), .CIN(n8328), 
          .COUT(n8329), .S0(det_q4_28_31__N_551[29]), .S1(det_q4_28_31__N_551[30]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_30 (.A0(n74), .B0(n41), .C0(GND_net), .D0(VCC_net), 
          .A1(n73), .B1(n40), .C1(GND_net), .D1(VCC_net), .CIN(n8327), 
          .COUT(n8328), .S0(det_q4_28_31__N_551[27]), .S1(det_q4_28_31__N_551[28]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_28 (.A0(n76), .B0(n43), .C0(GND_net), .D0(VCC_net), 
          .A1(n75), .B1(n42), .C1(GND_net), .D1(VCC_net), .CIN(n8326), 
          .COUT(n8327), .S0(det_q4_28_31__N_551[25]), .S1(det_q4_28_31__N_551[26]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_26 (.A0(n78), .B0(n45), .C0(GND_net), .D0(VCC_net), 
          .A1(n77), .B1(n44), .C1(GND_net), .D1(VCC_net), .CIN(n8325), 
          .COUT(n8326), .S0(det_q4_28_31__N_551[23]), .S1(det_q4_28_31__N_551[24]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_24 (.A0(n80), .B0(n47), .C0(GND_net), .D0(VCC_net), 
          .A1(n79), .B1(n46), .C1(GND_net), .D1(VCC_net), .CIN(n8324), 
          .COUT(n8325), .S0(det_q4_28_31__N_551[21]), .S1(det_q4_28_31__N_551[22]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_22 (.A0(n82), .B0(n49), .C0(GND_net), .D0(VCC_net), 
          .A1(n81), .B1(n48), .C1(GND_net), .D1(VCC_net), .CIN(n8323), 
          .COUT(n8324), .S0(det_q4_28_31__N_551[19]), .S1(det_q4_28_31__N_551[20]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_20 (.A0(n84), .B0(n51), .C0(GND_net), .D0(VCC_net), 
          .A1(n83), .B1(n50), .C1(GND_net), .D1(VCC_net), .CIN(n8322), 
          .COUT(n8323), .S0(det_q4_28_31__N_551[17]), .S1(det_q4_28_31__N_551[18]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_18 (.A0(n86), .B0(n53), .C0(GND_net), .D0(VCC_net), 
          .A1(n85), .B1(n52), .C1(GND_net), .D1(VCC_net), .CIN(n8321), 
          .COUT(n8322), .S0(det_q4_28_31__N_551[15]), .S1(det_q4_28_31__N_551[16]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_16 (.A0(n88), .B0(n55), .C0(GND_net), .D0(VCC_net), 
          .A1(n87), .B1(n54), .C1(GND_net), .D1(VCC_net), .CIN(n8320), 
          .COUT(n8321), .S0(det_q4_28_31__N_551[13]), .S1(det_q4_28_31__N_551[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_14 (.A0(n90), .B0(n57), .C0(GND_net), .D0(VCC_net), 
          .A1(n89), .B1(n56), .C1(GND_net), .D1(VCC_net), .CIN(n8319), 
          .COUT(n8320), .S0(det_q4_28_31__N_551[11]), .S1(det_q4_28_31__N_551[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_12 (.A0(n92), .B0(n59), .C0(GND_net), .D0(VCC_net), 
          .A1(n91), .B1(n58), .C1(GND_net), .D1(VCC_net), .CIN(n8318), 
          .COUT(n8319), .S0(det_q4_28_31__N_551[9]), .S1(det_q4_28_31__N_551[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_10 (.A0(n94), .B0(n61), .C0(GND_net), .D0(VCC_net), 
          .A1(n93), .B1(n60), .C1(GND_net), .D1(VCC_net), .CIN(n8317), 
          .COUT(n8318), .S0(det_q4_28_31__N_551[7]), .S1(det_q4_28_31__N_551[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_8 (.A0(n96), .B0(n63), .C0(GND_net), .D0(VCC_net), 
          .A1(n95), .B1(n62), .C1(GND_net), .D1(VCC_net), .CIN(n8316), 
          .COUT(n8317), .S0(det_q4_28_31__N_551[5]), .S1(det_q4_28_31__N_551[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_6 (.A0(n98), .B0(n65), .C0(GND_net), .D0(VCC_net), 
          .A1(n97), .B1(n64), .C1(GND_net), .D1(VCC_net), .CIN(n8315), 
          .COUT(n8316), .S0(det_q4_28_31__N_551[3]), .S1(det_q4_28_31__N_551[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_4 (.A0(n100), .B0(n67), .C0(GND_net), .D0(VCC_net), 
          .A1(n99), .B1(n66), .C1(GND_net), .D1(VCC_net), .CIN(n8314), 
          .COUT(n8315), .S0(det_q4_28_31__N_551[1]), .S1(det_q4_28_31__N_551[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_455_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_455_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n101), .B1(n68), .C1(GND_net), .D1(VCC_net), 
          .COUT(n8314), .S1(det_q4_28_31__N_551[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(89[37:70])
    defparam _add_1_455_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_455_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_455_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_455_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_32 (.A0(prod_b[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8312), .S0(b_inv_15__N_503[46]), .S1(b_inv_15__N_503[47]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_32.INIT0 = 16'haaa0;
    defparam _add_1_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_30 (.A0(prod_b[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8311), .COUT(n8312), .S0(b_inv_15__N_503[44]), 
          .S1(b_inv_15__N_503[45]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_30.INIT0 = 16'haaa0;
    defparam _add_1_add_4_30.INIT1 = 16'haaa0;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(prod_b[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8310), .COUT(n8311), .S0(b_inv_15__N_503[42]), 
          .S1(b_inv_15__N_503[43]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_28.INIT0 = 16'haaa0;
    defparam _add_1_add_4_28.INIT1 = 16'haaa0;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(prod_b[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8309), .COUT(n8310), .S0(b_inv_15__N_503[40]), 
          .S1(b_inv_15__N_503[41]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_26.INIT0 = 16'haaa0;
    defparam _add_1_add_4_26.INIT1 = 16'haaa0;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_24 (.A0(prod_b[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8308), .COUT(n8309), .S0(b_inv_15__N_503[38]), 
          .S1(b_inv_15__N_503[39]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_24.INIT0 = 16'haaa0;
    defparam _add_1_add_4_24.INIT1 = 16'haaa0;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_22 (.A0(prod_b[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8307), .COUT(n8308), .S0(b_inv_15__N_503[36]), 
          .S1(b_inv_15__N_503[37]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_add_4_22.INIT1 = 16'haaa0;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_20 (.A0(prod_b[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8306), .COUT(n8307), .S0(b_inv_15__N_503[34]), 
          .S1(b_inv_15__N_503[35]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_18 (.A0(prod_b[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8305), .COUT(n8306), .S0(b_inv_15__N_503[32]), 
          .S1(b_inv_15__N_503[33]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_16 (.A0(prod_b[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8304), .COUT(n8305));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_14 (.A0(prod_b[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8303), .COUT(n8304));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_12 (.A0(prod_b[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8302), .COUT(n8303));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_10 (.A0(prod_b[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8301), .COUT(n8302));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_8 (.A0(prod_b[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8300), .COUT(n8301));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_6 (.A0(prod_b[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8299), .COUT(n8300));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_4 (.A0(prod_b[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n8298), .COUT(n8299));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_2 (.A0(prod_b[15]), .B0(prod_b[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(prod_b[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n8298));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(50[19:38])
    defparam _add_1_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    LUT4 i701_3_lut (.A(n8033), .B(n3860), .C(n3863), .Z(n8040)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i701_3_lut.init = 16'h5454;
    LUT4 det_zero_reg_I_0_1_lut (.A(det_zero_reg), .Z(det_zero_reg_N_905)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(93[25:38])
    defparam det_zero_reg_I_0_1_lut.init = 16'h5555;
    LUT4 i279_2_lut (.A(n2809), .B(reset_c), .Z(clk_c_enable_410)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam i279_2_lut.init = 16'h2222;
    FD1S3AX state_FSM_i2_rep_23 (.D(n2820), .CK(clk_c), .Q(clk_c_enable_411));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(125[9] 134[16])
    defparam state_FSM_i2_rep_23.GSR = "ENABLED";
    LUT4 i274_2_lut (.A(n2808), .B(reset_c), .Z(clk_c_enable_395)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam i274_2_lut.init = 16'h2222;
    FD1P3AX a_reg_i0_i2 (.D(a_c_2), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i3 (.D(a_c_3), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[3]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i3.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i4 (.D(a_c_4), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i4.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i5 (.D(a_c_5), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i5.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i6 (.D(a_c_6), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[6]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i6.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i7 (.D(a_c_7), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[7]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i7.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i8 (.D(a_c_8), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[8]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i8.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i9 (.D(a_c_9), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[9]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i9.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i10 (.D(a_c_10), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[10]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i10.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i11 (.D(a_c_11), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[11]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i11.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i12 (.D(a_c_12), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[12]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i12.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i13 (.D(a_c_13), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[13]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i13.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i14 (.D(a_c_14), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[14]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i14.GSR = "ENABLED";
    FD1P3AX a_reg_i0_i15 (.D(a_c_15), .SP(clk_c_enable_431), .CK(clk_c), 
            .Q(a_reg[15]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam a_reg_i0_i15.GSR = "ENABLED";
    FD1S3IX start_NRDA_84 (.D(det_zero_reg_N_905), .CK(clk_c), .CD(n8032), 
            .Q(proximo_estado_2__N_952[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(77[18] 120[12])
    defparam start_NRDA_84.GSR = "ENABLED";
    LUT4 i1109_4_lut (.A(n49_adj_1230), .B(n62_adj_1298), .C(n58_adj_1236), 
         .D(n50_adj_1229), .Z(det_zero_reg_N_907)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i1109_4_lut.init = 16'h0001;
    LUT4 i17_4_lut (.A(det_q4_28_31__N_551[0]), .B(det_q4_28_31__N_551[25]), 
         .C(det_q4_28_31__N_551[27]), .D(det_q4_28_31__N_551[10]), .Z(n49_adj_1230)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(90[37:77])
    defparam i17_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module divNRDA_FSM
//

module divNRDA_FSM (regA, n4577, clk_c, n168, clk_c_enable_239, det_q4_28, 
            quotient_31__N_908, n3859, n3860, n7851, \next_state_2__N_65[2] , 
            n7891, n7885, n7887, n7865, n7867, n3861, n7883, n7877, 
            n7873, n7879, n7875, n8724, n3863, n4646, n7899, n7897, 
            n7909, n7911, n165, n162, n159, n156, n153, n150, 
            n147, n144, n141, n138, n135, n132, n129, n126, 
            n123, n120, n117, n114, n111, n108, n105, n102, 
            n99, n96, n93, n90, n87, n84, n81, n78, n75, n72, 
            n7881, \proximo_estado_2__N_952[0] , n7889, n8033, GND_net, 
            VCC_net, n7905, n7869, n7871, n7893, n7895, n7907, 
            n7861, n8040, clk_c_enable_432, n7863, n7857, n7859, 
            n7901, n7853, n7855, n7903, n7849);
    output [32:0]regA;
    output [32:0]n4577;
    input clk_c;
    input n168;
    output clk_c_enable_239;
    input [31:0]det_q4_28;
    output [31:0]quotient_31__N_908;
    output n3859;
    output n3860;
    output n7851;
    output \next_state_2__N_65[2] ;
    output n7891;
    output n7885;
    output n7887;
    output n7865;
    output n7867;
    output n3861;
    output n7883;
    output n7877;
    output n7873;
    output n7879;
    output n7875;
    output n8724;
    output n3863;
    output n4646;
    output n7899;
    output n7897;
    output n7909;
    output n7911;
    input n165;
    input n162;
    input n159;
    input n156;
    input n153;
    input n150;
    input n147;
    input n144;
    input n141;
    input n138;
    input n135;
    input n132;
    input n129;
    input n126;
    input n123;
    input n120;
    input n117;
    input n114;
    input n111;
    input n108;
    input n105;
    input n102;
    input n99;
    input n96;
    input n93;
    input n90;
    input n87;
    input n84;
    input n81;
    input n78;
    input n75;
    input n72;
    output n7881;
    input \proximo_estado_2__N_952[0] ;
    output n7889;
    output n8033;
    input GND_net;
    input VCC_net;
    output n7905;
    output n7869;
    output n7871;
    output n7893;
    output n7895;
    output n7907;
    output n7861;
    input n8040;
    input clk_c_enable_432;
    output n7863;
    output n7857;
    output n7859;
    output n7901;
    output n7853;
    output n7855;
    output n7903;
    output n7849;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(2[35:38])
    wire [7:0]n3858;
    
    wire clk_c_enable_192;
    wire [32:0]regM;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(27[14:18])
    wire [31:0]inv_det;   // d:/ci/rtl_fpga/projeto_final/kalman_core/matrix_inv.v(41[35:42])
    
    wire clk_c_enable_11, ready_N_1109;
    wire [5:0]i;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(25[8:9])
    
    wire n8726, n8562, clk_c_enable_417, n8729, n8723, n8554, n8532, 
        n8728, n8406;
    wire [2:0]proximo_estado_2__N_946;
    
    wire n3887, n7, n3888, n3892, n8452, n8528, n8399, n8448, 
        n8429, n3883, n38, n52, n46, n56, n42, n54, n60, n49, 
        n62, n58, n50, n41, n8550, n8526, n8297;
    wire [5:0]n29;
    
    wire n8296, n8295, n8568, n8034, A0_N_1113, n8524;
    
    LUT4 i782_2_lut (.A(regA[27]), .B(n3858[2]), .Z(n4577[28])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i782_2_lut.init = 16'h8888;
    FD1P3AX regA_i0_i0 (.D(n168), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i0.GSR = "ENABLED";
    FD1P3AX regM__i1 (.D(det_q4_28[0]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i1.GSR = "ENABLED";
    FD1S3AX regQ_i0 (.D(quotient_31__N_908[0]), .CK(clk_c), .Q(inv_det[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i0.GSR = "ENABLED";
    LUT4 i512_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[15]), .Z(n7851)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i512_2_lut_3_lut.init = 16'he1e1;
    FD1P3AX ready_61 (.D(ready_N_1109), .SP(clk_c_enable_11), .CK(clk_c), 
            .Q(\next_state_2__N_65[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam ready_61.GSR = "ENABLED";
    LUT4 i552_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[13]), .Z(n7891)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i552_2_lut_3_lut.init = 16'he1e1;
    LUT4 i546_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[10]), .Z(n7885)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i546_2_lut_3_lut.init = 16'he1e1;
    LUT4 i548_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[11]), .Z(n7887)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i548_2_lut_3_lut.init = 16'he1e1;
    LUT4 i526_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[0]), .Z(n7865)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i526_2_lut_3_lut.init = 16'he1e1;
    LUT4 i528_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[1]), .Z(n7867)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i528_2_lut_3_lut.init = 16'he1e1;
    LUT4 i3_2_lut_rep_20 (.A(i[3]), .B(i[4]), .Z(n8726)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(129[10:21])
    defparam i3_2_lut_rep_20.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(i[3]), .B(i[4]), .C(i[5]), .Z(n8562)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(129[10:21])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_21 (.A(clk_c_enable_239), .B(n3858[2]), .Z(clk_c_enable_417)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_21.init = 16'heeee;
    LUT4 i615_3_lut_4_lut_then_1_lut (.A(inv_det[16]), .Z(n8729)) /* synthesis lut_function=(A) */ ;
    defparam i615_3_lut_4_lut_then_1_lut.init = 16'haaaa;
    LUT4 i689_2_lut_rep_17_3_lut (.A(clk_c_enable_239), .B(n3858[2]), .C(n3861), 
         .Z(n8723)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i689_2_lut_rep_17_3_lut.init = 16'hf1f1;
    LUT4 i1_2_lut_3_lut_adj_4 (.A(i[5]), .B(regA[32]), .C(n3861), .Z(n8554)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_4.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_5 (.A(i[5]), .B(regA[32]), .C(i[1]), .Z(n8532)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_5.init = 16'h0808;
    LUT4 i783_2_lut (.A(regA[28]), .B(n3858[2]), .Z(n4577[29])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i783_2_lut.init = 16'h8888;
    LUT4 i544_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[9]), .Z(n7883)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i544_2_lut_3_lut.init = 16'he1e1;
    LUT4 i538_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[6]), .Z(n7877)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i538_2_lut_3_lut.init = 16'he1e1;
    LUT4 i534_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[4]), .Z(n7873)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i534_2_lut_3_lut.init = 16'he1e1;
    LUT4 i615_3_lut_4_lut_else_1_lut (.A(inv_det[16]), .B(n3858[2]), .C(inv_det[15]), 
         .D(clk_c_enable_239), .Z(n8728)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B (D))) */ ;
    defparam i615_3_lut_4_lut_else_1_lut.init = 16'hf3e2;
    LUT4 i540_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[7]), .Z(n7879)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i540_2_lut_3_lut.init = 16'he1e1;
    LUT4 i536_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[5]), .Z(n7875)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i536_2_lut_3_lut.init = 16'he1e1;
    LUT4 i1145_2_lut_rep_18 (.A(n3859), .B(n3860), .Z(n8724)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i1145_2_lut_rep_18.init = 16'h1111;
    LUT4 i354_2_lut_3_lut (.A(n3859), .B(n3860), .C(n3863), .Z(n4646)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i354_2_lut_3_lut.init = 16'hfefe;
    LUT4 i560_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[25]), .Z(n7899)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i560_2_lut_3_lut.init = 16'he1e1;
    LUT4 i558_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[24]), .Z(n7897)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i558_2_lut_3_lut.init = 16'he1e1;
    LUT4 i776_2_lut (.A(regA[21]), .B(n3858[2]), .Z(n4577[22])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i776_2_lut.init = 16'h8888;
    LUT4 i777_2_lut (.A(regA[22]), .B(n3858[2]), .Z(n4577[23])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i777_2_lut.init = 16'h8888;
    LUT4 i774_2_lut (.A(regA[19]), .B(n3858[2]), .Z(n4577[20])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i774_2_lut.init = 16'h8888;
    LUT4 i775_2_lut (.A(regA[20]), .B(n3858[2]), .Z(n4577[21])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i775_2_lut.init = 16'h8888;
    LUT4 i772_2_lut (.A(regA[17]), .B(n3858[2]), .Z(n4577[18])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i772_2_lut.init = 16'h8888;
    LUT4 i773_2_lut (.A(regA[18]), .B(n3858[2]), .Z(n4577[19])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i773_2_lut.init = 16'h8888;
    LUT4 i770_2_lut (.A(regA[15]), .B(n3858[2]), .Z(n4577[16])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i770_2_lut.init = 16'h8888;
    LUT4 i771_2_lut (.A(regA[16]), .B(n3858[2]), .Z(n4577[17])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i771_2_lut.init = 16'h8888;
    LUT4 i768_2_lut (.A(regA[13]), .B(n3858[2]), .Z(n4577[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i768_2_lut.init = 16'h8888;
    LUT4 i769_2_lut (.A(regA[14]), .B(n3858[2]), .Z(n4577[15])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i769_2_lut.init = 16'h8888;
    LUT4 i766_2_lut (.A(regA[11]), .B(n3858[2]), .Z(n4577[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i766_2_lut.init = 16'h8888;
    LUT4 i767_2_lut (.A(regA[12]), .B(n3858[2]), .Z(n4577[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i767_2_lut.init = 16'h8888;
    LUT4 i764_2_lut (.A(regA[9]), .B(n3858[2]), .Z(n4577[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i764_2_lut.init = 16'h8888;
    LUT4 i765_2_lut (.A(regA[10]), .B(n3858[2]), .Z(n4577[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i765_2_lut.init = 16'h8888;
    LUT4 i762_2_lut (.A(regA[7]), .B(n3858[2]), .Z(n4577[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i762_2_lut.init = 16'h8888;
    LUT4 i763_2_lut (.A(regA[8]), .B(n3858[2]), .Z(n4577[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i763_2_lut.init = 16'h8888;
    LUT4 i760_2_lut (.A(regA[5]), .B(n3858[2]), .Z(n4577[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i760_2_lut.init = 16'h8888;
    LUT4 i761_2_lut (.A(regA[6]), .B(n3858[2]), .Z(n4577[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i761_2_lut.init = 16'h8888;
    LUT4 i758_2_lut (.A(regA[3]), .B(n3858[2]), .Z(n4577[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i758_2_lut.init = 16'h8888;
    LUT4 i759_2_lut (.A(regA[4]), .B(n3858[2]), .Z(n4577[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i759_2_lut.init = 16'h8888;
    LUT4 i756_2_lut (.A(regA[1]), .B(n3858[2]), .Z(n4577[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i756_2_lut.init = 16'h8888;
    LUT4 i757_2_lut (.A(regA[2]), .B(n3858[2]), .Z(n4577[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i757_2_lut.init = 16'h8888;
    LUT4 i753_2_lut (.A(inv_det[31]), .B(n3858[2]), .Z(n4577[0])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i753_2_lut.init = 16'h8888;
    LUT4 i755_2_lut (.A(regA[0]), .B(n3858[2]), .Z(n4577[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i755_2_lut.init = 16'h8888;
    LUT4 i1_3_lut (.A(clk_c_enable_239), .B(n3861), .C(i[5]), .Z(n8406)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i1_3_lut.init = 16'haeae;
    LUT4 i232_2_lut (.A(proximo_estado_2__N_946[2]), .B(n3858[4]), .Z(n3887)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i232_2_lut.init = 16'h4444;
    LUT4 i233_4_lut (.A(n8562), .B(n3858[2]), .C(n7), .D(i[1]), .Z(n3888)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i233_4_lut.init = 16'hccc8;
    LUT4 i237_2_lut (.A(proximo_estado_2__N_946[2]), .B(n3858[4]), .Z(n3892)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i237_2_lut.init = 16'h8888;
    LUT4 i570_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[30]), .Z(n7909)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i570_2_lut_3_lut.init = 16'he1e1;
    LUT4 i572_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[31]), .Z(n7911)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i572_2_lut_3_lut.init = 16'he1e1;
    LUT4 i1_4_lut (.A(n7), .B(n8726), .C(i[1]), .D(n8554), .Z(n8452)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    FD1P3AX regA_i0_i1 (.D(n165), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i1.GSR = "ENABLED";
    FD1P3AX regA_i0_i2 (.D(n162), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i2.GSR = "ENABLED";
    FD1P3AX regA_i0_i3 (.D(n159), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i3.GSR = "ENABLED";
    FD1P3AX regA_i0_i4 (.D(n156), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i4.GSR = "ENABLED";
    FD1P3AX regA_i0_i5 (.D(n153), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i5.GSR = "ENABLED";
    FD1P3AX regA_i0_i6 (.D(n150), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i6.GSR = "ENABLED";
    FD1P3AX regA_i0_i7 (.D(n147), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i7.GSR = "ENABLED";
    FD1P3AX regA_i0_i8 (.D(n144), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i8.GSR = "ENABLED";
    FD1P3AX regA_i0_i9 (.D(n141), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i9.GSR = "ENABLED";
    FD1P3AX regA_i0_i10 (.D(n138), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i10.GSR = "ENABLED";
    FD1P3AX regA_i0_i11 (.D(n135), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i11.GSR = "ENABLED";
    FD1P3AX regA_i0_i12 (.D(n132), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i12.GSR = "ENABLED";
    FD1P3AX regA_i0_i13 (.D(n129), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i13.GSR = "ENABLED";
    FD1P3AX regA_i0_i14 (.D(n126), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i14.GSR = "ENABLED";
    FD1P3AX regA_i0_i15 (.D(n123), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i15.GSR = "ENABLED";
    FD1P3AX regA_i0_i16 (.D(n120), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i16.GSR = "ENABLED";
    FD1P3AX regA_i0_i17 (.D(n117), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i17.GSR = "ENABLED";
    FD1P3AX regA_i0_i18 (.D(n114), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i18.GSR = "ENABLED";
    FD1P3AX regA_i0_i19 (.D(n111), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i19.GSR = "ENABLED";
    FD1P3AX regA_i0_i20 (.D(n108), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i20.GSR = "ENABLED";
    FD1P3AX regA_i0_i21 (.D(n105), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i21.GSR = "ENABLED";
    FD1P3AX regA_i0_i22 (.D(n102), .SP(clk_c_enable_192), .CK(clk_c), 
            .Q(regA[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i22.GSR = "ENABLED";
    FD1P3AX regA_i0_i23 (.D(n99), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i23.GSR = "ENABLED";
    FD1P3AX regA_i0_i24 (.D(n96), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i24.GSR = "ENABLED";
    FD1P3AX regA_i0_i25 (.D(n93), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i25.GSR = "ENABLED";
    FD1P3AX regA_i0_i26 (.D(n90), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i26.GSR = "ENABLED";
    FD1P3AX regA_i0_i27 (.D(n87), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i27.GSR = "ENABLED";
    FD1P3AX regA_i0_i28 (.D(n84), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i28.GSR = "ENABLED";
    FD1P3AX regA_i0_i29 (.D(n81), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i29.GSR = "ENABLED";
    FD1P3AX regA_i0_i30 (.D(n78), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i30.GSR = "ENABLED";
    FD1P3AX regA_i0_i31 (.D(n75), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i31.GSR = "ENABLED";
    FD1P3AX regA_i0_i32 (.D(n72), .SP(clk_c_enable_192), .CK(clk_c), .Q(regA[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regA_i0_i32.GSR = "ENABLED";
    FD1P3AX regM__i2 (.D(det_q4_28[1]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i2.GSR = "ENABLED";
    FD1P3AX regM__i3 (.D(det_q4_28[2]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i3.GSR = "ENABLED";
    FD1P3AX regM__i4 (.D(det_q4_28[3]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i4.GSR = "ENABLED";
    FD1P3AX regM__i5 (.D(det_q4_28[4]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i5.GSR = "ENABLED";
    FD1P3AX regM__i6 (.D(det_q4_28[5]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i6.GSR = "ENABLED";
    FD1P3AX regM__i7 (.D(det_q4_28[6]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i7.GSR = "ENABLED";
    FD1P3AX regM__i8 (.D(det_q4_28[7]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i8.GSR = "ENABLED";
    FD1P3AX regM__i9 (.D(det_q4_28[8]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i9.GSR = "ENABLED";
    FD1P3AX regM__i10 (.D(det_q4_28[9]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i10.GSR = "ENABLED";
    FD1P3AX regM__i11 (.D(det_q4_28[10]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i11.GSR = "ENABLED";
    FD1P3AX regM__i12 (.D(det_q4_28[11]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i12.GSR = "ENABLED";
    FD1P3AX regM__i13 (.D(det_q4_28[12]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i13.GSR = "ENABLED";
    FD1P3AX regM__i14 (.D(det_q4_28[13]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i14.GSR = "ENABLED";
    FD1P3AX regM__i15 (.D(det_q4_28[14]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i15.GSR = "ENABLED";
    FD1P3AX regM__i16 (.D(det_q4_28[15]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i16.GSR = "ENABLED";
    FD1P3AX regM__i17 (.D(det_q4_28[16]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i17.GSR = "ENABLED";
    FD1P3AX regM__i18 (.D(det_q4_28[17]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i18.GSR = "ENABLED";
    FD1P3AX regM__i19 (.D(det_q4_28[18]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i19.GSR = "ENABLED";
    FD1P3AX regM__i20 (.D(det_q4_28[19]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i20.GSR = "ENABLED";
    FD1P3AX regM__i21 (.D(det_q4_28[20]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i21.GSR = "ENABLED";
    FD1P3AX regM__i22 (.D(det_q4_28[21]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i22.GSR = "ENABLED";
    FD1P3AX regM__i23 (.D(det_q4_28[22]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i23.GSR = "ENABLED";
    FD1P3AX regM__i24 (.D(det_q4_28[23]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i24.GSR = "ENABLED";
    FD1P3AX regM__i25 (.D(det_q4_28[24]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i25.GSR = "ENABLED";
    FD1P3AX regM__i26 (.D(det_q4_28[25]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i26.GSR = "ENABLED";
    FD1P3AX regM__i27 (.D(det_q4_28[26]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i27.GSR = "ENABLED";
    FD1P3AX regM__i28 (.D(det_q4_28[27]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i28.GSR = "ENABLED";
    FD1P3AX regM__i29 (.D(det_q4_28[28]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i29.GSR = "ENABLED";
    FD1P3AX regM__i30 (.D(det_q4_28[29]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i30.GSR = "ENABLED";
    FD1P3AX regM__i31 (.D(det_q4_28[30]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i31.GSR = "ENABLED";
    FD1P3AX regM__i32 (.D(det_q4_28[31]), .SP(clk_c_enable_239), .CK(clk_c), 
            .Q(regM[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regM__i32.GSR = "ENABLED";
    FD1S3AX regQ_i1 (.D(quotient_31__N_908[1]), .CK(clk_c), .Q(inv_det[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i1.GSR = "ENABLED";
    FD1S3AX regQ_i2 (.D(quotient_31__N_908[2]), .CK(clk_c), .Q(inv_det[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i2.GSR = "ENABLED";
    FD1S3AX regQ_i3 (.D(quotient_31__N_908[3]), .CK(clk_c), .Q(inv_det[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i3.GSR = "ENABLED";
    FD1S3AX regQ_i4 (.D(quotient_31__N_908[4]), .CK(clk_c), .Q(inv_det[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i4.GSR = "ENABLED";
    FD1S3AX regQ_i5 (.D(quotient_31__N_908[5]), .CK(clk_c), .Q(inv_det[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i5.GSR = "ENABLED";
    FD1S3AX regQ_i6 (.D(quotient_31__N_908[6]), .CK(clk_c), .Q(inv_det[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i6.GSR = "ENABLED";
    FD1S3AX regQ_i7 (.D(quotient_31__N_908[7]), .CK(clk_c), .Q(inv_det[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i7.GSR = "ENABLED";
    FD1S3AX regQ_i8 (.D(quotient_31__N_908[8]), .CK(clk_c), .Q(inv_det[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i8.GSR = "ENABLED";
    FD1S3AX regQ_i9 (.D(quotient_31__N_908[9]), .CK(clk_c), .Q(inv_det[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i9.GSR = "ENABLED";
    FD1S3AX regQ_i10 (.D(quotient_31__N_908[10]), .CK(clk_c), .Q(inv_det[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i10.GSR = "ENABLED";
    FD1S3AX regQ_i11 (.D(quotient_31__N_908[11]), .CK(clk_c), .Q(inv_det[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i11.GSR = "ENABLED";
    FD1S3AX regQ_i12 (.D(quotient_31__N_908[12]), .CK(clk_c), .Q(inv_det[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i12.GSR = "ENABLED";
    FD1S3AX regQ_i13 (.D(quotient_31__N_908[13]), .CK(clk_c), .Q(inv_det[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i13.GSR = "ENABLED";
    FD1S3AX regQ_i14 (.D(quotient_31__N_908[14]), .CK(clk_c), .Q(inv_det[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i14.GSR = "ENABLED";
    FD1S3AX regQ_i15 (.D(quotient_31__N_908[15]), .CK(clk_c), .Q(inv_det[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i15.GSR = "ENABLED";
    FD1S3AX regQ_i16 (.D(quotient_31__N_908[16]), .CK(clk_c), .Q(inv_det[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i16.GSR = "ENABLED";
    FD1S3AX regQ_i17 (.D(quotient_31__N_908[17]), .CK(clk_c), .Q(inv_det[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i17.GSR = "ENABLED";
    FD1S3AX regQ_i18 (.D(quotient_31__N_908[18]), .CK(clk_c), .Q(inv_det[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i18.GSR = "ENABLED";
    FD1S3AX regQ_i19 (.D(quotient_31__N_908[19]), .CK(clk_c), .Q(inv_det[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i19.GSR = "ENABLED";
    FD1S3AX regQ_i20 (.D(quotient_31__N_908[20]), .CK(clk_c), .Q(inv_det[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i20.GSR = "ENABLED";
    FD1S3AX regQ_i21 (.D(quotient_31__N_908[21]), .CK(clk_c), .Q(inv_det[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i21.GSR = "ENABLED";
    FD1S3AX regQ_i22 (.D(quotient_31__N_908[22]), .CK(clk_c), .Q(inv_det[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i22.GSR = "ENABLED";
    FD1S3AX regQ_i23 (.D(quotient_31__N_908[23]), .CK(clk_c), .Q(inv_det[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i23.GSR = "ENABLED";
    FD1S3AX regQ_i24 (.D(quotient_31__N_908[24]), .CK(clk_c), .Q(inv_det[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i24.GSR = "ENABLED";
    FD1S3AX regQ_i25 (.D(quotient_31__N_908[25]), .CK(clk_c), .Q(inv_det[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i25.GSR = "ENABLED";
    FD1S3AX regQ_i26 (.D(quotient_31__N_908[26]), .CK(clk_c), .Q(inv_det[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i26.GSR = "ENABLED";
    FD1S3AX regQ_i27 (.D(quotient_31__N_908[27]), .CK(clk_c), .Q(inv_det[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i27.GSR = "ENABLED";
    FD1S3AX regQ_i28 (.D(quotient_31__N_908[28]), .CK(clk_c), .Q(inv_det[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i28.GSR = "ENABLED";
    FD1S3AX regQ_i29 (.D(quotient_31__N_908[29]), .CK(clk_c), .Q(inv_det[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i29.GSR = "ENABLED";
    FD1S3AX regQ_i30 (.D(quotient_31__N_908[30]), .CK(clk_c), .Q(inv_det[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i30.GSR = "ENABLED";
    FD1S3AX regQ_i31 (.D(quotient_31__N_908[31]), .CK(clk_c), .Q(inv_det[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam regQ_i31.GSR = "ENABLED";
    LUT4 i781_2_lut (.A(regA[26]), .B(n3858[2]), .Z(n4577[27])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i781_2_lut.init = 16'h8888;
    LUT4 i542_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[8]), .Z(n7881)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i542_2_lut_3_lut.init = 16'he1e1;
    LUT4 i786_2_lut (.A(regA[31]), .B(n3858[2]), .Z(n4577[32])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i786_2_lut.init = 16'h8888;
    LUT4 i784_2_lut (.A(regA[29]), .B(n3858[2]), .Z(n4577[30])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i784_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_6 (.A(n8528), .B(n8399), .C(n3861), .D(n8448), 
         .Z(n8429)) /* synthesis lut_function=(A+(B (C)+!B !((D)+!C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i1_4_lut_adj_6.init = 16'heafa;
    LUT4 i228_2_lut (.A(\proximo_estado_2__N_952[0] ), .B(n3858[0]), .Z(n3883)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i228_2_lut.init = 16'h8888;
    LUT4 i785_2_lut (.A(regA[30]), .B(n3858[2]), .Z(n4577[31])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i785_2_lut.init = 16'h8888;
    LUT4 i778_2_lut (.A(regA[23]), .B(n3858[2]), .Z(n4577[24])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i778_2_lut.init = 16'h8888;
    LUT4 i6_2_lut (.A(det_q4_28[20]), .B(det_q4_28[19]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i550_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[12]), .Z(n7889)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i550_2_lut_3_lut.init = 16'he1e1;
    LUT4 i779_2_lut (.A(regA[24]), .B(n3858[2]), .Z(n4577[25])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i779_2_lut.init = 16'h8888;
    LUT4 i20_4_lut (.A(det_q4_28[5]), .B(det_q4_28[6]), .C(det_q4_28[7]), 
         .D(det_q4_28[22]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(det_q4_28[11]), .B(det_q4_28[18]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(det_q4_28[21]), .B(det_q4_28[2]), .C(det_q4_28[16]), 
         .D(det_q4_28[28]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(det_q4_28[17]), .B(det_q4_28[1]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(det_q4_28[9]), .B(det_q4_28[26]), .C(det_q4_28[12]), 
         .D(det_q4_28[4]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i28_4_lut (.A(det_q4_28[24]), .B(n56), .C(n46), .D(det_q4_28[8]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i617_4_lut (.A(inv_det[16]), .B(inv_det[17]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i617_4_lut.init = 16'hcac0;
    LUT4 i1149_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n8033)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i1149_4_lut.init = 16'h0001;
    LUT4 i9_2_lut (.A(det_q4_28[14]), .B(det_q4_28[30]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(det_q4_28[0]), .B(det_q4_28[10]), .C(det_q4_28[27]), 
         .D(det_q4_28[29]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i17_4_lut.init = 16'hfffe;
    FD1S3IX estado_atual_FSM_i1 (.D(n3883), .CK(clk_c), .CD(n8033), .Q(clk_c_enable_239));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i1.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(det_q4_28[13]), .B(n52), .C(n38), .D(det_q4_28[23]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i26_4_lut.init = 16'hfffe;
    PFUMX i1200 (.BLUT(n8728), .ALUT(n8729), .C0(n3861), .Z(quotient_31__N_908[16]));
    LUT4 i18_4_lut (.A(det_q4_28[3]), .B(det_q4_28[31]), .C(det_q4_28[15]), 
         .D(det_q4_28[25]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(42[8:21])
    defparam i18_4_lut.init = 16'hfffe;
    FD1S3IX estado_atual_FSM_i2 (.D(n8406), .CK(clk_c), .CD(n8033), .Q(n3858[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i2.GSR = "ENABLED";
    FD1S3IX estado_atual_FSM_i3 (.D(n3887), .CK(clk_c), .CD(n8033), .Q(n3863));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i3.GSR = "ENABLED";
    FD1S3IX estado_atual_FSM_i4 (.D(n3888), .CK(clk_c), .CD(n8033), .Q(n3858[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i4.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_7 (.A(n8550), .B(n8526), .C(i[1]), .D(i[4]), .Z(n8528)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i1_4_lut_adj_7.init = 16'hccce;
    FD1S3IX estado_atual_FSM_i6 (.D(n3892), .CK(clk_c), .CD(n8033), .Q(n3860));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i6.GSR = "ENABLED";
    FD1S3IX estado_atual_FSM_i7 (.D(n8452), .CK(clk_c), .CD(n8033), .Q(n3859));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_8 (.A(i[5]), .B(n7), .C(n8726), .D(n8532), .Z(n8399)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_8.init = 16'ha8aa;
    CCU2C i_418_add_4_7 (.A0(i[5]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n8297), 
          .S0(n29[5]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418_add_4_7.INIT0 = 16'haaa0;
    defparam i_418_add_4_7.INIT1 = 16'h0000;
    defparam i_418_add_4_7.INJECT1_0 = "NO";
    defparam i_418_add_4_7.INJECT1_1 = "NO";
    CCU2C i_418_add_4_5 (.A0(i[3]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n8296), 
          .COUT(n8297), .S0(n29[3]), .S1(n29[4]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418_add_4_5.INIT0 = 16'haaa0;
    defparam i_418_add_4_5.INIT1 = 16'haaa0;
    defparam i_418_add_4_5.INJECT1_0 = "NO";
    defparam i_418_add_4_5.INJECT1_1 = "NO";
    CCU2C i_418_add_4_3 (.A0(i[1]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n8295), 
          .COUT(n8296), .S0(n29[1]), .S1(n29[2]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418_add_4_3.INIT0 = 16'haaa0;
    defparam i_418_add_4_3.INIT1 = 16'haaa0;
    defparam i_418_add_4_3.INJECT1_0 = "NO";
    defparam i_418_add_4_3.INJECT1_1 = "NO";
    CCU2C i_418_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .COUT(n8295), 
          .S1(n29[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418_add_4_1.INIT0 = 16'h0000;
    defparam i_418_add_4_1.INIT1 = 16'h555f;
    defparam i_418_add_4_1.INJECT1_0 = "NO";
    defparam i_418_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_9 (.A(i[2]), .B(n8568), .C(n3858[2]), .D(i[5]), 
         .Z(n8550)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_9.init = 16'h1000;
    LUT4 i1_3_lut_adj_10 (.A(n3858[0]), .B(n3859), .C(\proximo_estado_2__N_952[0] ), 
         .Z(n8526)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i1_3_lut_adj_10.init = 16'hcece;
    LUT4 i1105_2_lut (.A(i[0]), .B(i[3]), .Z(n8568)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1105_2_lut.init = 16'heeee;
    FD1S3JX estado_atual_FSM_i0 (.D(n8429), .CK(clk_c), .PD(n8033), .Q(n3858[0]));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i0.GSR = "ENABLED";
    FD1P3IX i_418__i5 (.D(n29[5]), .SP(clk_c_enable_417), .CD(n8034), 
            .CK(clk_c), .Q(i[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418__i5.GSR = "ENABLED";
    FD1P3IX i_418__i4 (.D(n29[4]), .SP(clk_c_enable_417), .CD(n8034), 
            .CK(clk_c), .Q(i[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418__i4.GSR = "ENABLED";
    FD1P3IX i_418__i3 (.D(n29[3]), .SP(clk_c_enable_417), .CD(n8034), 
            .CK(clk_c), .Q(i[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418__i3.GSR = "ENABLED";
    FD1P3IX i_418__i2 (.D(n29[2]), .SP(clk_c_enable_417), .CD(n8034), 
            .CK(clk_c), .Q(i[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418__i2.GSR = "ENABLED";
    FD1P3IX i_418__i1 (.D(n29[1]), .SP(clk_c_enable_417), .CD(n8034), 
            .CK(clk_c), .Q(i[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418__i1.GSR = "ENABLED";
    FD1P3IX i_418__i0 (.D(n29[0]), .SP(clk_c_enable_417), .CD(n8034), 
            .CK(clk_c), .Q(i[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i_418__i0.GSR = "ENABLED";
    LUT4 i696_2_lut (.A(clk_c_enable_239), .B(n3858[2]), .Z(n8034)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(116[26:27])
    defparam i696_2_lut.init = 16'h2222;
    LUT4 i754_2_lut (.A(regA[32]), .B(n3861), .Z(A0_N_1113)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i754_2_lut.init = 16'h8888;
    LUT4 i619_4_lut (.A(inv_det[17]), .B(inv_det[18]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i619_4_lut.init = 16'hcac0;
    LUT4 i621_4_lut (.A(inv_det[18]), .B(inv_det[19]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i621_4_lut.init = 16'hcac0;
    LUT4 i623_4_lut (.A(inv_det[19]), .B(inv_det[20]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i623_4_lut.init = 16'hcac0;
    LUT4 i625_4_lut (.A(inv_det[20]), .B(inv_det[21]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i625_4_lut.init = 16'hcac0;
    LUT4 i627_4_lut (.A(inv_det[21]), .B(inv_det[22]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i627_4_lut.init = 16'hcac0;
    LUT4 i629_4_lut (.A(inv_det[22]), .B(inv_det[23]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i629_4_lut.init = 16'hcac0;
    LUT4 i631_4_lut (.A(inv_det[23]), .B(inv_det[24]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i631_4_lut.init = 16'hcac0;
    LUT4 i633_4_lut (.A(inv_det[24]), .B(inv_det[25]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i633_4_lut.init = 16'hcac0;
    LUT4 i635_4_lut (.A(inv_det[25]), .B(inv_det[26]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i635_4_lut.init = 16'hcac0;
    LUT4 i637_4_lut (.A(inv_det[26]), .B(inv_det[27]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i637_4_lut.init = 16'hcac0;
    LUT4 i639_4_lut (.A(inv_det[27]), .B(inv_det[28]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i639_4_lut.init = 16'hcac0;
    LUT4 i641_4_lut (.A(inv_det[28]), .B(inv_det[29]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i641_4_lut.init = 16'hcac0;
    LUT4 i643_4_lut (.A(inv_det[29]), .B(inv_det[30]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i643_4_lut.init = 16'hcac0;
    LUT4 i645_4_lut (.A(inv_det[30]), .B(inv_det[31]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i645_4_lut.init = 16'hcac0;
    LUT4 i1152_3_lut (.A(n3858[0]), .B(n3861), .C(n3858[4]), .Z(clk_c_enable_192)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i1152_3_lut.init = 16'h0101;
    LUT4 i566_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[28]), .Z(n7905)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i566_2_lut_3_lut.init = 16'he1e1;
    LUT4 i581_4_lut (.A(n8524), .B(regA[32]), .C(n3861), .D(n3858[2]), 
         .Z(quotient_31__N_908[0])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i581_4_lut.init = 16'h303a;
    LUT4 i1_2_lut (.A(clk_c_enable_239), .B(inv_det[0]), .Z(n8524)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i585_4_lut (.A(inv_det[0]), .B(inv_det[1]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i585_4_lut.init = 16'hcac0;
    LUT4 i587_4_lut (.A(inv_det[1]), .B(inv_det[2]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i587_4_lut.init = 16'hcac0;
    LUT4 i589_4_lut (.A(inv_det[2]), .B(inv_det[3]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i589_4_lut.init = 16'hcac0;
    LUT4 i591_4_lut (.A(inv_det[3]), .B(inv_det[4]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i591_4_lut.init = 16'hcac0;
    LUT4 i593_4_lut (.A(inv_det[4]), .B(inv_det[5]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i593_4_lut.init = 16'hcac0;
    LUT4 i595_4_lut (.A(inv_det[5]), .B(inv_det[6]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i595_4_lut.init = 16'hcac0;
    LUT4 i597_4_lut (.A(inv_det[6]), .B(inv_det[7]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i597_4_lut.init = 16'hcac0;
    LUT4 i599_4_lut (.A(inv_det[7]), .B(inv_det[8]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i599_4_lut.init = 16'hcac0;
    LUT4 i601_4_lut (.A(inv_det[8]), .B(inv_det[9]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i601_4_lut.init = 16'hcac0;
    LUT4 i603_4_lut (.A(inv_det[9]), .B(inv_det[10]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i603_4_lut.init = 16'hcac0;
    LUT4 i530_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[2]), .Z(n7869)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i530_2_lut_3_lut.init = 16'he1e1;
    LUT4 i532_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[3]), .Z(n7871)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i532_2_lut_3_lut.init = 16'he1e1;
    LUT4 i554_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[22]), .Z(n7893)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i554_2_lut_3_lut.init = 16'he1e1;
    LUT4 i1_4_lut_adj_11 (.A(n3859), .B(n3858[0]), .C(n8448), .D(n3861), 
         .Z(clk_c_enable_11)) /* synthesis lut_function=(A+!(B (C (D))+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_11.init = 16'hafee;
    LUT4 i261_2_lut (.A(n3861), .B(n3859), .Z(ready_N_1109)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i261_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_12 (.A(n8562), .B(n7), .C(regA[32]), .D(i[1]), 
         .Z(n8448)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(129[10:21])
    defparam i1_4_lut_adj_12.init = 16'hfffe;
    LUT4 i556_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[23]), .Z(n7895)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i556_2_lut_3_lut.init = 16'he1e1;
    LUT4 i568_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[29]), .Z(n7907)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i568_2_lut_3_lut.init = 16'he1e1;
    LUT4 i522_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[20]), .Z(n7861)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i522_2_lut_3_lut.init = 16'he1e1;
    LUT4 i605_4_lut (.A(inv_det[10]), .B(inv_det[11]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i605_4_lut.init = 16'hcac0;
    FD1S3AX estado_atual_FSM_i5 (.D(n8040), .CK(clk_c), .Q(n3861));   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam estado_atual_FSM_i5.GSR = "ENABLED";
    FD1P3AX A0_63 (.D(A0_N_1113), .SP(clk_c_enable_432), .CK(clk_c), .Q(proximo_estado_2__N_946[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=56, LSE_RLINE=64 */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(96[9] 140[16])
    defparam A0_63.GSR = "DISABLED";
    LUT4 i524_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[21]), .Z(n7863)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i524_2_lut_3_lut.init = 16'he1e1;
    LUT4 i518_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[18]), .Z(n7857)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i518_2_lut_3_lut.init = 16'he1e1;
    LUT4 i1_2_lut_adj_13 (.A(i[2]), .B(i[0]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(129[10:21])
    defparam i1_2_lut_adj_13.init = 16'heeee;
    LUT4 i520_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[19]), .Z(n7859)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i520_2_lut_3_lut.init = 16'he1e1;
    LUT4 i780_2_lut (.A(regA[25]), .B(n3858[2]), .Z(n4577[26])) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i780_2_lut.init = 16'h8888;
    LUT4 i562_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[26]), .Z(n7901)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i562_2_lut_3_lut.init = 16'he1e1;
    LUT4 i607_4_lut (.A(inv_det[11]), .B(inv_det[12]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i607_4_lut.init = 16'hcac0;
    LUT4 i514_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[16]), .Z(n7853)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i514_2_lut_3_lut.init = 16'he1e1;
    LUT4 i609_4_lut (.A(inv_det[12]), .B(inv_det[13]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i609_4_lut.init = 16'hcac0;
    LUT4 i516_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[17]), .Z(n7855)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i516_2_lut_3_lut.init = 16'he1e1;
    LUT4 i564_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[27]), .Z(n7903)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i564_2_lut_3_lut.init = 16'he1e1;
    LUT4 i611_4_lut (.A(inv_det[13]), .B(inv_det[14]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i611_4_lut.init = 16'hcac0;
    LUT4 i510_2_lut_3_lut (.A(n3859), .B(n3860), .C(regM[14]), .Z(n7849)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(103[13] 139[22])
    defparam i510_2_lut_3_lut.init = 16'he1e1;
    LUT4 i613_4_lut (.A(inv_det[14]), .B(inv_det[15]), .C(n8723), .D(n3858[2]), 
         .Z(quotient_31__N_908[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/projeto_final/kalman_core/divnrda_fsm.vhd(51[9] 90[18])
    defparam i613_4_lut.init = 16'hcac0;
    
endmodule
