// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Fri Sep 26 14:45:07 2025
//
// Verilog Description of module backward
//

module backward (clk, rst, start, U_in, y_in, done, x_out) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(4[8:16])
    input clk;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(5[24:27])
    input rst;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    input start;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(7[24:29])
    input [511:0]U_in;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    input [127:0]y_in;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    output done;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(12[24:28])
    output [127:0]x_out;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    
    wire clk_c /* synthesis is_clock=1, SET_AS_NETWORK=clk_c */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(5[24:27])
    
    wire GND_net, VCC_net, rst_c, start_c, U_in_c_511, U_in_c_510, 
        U_in_c_509, U_in_c_508, U_in_c_507, U_in_c_506, U_in_c_505, 
        U_in_c_504, U_in_c_503, U_in_c_502, U_in_c_501, U_in_c_500, 
        U_in_c_499, U_in_c_498, U_in_c_497, U_in_c_496, U_in_c_495, 
        U_in_c_494, U_in_c_493, U_in_c_492, U_in_c_491, U_in_c_490, 
        U_in_c_489, U_in_c_488, U_in_c_487, U_in_c_486, U_in_c_485, 
        U_in_c_484, U_in_c_483, U_in_c_482, U_in_c_481, U_in_c_480, 
        U_in_c_479, U_in_c_478, U_in_c_477, U_in_c_476, U_in_c_475, 
        U_in_c_474, U_in_c_473, U_in_c_472, U_in_c_471, U_in_c_470, 
        U_in_c_469, U_in_c_468, U_in_c_467, U_in_c_466, U_in_c_465, 
        U_in_c_464, U_in_c_463, U_in_c_462, U_in_c_461, U_in_c_460, 
        U_in_c_459, U_in_c_458, U_in_c_457, U_in_c_456, U_in_c_455, 
        U_in_c_454, U_in_c_453, U_in_c_452, U_in_c_451, U_in_c_450, 
        U_in_c_449, U_in_c_448, U_in_c_447, U_in_c_446, U_in_c_445, 
        U_in_c_444, U_in_c_443, U_in_c_442, U_in_c_441, U_in_c_440, 
        U_in_c_439, U_in_c_438, U_in_c_437, U_in_c_436, U_in_c_435, 
        U_in_c_434, U_in_c_433, U_in_c_432, U_in_c_431, U_in_c_430, 
        U_in_c_429, U_in_c_428, U_in_c_427, U_in_c_426, U_in_c_425, 
        U_in_c_424, U_in_c_423, U_in_c_422, U_in_c_421, U_in_c_420, 
        U_in_c_419, U_in_c_418, U_in_c_417, U_in_c_416, U_in_c_415, 
        U_in_c_414, U_in_c_413, U_in_c_412, U_in_c_411, U_in_c_410, 
        U_in_c_409, U_in_c_408, U_in_c_407, U_in_c_406, U_in_c_405, 
        U_in_c_404, U_in_c_403, U_in_c_402, U_in_c_401, U_in_c_400, 
        U_in_c_399, U_in_c_398, U_in_c_397, U_in_c_396, U_in_c_395, 
        U_in_c_394, U_in_c_393, U_in_c_392, U_in_c_391, U_in_c_390, 
        U_in_c_389, U_in_c_388, U_in_c_387, U_in_c_386, U_in_c_385, 
        U_in_c_384, U_in_c_383, U_in_c_382, U_in_c_381, U_in_c_380, 
        U_in_c_379, U_in_c_378, U_in_c_377, U_in_c_376, U_in_c_375, 
        U_in_c_374, U_in_c_373, U_in_c_372, U_in_c_371, U_in_c_370, 
        U_in_c_369, U_in_c_368, U_in_c_367, U_in_c_366, U_in_c_365, 
        U_in_c_364, U_in_c_363, U_in_c_362, U_in_c_361, U_in_c_360, 
        U_in_c_359, U_in_c_358, U_in_c_357, U_in_c_356, U_in_c_355, 
        U_in_c_354, U_in_c_353, U_in_c_352, U_in_c_351, U_in_c_350, 
        U_in_c_349, U_in_c_348, U_in_c_347, U_in_c_346, U_in_c_345, 
        U_in_c_344, U_in_c_343, U_in_c_342, U_in_c_341, U_in_c_340, 
        U_in_c_339, U_in_c_338, U_in_c_337, U_in_c_336, U_in_c_335, 
        U_in_c_334, U_in_c_333, U_in_c_332, U_in_c_331, U_in_c_330, 
        U_in_c_329, U_in_c_328, U_in_c_327, U_in_c_326, U_in_c_325, 
        U_in_c_324, U_in_c_323, U_in_c_322, U_in_c_321, U_in_c_320, 
        U_in_c_319, U_in_c_318, U_in_c_317, U_in_c_316, U_in_c_315, 
        U_in_c_314, U_in_c_313, U_in_c_312, U_in_c_311, U_in_c_310, 
        U_in_c_309, U_in_c_308, U_in_c_307, U_in_c_306, U_in_c_305, 
        U_in_c_304, U_in_c_303, U_in_c_302, U_in_c_301, U_in_c_300, 
        U_in_c_299, U_in_c_298, U_in_c_297, U_in_c_296, U_in_c_295, 
        U_in_c_294, U_in_c_293, U_in_c_292, U_in_c_291, U_in_c_290, 
        U_in_c_289, U_in_c_288, U_in_c_287, U_in_c_286, U_in_c_285, 
        U_in_c_284, U_in_c_283, U_in_c_282, U_in_c_281, U_in_c_280, 
        U_in_c_279, U_in_c_278, U_in_c_277, U_in_c_276, U_in_c_275, 
        U_in_c_274, U_in_c_273, U_in_c_272, U_in_c_271, U_in_c_270, 
        U_in_c_269, U_in_c_268, U_in_c_267, U_in_c_266, U_in_c_265, 
        U_in_c_264, U_in_c_263, U_in_c_262, U_in_c_261, U_in_c_260, 
        U_in_c_259, U_in_c_258, U_in_c_257, U_in_c_256, U_in_c_255, 
        U_in_c_254, U_in_c_253, U_in_c_252, U_in_c_251, U_in_c_250, 
        U_in_c_249, U_in_c_248, U_in_c_247, U_in_c_246, U_in_c_245, 
        U_in_c_244, U_in_c_243, U_in_c_242, U_in_c_241, U_in_c_240, 
        U_in_c_239, U_in_c_238, U_in_c_237, U_in_c_236, U_in_c_235, 
        U_in_c_234, U_in_c_233, U_in_c_232, U_in_c_231, U_in_c_230, 
        U_in_c_229, U_in_c_228, U_in_c_227, U_in_c_226, U_in_c_225, 
        U_in_c_224, U_in_c_223, U_in_c_222, U_in_c_221, U_in_c_220, 
        U_in_c_219, U_in_c_218, U_in_c_217, U_in_c_216, U_in_c_215, 
        U_in_c_214, U_in_c_213, U_in_c_212, U_in_c_211, U_in_c_210, 
        U_in_c_209, U_in_c_208, U_in_c_207, U_in_c_206, U_in_c_205, 
        U_in_c_204, U_in_c_203, U_in_c_202, U_in_c_201, U_in_c_200, 
        U_in_c_199, U_in_c_198, U_in_c_197, U_in_c_196, U_in_c_195, 
        U_in_c_194, U_in_c_193, U_in_c_192, U_in_c_191, U_in_c_190, 
        U_in_c_189, U_in_c_188, U_in_c_187, U_in_c_186, U_in_c_185, 
        U_in_c_184, U_in_c_183, U_in_c_182, U_in_c_181, U_in_c_180, 
        U_in_c_179, U_in_c_178, U_in_c_177, U_in_c_176, U_in_c_175, 
        U_in_c_174, U_in_c_173, U_in_c_172, U_in_c_171, U_in_c_170, 
        U_in_c_169, U_in_c_168, U_in_c_167, U_in_c_166, U_in_c_165, 
        U_in_c_164, U_in_c_163, U_in_c_162, U_in_c_161, U_in_c_160, 
        U_in_c_159, U_in_c_158, U_in_c_157, U_in_c_156, U_in_c_155, 
        U_in_c_154, U_in_c_153, U_in_c_152, U_in_c_151, U_in_c_150, 
        U_in_c_149, U_in_c_148, U_in_c_147, U_in_c_146, U_in_c_145, 
        U_in_c_144, U_in_c_143, U_in_c_142, U_in_c_141, U_in_c_140, 
        U_in_c_139, U_in_c_138, U_in_c_137, U_in_c_136, U_in_c_135, 
        U_in_c_134, U_in_c_133, U_in_c_132, U_in_c_131, U_in_c_130, 
        U_in_c_129, U_in_c_128, U_in_c_127, U_in_c_126, U_in_c_125, 
        U_in_c_124, U_in_c_123, U_in_c_122, U_in_c_121, U_in_c_120, 
        U_in_c_119, U_in_c_118, U_in_c_117, U_in_c_116, U_in_c_115, 
        U_in_c_114, U_in_c_113, U_in_c_112, U_in_c_111, U_in_c_110, 
        U_in_c_109, U_in_c_108, U_in_c_107, U_in_c_106, U_in_c_105, 
        U_in_c_104, U_in_c_103, U_in_c_102, U_in_c_101, U_in_c_100, 
        U_in_c_99, U_in_c_98, U_in_c_97, U_in_c_96, U_in_c_95, U_in_c_94, 
        U_in_c_93, U_in_c_92, U_in_c_91, U_in_c_90, U_in_c_89, U_in_c_88, 
        U_in_c_87, U_in_c_86, U_in_c_85, U_in_c_84, U_in_c_83, U_in_c_82, 
        U_in_c_81, U_in_c_80, U_in_c_79, U_in_c_78, U_in_c_77, U_in_c_76, 
        U_in_c_75, U_in_c_74, U_in_c_73, U_in_c_72, U_in_c_71, U_in_c_70, 
        U_in_c_69, U_in_c_68, U_in_c_67, U_in_c_66, U_in_c_65, U_in_c_64, 
        U_in_c_63, U_in_c_62, U_in_c_61, U_in_c_60, U_in_c_59, U_in_c_58, 
        U_in_c_57, U_in_c_56, U_in_c_55, U_in_c_54, U_in_c_53, U_in_c_52, 
        U_in_c_51, U_in_c_50, U_in_c_49, U_in_c_48, U_in_c_47, U_in_c_46, 
        U_in_c_45, U_in_c_44, U_in_c_43, U_in_c_42, U_in_c_41, U_in_c_40, 
        U_in_c_39, U_in_c_38, U_in_c_37, U_in_c_36, U_in_c_35, U_in_c_34, 
        U_in_c_33, U_in_c_32, U_in_c_31, U_in_c_30, U_in_c_29, U_in_c_28, 
        U_in_c_27, U_in_c_26, U_in_c_25, U_in_c_24, U_in_c_23, U_in_c_22, 
        U_in_c_21, U_in_c_20, U_in_c_19, U_in_c_18, U_in_c_17, U_in_c_16, 
        U_in_c_15, U_in_c_14, U_in_c_13, U_in_c_12, U_in_c_11, U_in_c_10, 
        U_in_c_9, U_in_c_8, U_in_c_7, U_in_c_6, U_in_c_5, U_in_c_4, 
        U_in_c_3, U_in_c_2, U_in_c_1, U_in_c_0, y_in_c_127, y_in_c_126, 
        y_in_c_125, y_in_c_124, y_in_c_123, y_in_c_122, y_in_c_121, 
        y_in_c_120, y_in_c_119, y_in_c_118, y_in_c_117, y_in_c_116, 
        y_in_c_115, y_in_c_114, y_in_c_113, y_in_c_112, y_in_c_111, 
        y_in_c_110, y_in_c_109, y_in_c_108, y_in_c_107, y_in_c_106, 
        y_in_c_105, y_in_c_104, y_in_c_103, y_in_c_102, y_in_c_101, 
        y_in_c_100, y_in_c_99, y_in_c_98, y_in_c_97, y_in_c_96, y_in_c_95, 
        y_in_c_94, y_in_c_93, y_in_c_92, y_in_c_91, y_in_c_90, y_in_c_89, 
        y_in_c_88, y_in_c_87, y_in_c_86, y_in_c_85, y_in_c_84, y_in_c_83, 
        y_in_c_82, y_in_c_81, y_in_c_80, y_in_c_79, y_in_c_78, y_in_c_77, 
        y_in_c_76, y_in_c_75, y_in_c_74, y_in_c_73, y_in_c_72, y_in_c_71, 
        y_in_c_70, y_in_c_69, y_in_c_68, y_in_c_67, y_in_c_66, y_in_c_65, 
        y_in_c_64, y_in_c_63, y_in_c_62, y_in_c_61, y_in_c_60, y_in_c_59, 
        y_in_c_58, y_in_c_57, y_in_c_56, y_in_c_55, y_in_c_54, y_in_c_53, 
        y_in_c_52, y_in_c_51, y_in_c_50, y_in_c_49, y_in_c_48, y_in_c_47, 
        y_in_c_46, y_in_c_45, y_in_c_44, y_in_c_43, y_in_c_42, y_in_c_41, 
        y_in_c_40, y_in_c_39, y_in_c_38, y_in_c_37, y_in_c_36, y_in_c_35, 
        y_in_c_34, y_in_c_33, y_in_c_32, y_in_c_31, y_in_c_30, y_in_c_29, 
        y_in_c_28, y_in_c_27, y_in_c_26, y_in_c_25, y_in_c_24, y_in_c_23, 
        y_in_c_22, y_in_c_21, y_in_c_20, y_in_c_19, y_in_c_18, y_in_c_17, 
        y_in_c_16, y_in_c_15, y_in_c_14, y_in_c_13, y_in_c_12, y_in_c_11, 
        y_in_c_10, y_in_c_9, y_in_c_8, y_in_c_7, y_in_c_6, y_in_c_5, 
        y_in_c_4, y_in_c_3, y_in_c_2, y_in_c_1, y_in_c_0, done_c, 
        x_out_c_127, x_out_c_126, x_out_c_125, x_out_c_124, x_out_c_123, 
        x_out_c_122, x_out_c_121, x_out_c_120, x_out_c_119, x_out_c_118, 
        x_out_c_117, x_out_c_116, x_out_c_115, x_out_c_114, x_out_c_113, 
        x_out_c_112, x_out_c_111, x_out_c_110, x_out_c_109, x_out_c_108, 
        x_out_c_107, x_out_c_106, x_out_c_105, x_out_c_104, x_out_c_103, 
        x_out_c_102, x_out_c_101, x_out_c_100, x_out_c_99, x_out_c_98, 
        x_out_c_97, x_out_c_96, x_out_c_95, x_out_c_94, x_out_c_93, 
        x_out_c_92, x_out_c_91, x_out_c_90, x_out_c_89, x_out_c_88, 
        x_out_c_87, x_out_c_86, x_out_c_85, x_out_c_84, x_out_c_83, 
        x_out_c_82, x_out_c_81, x_out_c_80, x_out_c_79, x_out_c_78, 
        x_out_c_77, x_out_c_76, x_out_c_75, x_out_c_74, x_out_c_73, 
        x_out_c_72, x_out_c_71, x_out_c_70, x_out_c_69, x_out_c_68, 
        x_out_c_67, x_out_c_66, x_out_c_65, x_out_c_64, x_out_c_63, 
        x_out_c_62, x_out_c_61, x_out_c_60, x_out_c_59, x_out_c_58, 
        x_out_c_57, x_out_c_56, x_out_c_55, x_out_c_54, x_out_c_53, 
        x_out_c_52, x_out_c_51, x_out_c_50, x_out_c_49, x_out_c_48, 
        x_out_c_47, x_out_c_46, x_out_c_45, x_out_c_44, x_out_c_43, 
        x_out_c_42, x_out_c_41, x_out_c_40, x_out_c_39, x_out_c_38, 
        x_out_c_37, x_out_c_36, x_out_c_35, x_out_c_34, x_out_c_33, 
        x_out_c_32, x_out_c_31, x_out_c_30, x_out_c_29, x_out_c_28, 
        x_out_c_27, x_out_c_26, x_out_c_25, x_out_c_24, x_out_c_23, 
        x_out_c_22, x_out_c_21, x_out_c_20, x_out_c_19, x_out_c_18, 
        x_out_c_17, x_out_c_16, x_out_c_15, x_out_c_14, x_out_c_13, 
        x_out_c_12, x_out_c_11, x_out_c_10, x_out_c_9, x_out_c_8, 
        x_out_c_7, x_out_c_6, x_out_c_5, x_out_c_4, x_out_c_3, x_out_c_2, 
        x_out_c_1, x_out_c_0;
    wire [31:0]\U[0] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[1] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[2] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[3] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[4] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[5] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[6] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[7] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[8] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[9] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[10] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[11] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[12] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[13] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[14] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    wire [31:0]\U[15] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(18[21:22])
    
    wire n42497, n39796, n39794, n42496;
    wire [31:0]\y[3] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(19[21:22])
    wire [31:0]\x[0] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(20[21:22])
    wire [31:0]\x[1] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(20[21:22])
    wire [31:0]\x[2] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(20[21:22])
    wire [31:0]\x[3] ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(20[21:22])
    wire [31:0]i;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(22[11:12])
    
    wire n20433, n38693, n39789, n42495, n18965, n38684, n31054, 
        n18720, n19277, n18719, n20383, n20392, n20393, n20394, 
        n20395, n20396, n20397, n20398, n18718, n18717, n19279, 
        n18716, n19278, n20391, n20384, n20385, n20386, n20387, 
        n20388, n20389, n20390, n37686, n18715, n19119, n18714, 
        n19280, n18713, n20399, n20376, n20377, n20378, n20379, 
        n20380, n20381, n20382, n18712, n31021, n18711, n19282, 
        n18710, n19281, n20343, n20368, n20369, n20370, n20371, 
        n20372, n20373, n20374, n39780, n42494, n38682, n37505, 
        n18709, n19114, n18708, n19283, n18707, n20351, n20360, 
        n20361, n20362, n20363, n20364, n20365, n20366, n38677, 
        n18954, n18706, n19285, n18705, n19284, n20359, n20352, 
        n20353, n20354, n20355, n20356, n20357, n20358, n18704, 
        n19109, n18703, n19286, n18702, n20367, n20344, n20345, 
        n20346, n20347, n20348, n20349, n20350, n42493, n18701, 
        n18700, n19288, n18699, n19287, n20311, n20336, n20337, 
        n20338, n20339, n20340, n20341, n20342, n18698, n193, 
        n19104, n18697, n19289, n18696, n20319, n20328, n20329, 
        n20330, n20331, n20332, n20333, n20334, n39773, n18695, 
        n188, n18592, n19291, n18694, n19290, n20327, n20320, 
        n20321, n20322, n20323, n20324, n20325, n20326, n18693, 
        n183, n18591, n18692, n19292, n18691, n20335, n20312, 
        n20313, n20314, n20315, n20316, n20317, n20318, n38668, 
        n19593, n18690, n178, n18590, n19294, n18689, n19293, 
        n20279, n20304, n20305, n20306, n20307, n20308, n20309, 
        n20310, n18688, n173, n18589, n18687, n19295, n18686, 
        n20287, n20296, n20297, n20298, n20299, n20300, n20301, 
        n20302, n18685, n168, n18588, n193_adj_1, n194, n19296, 
        n20295, n20288, n20289, n20290, n20291, n20292, n20293, 
        n20294, n18684, n163, n19097, n190, n191, n192, n20303, 
        n20280, n20281, n20282, n20283, n20284, n20285, n20286, 
        n18683, n18587, n18586, n187, n188_adj_2, n189, n20247, 
        n20272, n20273, n20274, n20275, n20276, n20277, n20278, 
        n19686, n18585, n18938, n184, n185, n186, n20255, n20264, 
        n20265, n20266, n20267, n20268, n20269, n20270, n18682, 
        n18584, n172, n181, n182, n183_adj_3, n20263, n20256, 
        n20257, n20258, n20259, n20260, n20261, n20262, n39760, 
        n19683, n18583, n178_adj_4, n178_adj_5, n179, n180, n20271, 
        n20248, n20249, n20250, n20251, n20252, n20253, n20254, 
        n38661, n18681, n18582, n184_adj_6, n175, n176, n177, 
        n20240, n20241, n20242, n20243, n20244, n20245, n20246, 
        n19680, n18581, n190_adj_7, n172_adj_8, n173_adj_9, n174, 
        n40592, n20238, n38655, n40591, n19677, n19009, n18976, 
        n169, n170, n171, n39756, n40590, n19675, n19070, n18975, 
        n166, n167, n168_adj_10, n20239, n163_adj_11, n19673, n19014, 
        n18974, n163_adj_12, n164, n165, n20183, n160, n157, n40589, 
        n19671, n19016, n18973, n18580, n18579, n18578, n20191, 
        n20200, n20201, n20202, n20203, n20204, n20205, n40588, 
        n40587, n40586, n39753, n19669, n19018, n19408, n18577, 
        n18576, n18575, n20199, n20192, n20193, n20194, n20195, 
        n20196, n20197, n20198, n19667, n19062, n18680, n18574, 
        n18573, n18572, n154, n20184, n20185, n20186, n20187, 
        n20188, n20189, n20190, n40585, n19664, n19021, n18679, 
        n18571, n18570, n18569, n20151, n20176, n20177, n20178, 
        n20179, n20180, n20181, n20182, n19661, n19059, n18678, 
        n18568, n18567, n18566, n20159, n20168, n20169, n20170, 
        n20171, n20172, n20173, n20174, n38644, n19658, n19057, 
        n18677, n18565, n18564, n18563, n20167, n20160, n20161, 
        n20162, n20163, n20164, n20165, n20166, n40584, n19655, 
        n19026, n18676, n18562, n18561, n18560, n20175, n20152, 
        n20153, n20154, n20155, n20156, n20157, n20158, n38641, 
        n40583, n19653, n19652, n19219, n19226, n18966, n18675, 
        n20075, n20103, n20090, n20125, n20080, n20078, n20102, 
        n20076, n39741, n19649, n19713, n18964, n19225, n18674, 
        n18963, n20081, n20101, n20089, n20123, n20050, n20074, 
        n20100, n20064, n40582, n19715, n19550, n19185, n19224, 
        n18673, n18961, n20071, n20098, n20088, n20121, n20047, 
        n20072, n20097, n20062, n19548, n19718, n19215, n19223, 
        n18672, n18959, n20069, n20095, n20087, n20119, n20044, 
        n20070, n20094, n20060, n19640, n19720, n19545, n19188, 
        n19222, n18671, n18957, n20067, n20092, n20086, n20117, 
        n20041, n20068, n20091, n20058, n40581, n40580, n19543, 
        n19723, n18670, n19221, n18955, n18669, n20073, n20079, 
        n20085, n20115, n20034, n20066, n20082, n20056, n40579, 
        n19540, n19726, n18953, n19220, n18668, n18952, n20035, 
        n20065, n20084, n20113, n20031, n20038, n20032, n20054, 
        n40577, n40576, n19538, n19728, n18667, n18950, n18666, 
        n18949, n20022, n20063, n20083, n20077, n20030, n19985, 
        n20025, n20052, n39733, n19536, n19730, n18665, n18947, 
        n18664, n18946, n20020, n20061, n20033, n20037, n20029, 
        n19979, n20023, n20049, n38629, n19733, n19532, n18663, 
        n18944, n18943, n18942, n20026, n20059, n20011, n20003, 
        n20028, n19978, n20021, n20046, n40575, n19679, n19526, 
        n191_adj_13, n192_adj_14, n193_adj_15, n20024, n20057, n20007, 
        n20000, n20027, n19977, n20019, n20043, n40574, n19681, 
        n19666, n185_adj_16, n186_adj_17, n187_adj_18, n20014, n20055, 
        n19990, n19997, n20010, n19976, n20017, n20040, n40573, 
        n39728, n18662, n19663, n179_adj_19, n180_adj_20, n181_adj_21, 
        n20004, n20053, n19962, n19994, n20006, n19975, n20015, 
        n20036, n38621, n40572, n19684, n19660, n173_adj_22, n174_adj_23, 
        n175_adj_24, n20018, n20051, n19960, n19988, n19991, n19974, 
        n20013, n19987, n18661, n19657, n168_adj_25, n169_adj_26, 
        n19089, n20016, n20048, n19958, n19984, n19947, n19973, 
        n20009, n19968, n37681, n19687, n18939, n163_adj_27, n164_adj_28, 
        n19092, n20008, n20045, n19956, n19983, n19936, n19969, 
        n20005, n19963, n40571, n40570, n38616, n19763, n19798, 
        n19651, n18937, n19992, n20042, n19950, n19982, n19935, 
        n19964, n20002, n19953, n40569, n19552, n19797, n19714, 
        n18936, n20001, n20039, n19946, n19981, n19934, n19961, 
        n19999, n19945, n40568, n19788, n19796, n19716, n19549, 
        n20012, n19986, n19944, n19980, n19933, n19959, n19996, 
        n19943, n40567, n40566, n40565, n19594, n19767, n19795, 
        n19547, n19719, n19995, n19971, n19942, n19970, n19932, 
        n19957, n19993, n19941, n19639, n19785, n19794, n19721, 
        n19544, n19911, n19966, n19940, n19965, n19931, n19955, 
        n19989, n19939, n40564, n19542, n19760, n19724, n19541, 
        n19922, n19952, n19938, n19954, n19930, n19951, n19949, 
        n19937, n40562, n18945, n19539, n19103, n19102, n19101, 
        n19998, n19923, n19924, n19925, n19926, n19927, n19928, 
        n19929, n40561, n18948, n19537, n19106, n18660, n19105, 
        n19948, n19912, n19913, n19914, n19915, n19916, n19917, 
        n19918, n18951, n19535, n18659, n19108, n18658, n19238, 
        n19901, n19902, n19903, n19904, n19905, n19906, n19907, 
        n39718, n18657, n19734, n19111, n18656, n19110, n19878, 
        n19890, n19891, n19892, n19893, n19894, n19895, n19896, 
        n40560, n40559, n40558, n36882, n39716, n19595, n18956, 
        n18920, n18655, n19113, n18654, n19889, n19879, n19880, 
        n19881, n19882, n19883, n19884, n19885, n39714, n40557, 
        n19638, n18958, n174_adj_29, n19116, n18653, n19115, n19900, 
        n19237, n19236, n19235, n19234, n19233, n39712, n40556, 
        n19596, n19637, n18960, n173_adj_30, n18652, n19118, n18651, 
        n19273, n19248, n19247, n19246, n19245, n19244, n19243, 
        n19242, n19597, n18962, n19121, n18650, n19120, n18649, 
        n19259, n19258, n19257, n19256, n19255, n19254, n19253, 
        n19636, n18648, n18647, n151, n18646, n19260, n19267, 
        n18645, n19266, n18644, n19265, n18643, n19264, n19598, 
        n18642, n19530, n18641, n19249, n18640, n19272, n18639, 
        n19271, n18638, n19270, n18637, n40555, n40554, n19635, 
        n19599, n19464, n19037, n19736, n19197, n19183, n19212, 
        n19176, n19207, n19206, n19218, n19205, n40553, n19634, 
        n19600, n19038, n19529, n19194, n19184, n19190, n19177, 
        n19160, n19204, n19217, n19167, n19633, n19601, n18999, 
        n19039, n19632, n19199, n19216, n19211, n19178, n19403, 
        n19203, n19186, n19166, n37339, n19602, n19468, n19040, 
        n19631, n19200, n19187, n19191, n19179, n19157, n19202, 
        n19214, n19165, n40552, n38597, n40551, n18996, n19457, 
        n19603, n19393, n19213, n19210, n19180, n19156, n19201, 
        n19189, n19164, n40550, n40549, n19630, n19604, n19629, 
        n19458, n19605, n19628, n19198, n19195, n19192, n19181, 
        n19409, n19168, n19208, n19163, n37338, n19606, n19459, 
        n19531, n19735, n148, n19394, n19209, n19182, n19155, 
        n19410, n19162, n40547, n39698, n19627, n37337, n40546, 
        n19731, n19534, n19732, n19415, n19395, n19193, n19196, 
        n19411, n19079, n19161, n39696, n19607, n19626, n181_adj_31, 
        n18636, n19608, n19416, n19396, n145, n19407, n19082, 
        n19402, n19625, n19793, n19609, n19413, n19397, n19420, 
        n19424, n19412, n19083, n142, n19158, n40545, n37334, 
        n38589, clk_c_enable_832, n19624, n19610, n167_adj_32, n18559, 
        n19623, n19611, n19418, n19400, n19474, n19074, n18918, 
        n19479, n19466, n40544, n19622, n19612, n166_adj_33, n19621, 
        n18558, n18982, n19399, n18992, n19073, n18917, n19090, 
        n19465, n19480, n36872, n19613, n19620, n19614, n19619, 
        n19738, n18985, n19467, n18993, n19006, n19615, n19088, 
        n19423, n18914, n38587, n19618, n19616, n167_adj_34, n190_adj_35, 
        n19742, n19417, n19000, n19472, n19007, n18557, n19087, 
        n19421, n18913, n40543, n19617, n19553, n171_adj_36, n19520, 
        n19741, n19414, n19001, n18994, n19008, n18556, n19086, 
        n18977, n40542, n40541, n40540, n39687, n19554, n19519, 
        n19555, n19518, n19740, n19739, n139, n19404, n19471, 
        n19041, n19525, n19085, n39685, n40539, n19556, n19517, 
        n169_adj_37, n18555, n19557, n136, n19159, n19784, n18916, 
        n19775, n19787, n19093, n40538, n40537, n19516, n19558, 
        n19772, n19559, n18554, n19398, n19473, n18986, n19084, 
        n133, n18978, n40536, n40535, n19560, n175_adj_38, n19561, 
        n130, n19776, n19766, n19098, n19042, n19524, n40534, 
        n40532, n40531, n19562, n127, n19563, n19528, n19564, 
        n19419, n19401, n18989, n19756, n18915, n19780, n19765, 
        n19565, n38582, n18940, n124, n19096, n19043, n19523, 
        n19566, n19091, n40530, n40529, n40528, n40527, n19567, 
        n178_adj_39, n19568, n19781, n121, n19095, n19044, n19773, 
        n18553, n19569, n19078, n40526, n39678, n19570, n32870, 
        n19571, n177_adj_40, n19094, n19081, n18925, n18552, n176_adj_41, 
        n118, n25246, n25250, n19572, n32869, n25252, n19573, 
        n115, n25254, n19574, n25256, n19575, n32868, n25258, 
        n19576, n112, n25260, n19577, n25262, n19578, n40525, 
        n32867, n25264, n19579, n32456, n40524, n32452, n32451, 
        n32450, n32449, n32444, n32443, n32442, n32438, n32437, 
        n32436, n109, n32435, n19580, n32434, n32433, n32432, 
        n19581, n32431, n19702, n32430, n32866, n19582, n106, 
        n19583, n192_adj_42, n19737, n19779, n19786, n19422, n19077, 
        n32865, n18922, n19584, n19778, n32864, n19768, n19297, 
        n19405, n19298, n19299, n19300, n19301, n19302, n19303, 
        n19304, n19305, n19306, n19307, n19308, n19309, n19310, 
        n19311, n19312, n39671, n19313, n19314, n19315, n19316, 
        n19317, n19318, n19769, n19319, n19320, n18551, n18984, 
        n19789, n19321, n40523, n19478, n18932, n19764, n19322, 
        n40522, n19323, n19324, n19325, n19326, n19327, n18921, 
        n19790, n19328, n18635, n19100, n18919, n19329, n18926, 
        n37374, n18550, n19449, n18634, n19330, n18633, n32429, 
        n32863, n19331, n39667, n18632, n19332, n18631, n38576, 
        n19333, n32428, n18630, n19334, n18629, n19783, n19335, 
        n18628, n19336, n18627, n19337, n18626, n70, n19521, n19338, 
        n18979, n18625, n170_adj_43, n19339, n193_adj_44, n32427, 
        n19099, n103, n18923, n18549, n18624, n19340, n18623, 
        n19341, n18622, n18548, n18981, n18980, n172_adj_45, n19712, 
        n19075, n19342, n13381, n40521, n40520, n40519, n40517, 
        n40516, n19477, n18621, n19743, clk_c_enable_780, n40515, 
        n19343, n18620, n168_adj_46, n191_adj_47, n18941, n19527, 
        n18988, n18987, n19782, n19759, n32862, n19483, n18995, 
        n19522, n40514, n39660, n38571, n19344, n18983, n19470, 
        n19771, n19758, n100, n19482, n19469, n19744, clk_c_enable_829, 
        n194_adj_48, n18547, n18927, n18997, n19770, n19757, n19481, 
        n18998, n19774, n30887, n40513, n40512, n18619, n19751, 
        n32861, n18546, n18931, n106_adj_49, n20127, n18928, n39656, 
        n20133, n19447, n40511, n20147, n19002, n37336, n19051, 
        n40510, n40509, n37513, n19463, n40508, n19052, n19791, 
        n18545, n40507, n112_adj_50, n187_adj_51, n19762, n18544, 
        n40506, clk_c_enable_812, n18618, n115_adj_52, n19345, n18617, 
        n19346, n19460, n18616, n20128, n19347, n18615, n19348, 
        n18614, n19349, n136_adj_53, n18613, n19350, n18612, n19351, 
        n18611, n19005, n19352, n18610, n20130, n19353, n18609, 
        n19354, n18608, n19355, n18607, n19356, n18543, n18606, 
        n19357, n20144, n18605, n19358, n18604, n19031, n25306, 
        n32426, n32425, n32391, n32385, n32384, n32383, n32382, 
        n32381, n32380, n32379, n32378, n32377, n32376, n40505, 
        n40504, n40502, n40501, n38562, n39646, n40500, n40499, 
        n40498, n40497, n40496, n40495, n40494, n40493, n40492, 
        n39641, n40491, n40490, n39636, n25266, n25268, n25270, 
        n25272, n25274, n25276, n25278, n16519, n19359, n18603, 
        n19360, n194_adj_54, n193_adj_55, n38555, n192_adj_56, n191_adj_57, 
        n190_adj_58, n32375, n189_adj_59, n188_adj_60, n187_adj_61, 
        n186_adj_62, n185_adj_63, n18542, n184_adj_64, n183_adj_65, 
        n182_adj_66, n32374, n181_adj_67, n20146, n180_adj_68, n179_adj_69, 
        n178_adj_70, n177_adj_71, n176_adj_72, n175_adj_73, n32373, 
        n174_adj_74, n173_adj_75, n172_adj_76, n171_adj_77, n19030, 
        n170_adj_78, n169_adj_79, n168_adj_80, n32372, n167_adj_81, 
        n166_adj_82, n165_adj_83, n164_adj_84, n19802, n19453, n36532, 
        n32371, n163_adj_85, n19451, n19443, n18541, n32370, n18540, 
        n19441, n39634, n18539, n19440, n32369, n18538, n19438, 
        n40489, n18537, n19437, n40487, n32368, n18536, n19752, 
        n19428, n40486, n19427, n40485, n32367, n18535, n19425, 
        n18534, n32366, n18533, n18532, n18531, n18530, n32365, 
        n18529, n18929, n18528, n18527, n18526, n32860, n18525, 
        n18524, n19456, n32364, n18523, n18522, n19455, n19454, 
        n18602, n19533, n19729, n32363, n19452, n20131, n19700, 
        n19727, n19725, n18601, n19722, n19546, n32362, n19442, 
        n18521, n19704, n19717, n19551, n19050, n18600, n19650, 
        n19654, n32361, n19439, n32859, n19705, n19656, n19659, 
        n18599, n19662, n19665, n32360, n19436, n19708, n19668, 
        n19670, n20135, n18598, n19672, n19674, n40484, n40483, 
        n32359, n32358, n32357, n40482, n25244, n39629, n40481, 
        n40480, n40479, n38551, n40478, n40477, n40476, n18520, 
        n15805, n18519, n18518, n18517, n18516, n18515, n18514, 
        n18513, n18512, n18511, n18510, n18509, n18508, n19809, 
        n32858, n19810, n97, n19435, n19433, n189_adj_86, n19811, 
        n19812, n19430, n32857, n19813, n19448, n94, n19814, n19429, 
        n19815, n32856, n40475, n40474, n38546, n40472, n40471, 
        n39618, n42492, n38536, n40470, n40469, n40468, n42491, 
        n39614, n37411, n42440, n40467, n37672, n40466, n37670, 
        n39609, n37298, n38533, n38531, n42439, n40465, n40464, 
        n40463, n40462, n39602, n42490, n40461, n40460, n40459, 
        n40457, n37417, n39593, n42438, n39591, n42437, n40456, 
        n40455, n40454, n40453, n40452, n40451, n42489, n40450, 
        n40449, n36832, n38517, n37286, n39576, n38515, n40448, 
        n37284, n40447, n40446, n40445, n39573, n40444, n37282, 
        n40442, n40441, n40440, n40439, n40438, n40437, n32855, 
        n91, n32854, n88, n32853, n85, n18794, n18795, n18796, 
        n18797, n18798, n18799, n18800, n18801, n18802, n18803, 
        n18804, n18805, n18806, n18807, n18808, n18809, n18810, 
        n18811, n18812, n18813, n18814, n18815, n18816, n32356, 
        n32355, n32354, n32390, n33, n32, n31, n30, n29, n28, 
        n27, n26, n25, n24, n23, n22, n21, n32852, n19816, 
        n82, n19817, n19753, n19818, n32851, n19819, n18753, n18754, 
        n18755, n18756, n18757, n18758, n18759, n18760, n18761, 
        n79, n32850, n76, n32849, n73, n32848, n70_adj_87, n39566, 
        n32847, n32846, n32845, n32844, n32843, n20, n32842, n19, 
        n18, n17, n16, n15, n14, n13, n18597, n19707, n12, 
        n11, n19820, n10, n40436, n9, n18817, n18818, n18819, 
        n18820, n18821, n18822, n18823, n18824, n18825, n18826, 
        n18827, n18828, n18829, n18830, n18831, n18832, n18833, 
        n18834, n18835, n18836, n18837, n18838, n18839, n18840, 
        n18841, n18842, n18843, n18844, n18845, n18846, n18847, 
        n18848, n40435, n19821, n32841, n19822, n19823, n32840, 
        n19824, n37276, n19825, n32839, n19826, n19827, n32838, 
        n18912, n18849, n18850, n18851, n18852, n18853, n18854, 
        n18855, n18856, n18857, n18858, n18859, n18860, n18861, 
        n18862, n18863, n18864, n18865, n18866, n18867, n18868, 
        n18869, n18870, n18871, n18872, n18873, n18874, n18875, 
        n18876, n18877, n18878, n18879, n18880, n19828, n32837, 
        n19829, n32836, n19830, n19003, n8, n7, n6, n5, n4, 
        n3, n32392, n19426, n19054, n19709, n19676, n19678, n18596, 
        n18721, n18722, n18723, n18724, n18725, n18726, n18727, 
        n18728, n18729, n18730, n18731, n18732, n18733, n18734, 
        n18735, n18736, n18737, n18738, n18739, n18740, n18741, 
        n18742, n18743, n18744, n18745, n18746, n18747, n18748, 
        n18749, n18750, n18751, n18752, n38502, n19831, n32835, 
        n18507, n180_adj_88, n19076, n19080, n18924, n19777, n179_adj_89, 
        n19406, n38499, n5193, n5194, n5195, n5196, n5197, n5198, 
        n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, 
        n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, 
        n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
        n5223, n5224, n19832, n25280, n25282, n25284, n25286, 
        n25288, n25290, n25292, n25294, n25296, n25298, n25300, 
        n25302, n25304, n19431, n19701, n19231, n133_adj_90, n19175, 
        n20142, n19803, n19434, n19799, n19230, n19047, n32834, 
        n20143, n19445, n32833, n19363, n19833, n18506, n32832, 
        n30987, n5325, n5326, n5327, n5328, n5329, n5330, n5331, 
        n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
        n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, 
        n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
        n5356, n32831, n32830, n40434, n5460, n5461, n5462, n5463, 
        n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
        n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
        n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, 
        n5488, n5489, n5490, n5491, n5494, n5495, n5496, n5497, 
        n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, 
        n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
        n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
        n5522, n5523, n5524, n5525, n85_adj_91, n40433, n19834, 
        n19462, n19055, n103_adj_92, n19792, n18505, n32829, n188_adj_93, 
        n19761, n18504, n32828, n19461, n20132, n32827, n37657, 
        n18503, n19004, n20134, n139_adj_94, n19169, n20148, n19028, 
        n19754, n18502, n20150, n19027, n37274, n19048, n73_adj_95, 
        n18501, n18935, n20108, n19032, n20136, n19053, n37272, 
        n20139, n18595, n142_adj_96, n32826, n164_adj_97, n19476, 
        n32825, n19046, n20107, n32824, n19706, n19232, n20137, 
        n19049, n79_adj_98, n20105, n19835, n19034, n130_adj_99, 
        n20145, n18990, n19432, n18594, n19228, n38491, n19172, 
        n20138, n32823, n19836, n19837, n19446, n19800, n19227, 
        n19029, n118_adj_100, n20140, n18911, n32822, n76_adj_101, 
        n19703, n19173, n127_adj_102, n19844, n19035, n20106, n145_adj_103, 
        n19801, n32821, n19174, n18933, n82_adj_104, n20112, n165_adj_105, 
        n19475, n19749, n40432, n19045, n20111, n19838, n19229, 
        n20141, n36818, n40431, n19804, n39557, n18934, n32820, 
        n20109, n19843, n19033, n32819, n20149, n18991, n19750, 
        n109_adj_106, n19839, n18593, n19170, n40430, n32818, n163_adj_107, 
        n19036, n20110, n32817, n19755, n32816, n18500, n19682, 
        n19842, n19710, n18499, n19685, n18498, n18497, n19688, 
        n19840, n40429, n19711, n19689, n19690, n186_adj_108, n19691, 
        n19692, n19841, n185_adj_109, n19693, n19694, n19171, n184_adj_110, 
        n18496, n19695, n18881, n19392, n183_adj_111, n18495, n19696, 
        n182_adj_112, n18494, n19697, n18882, n18493, n18492, n19698, 
        n19450, n18491, n18490, n19699, n19391, n18883, n19390, 
        n18884, n19389, n18930, n18885, n19388, n18886, n19387, 
        n18887, n19386, n18888, n32815, n19385, n18889, n19384, 
        n18890, n19383, n18891, n19382, n18892, n19381, n18893, 
        n19380, n18894, n19379, n18895, n19378, n18896, n19377, 
        n18897, n19376, n18898, n19375, n20129, n18899, n19374, 
        n18900, n19373, n18901, n19372, n18902, n19371, n19361, 
        n18903, n19641, n19592, n19642, n19591, n19643, n19590, 
        n19644, n19589, n19645, n19588, n19646, n19587, n19647, 
        n19586, n19648, n19585, n18489, n18488, n18487, n18486, 
        n18485, n18484, n18483, n18482, n18481, n18480, n18479, 
        n18478, n18477, n18476, n19370, n19444, n18904, n19369, 
        n18905, n148_adj_113, n19368, n18906, n19367, n32814, done_N_1929, 
        done_N_1931, done_N_1932, done_N_1934, n32813, n40427, done_N_1928, 
        n32812, n40426, n38479, n38474, n40425, n40424, n39546, 
        n39544, n37646, n38472;
    wire [511:0]U_0__31__N_967;
    
    wire n40423, n40422, n40421, n40420, n40419, n40418, n38467, 
        n39535, n38456, n40417, n40416, n40415, n40414, n40412, 
        n40411, n39531, n38452, n40410, n40409, n40408, n39525, 
        n38447, n37258, n40407, n40406, n40405, n40404, n39520, 
        n37256, n36802, n40403, n40402, n39514, n38440, n39511, 
        n40401;
    wire [31:0]i_31__N_1607;
    
    wire n37252, n40400, n40399, n38431, n40397, n40396, n40395, 
        n40394, n37250, n37462, n39504, n38429, n40393, n40392, 
        n39500, n40391, n40390, n40389, n40388, n40387, n40386, 
        n40385, n40384, n40382, n19252, n18475, n18474, n39493, 
        n40381, n37244, n39487, n40380, n40379, n40378, n37242, 
        n40377, n40376, n40375, n40374, n39482, n39480, n40373, 
        n40372, n37240, n36784, n40371, n40370, n40369, n40367, 
        n40366, n40365, n37238, n40364, n40363, n38414, n39466, 
        n38411, n38409, n40362, n40361, n40360, n40359, n40358, 
        n40357, n40356, n40355, n40354, n40352, n39458, n39456, 
        n40351, n40350, n40349, n40348, n40347, n40346, n39451, 
        n40345, n40344, n38397, n40343, n40342, n40341, n40340, 
        n40339, n39445, n40337, n40336, n40335, n40334, n40333, 
        n37480, n40332, n40331, n40330, n40329, n39440, n40328, 
        n38395, n40327, n40326, n40325, n40324, n40322, n40321, 
        n37218, n40320, n9902, n9901, n40319, n32811, n32810, 
        n20406, n20405, n20404, n20403, n20402, n20401, n20400, 
        n20375, n19275, n18473, n19276, n18472, n32809, n18967, 
        n32808, n32807, n32806, n32805, n32804, n32803, n32802, 
        n32801, n20414, n20413, n20412, n20411, n20410, n20409, 
        n20408, n20431, n18471, n19274, n18470, n18469, n18968, 
        n32800, n32799, n32798, n40318, n32797, n32796, n32795, 
        n32794, n40317, n20422, n20421, n20420, n20419, n20418, 
        n20417, n20416, n20423, n19268, n18468, n19269, n18467, 
        n18466, n18969, n32793, n32792, n32791, n32790, n32789, 
        n32788, n40316, n32787, n32786, n20430, n20429, n20428, 
        n20427, n20426, n20425, n20424, n20415, n19261, n19262, 
        n19263, n18465, n19122, n18970, n32785, n32784, n32783, 
        n32782, n32781, n40315, n20438, n20437, n20436, n20435, 
        n20434, n18907, n10098, n18971, n32780, n32779, n32778, 
        n32777, n20432, n20407, n19250, n19251, n32776, n19366, 
        n18908, n19365, n18909, n32775, n39431, n36760, n40314, 
        n37431, n40313, n40312, n37212, n40311, n40310, n40309, 
        n40307, n40306, n40305, n40304, n39424, n40303, n37210, 
        n40302, n36756, n39420, n38384, n38382, n37206, n25248, 
        n36752, n38373, n40301, n40300, n39415, n40299, n40298, 
        n40297, n32773, n20446, n20445, n20444, n20443, n20442, 
        n20441, n20440, n20463, n19239, n19240, n19241, n18464, 
        n19117, n18972, n32772, n32771, n32770, n40296, n32769, 
        n32768, n20454, n20453, n20452, n20451, n20450, n20449, 
        n20448, n20455, n19877, n32767, n18463, n18462, n18461, 
        n32766, n32765, n32764, n32763, n32762, n20462, n20461, 
        n20460, n20459, n20458, n20457, n20456, n20447, n19888, 
        n19887, n19886, n18460, n19112, n18459, n40295, n32761, 
        n60, n32760, n32759, n32756, n20470, n20469, n20468, n20467, 
        n20466, n20465, n20464, n20439, n19899, n19898, n19897, 
        n18458, n18457, n18456, n32755, n32754, n32753, n40294, 
        n32752, n32751, n20478, n20477, n20476, n20475, n20474, 
        n20473, n20472, n20505, n19910, n19909, n19908, n18455, 
        n19107, n18454, n32750, n32749, n32748, n32747, n32746, 
        n32745, n20486, n20485, n20484, n20483, n20482, n20481, 
        n20480, n20553, n19921, n19920, n19919, n194_adj_114, n18453, 
        n194_adj_115, n32744, n32743, n32742, n32738, n32737, n32736, 
        n32735, n32734, n32733, n32732, n32731, n32730, n32729, 
        n20494, n20506, n20508, n20487, n20511, n20495, n20509, 
        n20479, n192_adj_116, n191_adj_117, n190_adj_118, n189_adj_119, 
        n189_adj_120, n188_adj_121, n32728, n32727, n32726, n32725, 
        n32724, n32719, n32718, n32717, n32716, n32715, n32714, 
        n32713, n20496, n20544, n20512, n20488, n20522, n20497, 
        n20523, n20471, n187_adj_122, n186_adj_123, n185_adj_124, 
        n184_adj_125, n183_adj_126, n182_adj_127, n32712, n32711, 
        n32710, n32709, n32708, n32707, n32706, n36746, n32702, 
        n32701, n32700, n32699, n32698, n32697, n20498, n20548, 
        n20514, n20489, n20526, n20499, n20527, n20550, n182_adj_128, 
        n181_adj_129, n180_adj_130, n179_adj_131, n177_adj_132, n176_adj_133, 
        n38364, n32696, n32695, n32694, n32693, n32692, n32691, 
        n32690, n32689, n32684, n32683, n32682, n32681, n20500, 
        n20551, n20516, n20490, n20535, n20501, n20541, n32680, 
        n177_adj_134, n176_adj_135, n175_adj_136, n174_adj_137, n171_adj_138, 
        n170_adj_139, n32679, n32678, n32677, n32676, n32675, n32674, 
        n32673, n32672, n32668, n32667, n32666, n20502, n20554, 
        n20518, n20491, n20536, n20503, n32665, n20556, n172_adj_140, 
        n171_adj_141, n170_adj_142, n169_adj_143, n166_adj_144, n165_adj_145, 
        n32664, n32663, n32662, n32661, n32660, n32659, n32658, 
        n32657, n32656, n32651, n32650, n32649, n20510, n20557, 
        n20521, n20492, n20537, n20507, n20547, n167_adj_146, n166_adj_147, 
        n165_adj_148, n164_adj_149, n18452, n18451, n32648, n32647, 
        n32646, n32645, n32644, n32643, n32642, n32641, n161, 
        n32640, n158, n20520, n20560, n20525, n20493, n20538, 
        n20513, n20563, n19967, n18450, n18449, n18448, n18447, 
        n18446, n155, n32636, n152, n32635, n149, n32634, n146, 
        n32633, n143, n39405, n20524, n20564, n20528, n20504, 
        n20539, n20515, n32632, n19972, n18445, n18444, n18443, 
        n18442, n18441, n32631, n140, n32630, n137, n32629, n134, 
        n32628, n131, n40292, n32627, n128, n20542, n32626, n20529, 
        n20546, n20543, n20517, n32625, n18440, n18439, n18438, 
        n18437, n18436, n18435, n125, n122, n32620, n119, n32619, 
        n116, n38362, n32618, n113, n40291, n32617, n20530, n20561, 
        n20549, n20519, n20559, n18434, n18433, n32616, n32615, 
        n32614, n110, n32613, n107, n32612, n104, n32611, n101, 
        n32610, n98, n38360, n20531, n20565, n20552, n20545, n32606, 
        n32605, n32604, n31084, n32603, n95, n32602, n92, n32601, 
        n89, n32600, n86, n32599, n83, n32598, n32597, n20532, 
        n32596, n20555, n20562, n36744, n38357, n32591, n80, n32590, 
        n77, n32589, n74, n32588, n71, n32587, n68, n32586, 
        n20533, n20558, n20566, n32585, n32584, n32583, n32582, 
        n32578, n32577, n32576, n32575, n32574, n32573, n32572, 
        n32571, n32570, n32569, n20534, n32564, n32563, n32562, 
        n19072, n19010, n19071, n19011, n32561, n32560, n32559, 
        n32558, n32557, n32556, n32552, n32551, n20540, n40290, 
        n19012, n19069, n19013, n19068, n32550, n32549, n32548, 
        n32547, n32546, n32545, n32544, n32539, n32538, n32537, 
        n19067, n19015, n20114, n19066, n32536, n32535, n32534, 
        n32533, n32532, n32528, n32527, n32526, n32525, n121_adj_150, 
        n19065, n19017, n20116, n19064, n32524, n32523, n32522, 
        n32521, n40289, n32516, n32515, n32514, n32513, n32512, 
        n32511, n32510, n88_adj_151, n94_adj_152, n19063, n19019, 
        n20118, n20093, n32506, n32505, n32504, n32503, n32502, 
        n32501, n32500, n32495, n32494, n32493, n32492, n32491, 
        n32490, n32486, n40288, n19020, n19061, n20120, n20096, 
        n19745, n19808, n32485, n32484, n32483, n32482, n32481, 
        n32476, n32475, n32474, n40287, n32473, n97_adj_153, n32472, 
        n40286, n124_adj_154, n40285, n19060, n19022, n20122, n20099, 
        n19746, n19807, n39400, n32468, n163_adj_155, n32467, n160_adj_156, 
        n32466, n157_adj_157, n32465, n154_adj_158, n32464, n151_adj_159, 
        n91_adj_160, n100_adj_161, n19023, n19058, n20124, n19024, 
        n19747, n19806, n36740, n32459, n32458, n32457, n19025, 
        n19056, n20126, n20104, n19748, n19805, n40284, n40283, 
        n38346, n19362, n19364, n18910, n38337, n38335, n40282, 
        n40281, n40280, n40279, n40277, n40276, n40275, n40274, 
        n39386, n40273, n40272, n39384, n38330, n40271, n36734, 
        n40270, n38321, n40269, n40268, n40267, n40266, n38314, 
        n40265, n39371, n40264, n40262, n40261, n40260, n39368, 
        n37186, n23957, n40259, n40258, n40257, n40256, n38301, 
        n40255, n40254, n40253, n39360, n38297, n38294, n40252, 
        n40251, n40250, n40249, n39351, n39349, n32393, n32394, 
        n32395, n32396, n32397, n32398, n32399, n32400, n32401, 
        n32402, n32403, n32404, n32405, n32407, n40247, n32408, 
        n32409, n32410, n32411, n32412, n32413, n40246, n32414, 
        n32415, n32416, n32417, n32418, n32419, n32420, n60_adj_162, 
        n32421, n32422, n32423, n40245, n32424, n40244, n39340, 
        n38282, n40243, n40242, n40241, n40240, n40239, n39331, 
        n40238, n38274, clk_c_enable_541, n39328, n40237, n40236, 
        n37180, n39326, n39324, n40235, n40234, n40232, n40231, 
        n37178, n63, n38269, n40230, n40229, n37176, n40228, n40227, 
        n40226, n36720, n39311, n40225, n39308, n2, n3_adj_163, 
        n4_adj_164, n5_adj_165, n6_adj_166, n7_adj_167, n8_adj_168, 
        n9_adj_169, n10_adj_170, n11_adj_171, n12_adj_172, n13_adj_173, 
        n14_adj_174, n15_adj_175, n16_adj_176, n17_adj_177, n18_adj_178, 
        n19_adj_179, n20_adj_180, n21_adj_181, n22_adj_182, n23_adj_183, 
        n24_adj_184, n25_adj_185, n26_adj_186, n27_adj_187, n28_adj_188, 
        n29_adj_189, n30_adj_190, n31_adj_191, n32_adj_192, n33_adj_193, 
        n39306, n40224, n27528, n27533, n37172, n40223, n68_adj_194, 
        n69, n70_adj_195, n71_adj_196, n72, n73_adj_197, n74_adj_198, 
        n75, n76_adj_199, n77_adj_200, n78, n79_adj_201, n80_adj_202, 
        n81, n82_adj_203, n83_adj_204, n84, n85_adj_205, n86_adj_206, 
        n87, n88_adj_207, n89_adj_208, n90, n91_adj_209, n92_adj_210, 
        n93, n94_adj_211, n95_adj_212, n96, n97_adj_213, n98_adj_214, 
        n99, n102, n103_adj_215, n104_adj_216, n105, n106_adj_217, 
        n107_adj_218, n108, n109_adj_219, n110_adj_220, n111, n112_adj_221, 
        n113_adj_222, n114, n115_adj_223, n116_adj_224, n117, n118_adj_225, 
        n119_adj_226, n120, n121_adj_227, n122_adj_228, n123, n124_adj_229, 
        n125_adj_230, n126, n127_adj_231, n128_adj_232, n129, n130_adj_233, 
        n131_adj_234, n132, n40222, n40221, n40220, n40219, n40217, 
        n40216, n39296, n38257, n40215, n40214, n40213, n40212, 
        n40211, n40210, n35961, n39291, n40209, n39289, n40208, 
        n38255, n40207, n40206, n40205, n40204, n40202, n39284, 
        n38250, n38244, n40201, n40200, n40199, n40198, n39273, 
        n40197, n678, n682, n683, n684, n685, n40196, n36704, 
        n38239, n39269, n708, n30965, n30968, n40195, n36702, 
        n40194, n39264, n36700, n40193, n40192, n38230, n864, 
        n865, n872, n873, n874, n875, n876, n877, n878, n879, 
        n880, n881, n882, n883, n884, n885, n886, n887, n888, 
        n889, n890, n891, n892, n893, n40191, n40190, n36698, 
        n40189, n40187, n37154, n40186, n40185, n39257, n36696, 
        n38223, n1047, n1048, n1049, n40184, n36694, n40183, n1078, 
        n38219, n40182, n30872, n30944, n40181, n40180, n40179, 
        n39248, n40178, n39246, n40177, n40176, n1227, n1228, 
        n1229, n1230, n36692, n37148, n40175, n38214, n40174, 
        n40172, n40171, n40170, n40169, n36690, n40168, n1403, 
        n1404, n1405, n1406, n1407, n1408, n36688, n40167, n40166, 
        n37146, n36686, n40165, n39231, n1462, n30929, n30926, 
        n40164, n39228, n40163, n40162, n40161, n36684, n37144, 
        n40160, n40159, n40157, n39226, n1577, n1578, n1579, n1580, 
        n1581, n1582, n1583, n37370, n40156, clk_c_enable_677, n38204, 
        n40155, n1635, n30920, n30938, n40154, n40153, n40152, 
        n36682, n38199, n40151, n1748, n1749, n1750, n1751, n1752, 
        n1753, n1754, n1755, n40150, n39214, n38194, n39212, n36680, 
        n1805, n30914, n30932, n40149, n36678, n40148, n40147, 
        n40146, n36676, n1916, n1917, n1918, n1919, n1920, n1921, 
        n1922, n1923, n1924, n40145, n30917, n30923, n40144, n38185, 
        n39201, n38183, n39199, n40142, n40141, n40140, n36674, 
        n40139, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
        n2088, n2089, n2090, n36672, n40138, n40137, n30908, n2137, 
        n56, n2141, n2142, n39190, n40136, n40135, n40134, n2243, 
        n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, 
        n2252, n2253, n36670, n39186, n40133, n39184, n40132, 
        n30905, n2298, n40131, n40130, n38170, n36668, n40129, 
        n40127, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
        n2409, n2410, n2411, n2412, n2413, n37495, n36666, n40126, 
        n40125, n2455, n2456, n40124, n37122, n30890, n30950, 
        n40123, n40122, n39171, n40121, n36664, n40120, n39168, 
        n40119, n38167, n40118, n37120, n2558, n2559, n2560, n2561, 
        n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
        n2570, n40117, n40116, n40115, n40114, n30902, n30911, 
        n39166, n39164, n36662, n40110, n2711, n2712, n2713, n2714, 
        n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
        n2723, n2724, n40108, n38159, n36660, n2762, n55, n40104, 
        n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
        n2869, n2870, n2871, n2872, n2873, n2874, n2875, n36658, 
        n39150, n38150, n38148, n2911, n30896, n36656, n3008, 
        n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
        n3017, n3018, n3019, n3020, n3021, n3022, n3023, n40102, 
        n39146, n3057, n30893, n3060, n36654, n40100, n39143, 
        n36652, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
        n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
        n3167, n3168, n38137, n40096, n38136, n40094, n36650, 
        n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, 
        n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
        n3309, n3310, n40092, n39133, n39131, n39129, n3340, n38134, 
        n40090, n36648, n3431, n3432, n3433, n3434, n3435, n3436, 
        n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, 
        n3445, n3446, n3447, n3448, n3449, n40086, n35925, n3477, 
        n3479, n36646, n39126, n38127, n3566, n3567, n3568, n3569, 
        n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
        n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, 
        n38125, n36644, n3611, n40082, n38114, n3698, n3699, n3700, 
        n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, 
        n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, 
        n3717, n3718, n38111, n35922, n4_adj_235, n40080, n39115, 
        n37469, n42488, n40078, n3827, n3828, n3829, n3830, n3831, 
        n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, 
        n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
        n3848, n36642, n3870, n3871, n38101, n38099, n38096, clk_c_enable_708, 
        n40074, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
        n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
        n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, 
        n39106, n39104, n3995, n38087, n4076, n4077, n4078, n4079, 
        n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, 
        n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, 
        n4096, n4097, n4098, n4099, n4117, n39099, n4196, n4197, 
        n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, 
        n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
        n4214, n4215, n4216, n4217, n4218, n4219, n4220, n36636, 
        n38080, n37440, n4236, n4313, n4314, n4315, n4316, n4317, 
        n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, 
        n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
        n4334, n4335, n4336, n4337, n4338, n4352, n39090, n4427, 
        n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, 
        n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
        n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, 
        n4452, n4453, n35955, n4465, n39083, n37092, n40061, n4538, 
        n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
        n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, 
        n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
        n4563, n4564, n4565, n38067, n40059, n40057, n4646, n4647, 
        n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, 
        n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
        n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, 
        n4672, n4673, n4674, n35919, n4682, n4683, n42487, n22242, 
        n22243, n22244, n22245, n22246, n22247, n22248, n22249, 
        n22250, n22251, n22252, n22253, n22254, n22255, n22256, 
        n22257, n22258, n22259, n22260, n22261, n22262, n22263, 
        n22264, n22265, n22266, n22267, n22268, n22269, n22270, 
        n22271, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
        n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, 
        n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
        n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4783, 
        n40053, n39066, n22241, n39063, n4883, n4885, n22306, 
        n22305, n22304, n22303, n22302, n22301, n22300, n22299, 
        n22298, n22297, n22296, n22295, n22294, n22293, n22292, 
        n22291, n22290, n22289, n22288, n22287, n22286, n22285, 
        n22284, n22283, n22282, n22281, n22280, n22279, n22278, 
        n22277, n22276, n22275, n38058, n37364, n42486, n40043, 
        n42485, n42484, n37082, n38054, n39051, n38050, n36624, 
        n42483, n58, n60_adj_236, n62, n64, n40035, n39043, n42482, 
        n38041, n42481, n56_adj_237, n57, n58_adj_238, n60_adj_239, 
        n62_adj_240, n64_adj_241, n40033, n39038, n38036, n37508, 
        n38034, n54, n56_adj_242, n58_adj_243, n60_adj_244, n61, 
        n62_adj_245, n64_adj_246, n37380, n39028, n40027, n37482, 
        n52, n54_adj_247, n56_adj_248, n58_adj_249, n59, n60_adj_250, 
        n62_adj_251, n64_adj_252, n42480, n37379, n40021, n50, n52_adj_253, 
        n54_adj_254, n56_adj_255, n57_adj_256, n58_adj_257, n60_adj_258, 
        n62_adj_259, n64_adj_260, n37378, n38020, n39017, n37377, 
        n39015, n39011, n40017, n48, n49, n50_adj_261, n52_adj_262, 
        n54_adj_263, n55_adj_264, n56_adj_265, n58_adj_266, n60_adj_267, 
        n62_adj_268, n64_adj_269, n39004, n46, n48_adj_270, n50_adj_271, 
        n51, n52_adj_272, n53, n54_adj_273, n56_adj_274, n58_adj_275, 
        n60_adj_276, n62_adj_277, n64_adj_278, n40011, n38012, n36606, 
        n40007, n38999, n44, n45, n46_adj_279, n48_adj_280, n50_adj_281, 
        n51_adj_282, n52_adj_283, n54_adj_284, n56_adj_285, n58_adj_286, 
        n60_adj_287, n62_adj_288, n64_adj_289, n38990, n42, n44_adj_290, 
        n46_adj_291, n47, n48_adj_292, n49_adj_293, n50_adj_294, n52_adj_295, 
        n54_adj_296, n56_adj_297, n58_adj_298, n60_adj_299, n62_adj_300, 
        n64_adj_301, n39999, n38007, n40, n42_adj_302, n44_adj_303, 
        n45_adj_304, n46_adj_305, n47_adj_306, n48_adj_307, n50_adj_308, 
        n52_adj_309, n54_adj_310, n56_adj_311, n58_adj_312, n60_adj_313, 
        n62_adj_314, n64_adj_315, n39995, n38982, n38, n39, n40_adj_316, 
        n42_adj_317, n43, n44_adj_318, n46_adj_319, n48_adj_320, n50_adj_321, 
        n52_adj_322, n54_adj_323, n56_adj_324, n58_adj_325, n60_adj_326, 
        n62_adj_327, n64_adj_328, n38980, n39991, n38003, n36, n38_adj_329, 
        n40_adj_330, n41, n42_adj_331, n43_adj_332, n44_adj_333, n46_adj_334, 
        n48_adj_335, n50_adj_336, n52_adj_337, n54_adj_338, n56_adj_339, 
        n58_adj_340, n60_adj_341, n62_adj_342, n64_adj_343, n39989, 
        n37054, n39987, n39985, n34, n36_adj_344, n38_adj_345, n39_adj_346, 
        n40_adj_347, n41_adj_348, n42_adj_349, n44_adj_350, n46_adj_351, 
        n48_adj_352, n50_adj_353, n52_adj_354, n54_adj_355, n56_adj_356, 
        n58_adj_357, n60_adj_358, n62_adj_359, n64_adj_360, n38975, 
        n32_adj_361, n33_adj_362, n34_adj_363, n36_adj_364, n37, n38_adj_365, 
        n40_adj_366, n42_adj_367, n44_adj_368, n46_adj_369, n48_adj_370, 
        n50_adj_371, n52_adj_372, n54_adj_373, n56_adj_374, n58_adj_375, 
        n60_adj_376, n62_adj_377, n64_adj_378, n38969, n37998, n42479, 
        n30_adj_379, n31_adj_380, n32_adj_381, n34_adj_382, n35, n36_adj_383, 
        n37_adj_384, n38_adj_385, n40_adj_386, n42_adj_387, n44_adj_388, 
        n46_adj_389, n48_adj_390, n50_adj_391, n52_adj_392, n53_adj_393, 
        n54_adj_394, n56_adj_395, n58_adj_396, n60_adj_397, n62_adj_398, 
        n64_adj_399, n37988, n37985, n37637, n37635, n28_adj_400, 
        n30_adj_401, n32_adj_402, n33_adj_403, n34_adj_404, n35_adj_405, 
        n36_adj_406, n38_adj_407, n40_adj_408, n42_adj_409, n44_adj_410, 
        n46_adj_411, n48_adj_412, n50_adj_413, n51_adj_414, n52_adj_415, 
        n54_adj_416, n56_adj_417, n58_adj_418, n60_adj_419, n62_adj_420, 
        n64_adj_421, n42478, n37632, n26_adj_422, n28_adj_423, n30_adj_424, 
        n31_adj_425, n32_adj_426, n34_adj_427, n36_adj_428, n37_adj_429, 
        n38_adj_430, n40_adj_431, n42_adj_432, n44_adj_433, n46_adj_434, 
        n48_adj_435, n49_adj_436, n50_adj_437, n52_adj_438, n54_adj_439, 
        n56_adj_440, n58_adj_441, n60_adj_442, n62_adj_443, n64_adj_444, 
        n24_adj_445, n25_adj_446, n26_adj_447, n28_adj_448, n29_adj_449, 
        n30_adj_450, n32_adj_451, n34_adj_452, n35_adj_453, n36_adj_454, 
        n38_adj_455, n40_adj_456, n42_adj_457, n44_adj_458, n46_adj_459, 
        n47_adj_460, n48_adj_461, n50_adj_462, n52_adj_463, n54_adj_464, 
        n56_adj_465, n58_adj_466, n60_adj_467, n62_adj_468, n64_adj_469, 
        n38964, n22_adj_470, n24_adj_471, n26_adj_472, n28_adj_473, 
        n30_adj_474, n32_adj_475, n33_adj_476, n34_adj_477, n36_adj_478, 
        n38_adj_479, n40_adj_480, n42_adj_481, n44_adj_482, n45_adj_483, 
        n46_adj_484, n48_adj_485, n50_adj_486, n52_adj_487, n54_adj_488, 
        n56_adj_489, n58_adj_490, n60_adj_491, n62_adj_492, n64_adj_493, 
        n39975, n20_adj_494, n22_adj_495, n24_adj_496, n25_adj_497, 
        n26_adj_498, n28_adj_499, n30_adj_500, n31_adj_501, n32_adj_502, 
        n34_adj_503, n36_adj_504, n37_adj_505, n38_adj_506, n40_adj_507, 
        n42_adj_508, n43_adj_509, n44_adj_510, n46_adj_511, n48_adj_512, 
        n50_adj_513, n52_adj_514, n54_adj_515, n56_adj_516, n58_adj_517, 
        n60_adj_518, n62_adj_519, n64_adj_520, n37975, n18_adj_521, 
        n19_adj_522, n20_adj_523, n22_adj_524, n23_adj_525, n24_adj_526, 
        n26_adj_527, n28_adj_528, n29_adj_529, n30_adj_530, n32_adj_531, 
        n34_adj_532, n35_adj_533, n36_adj_534, n38_adj_535, n40_adj_536, 
        n41_adj_537, n42_adj_538, n44_adj_539, n46_adj_540, n48_adj_541, 
        n50_adj_542, n52_adj_543, n54_adj_544, n56_adj_545, n58_adj_546, 
        n60_adj_547, n62_adj_548, n64_adj_549, n37520, n16_adj_550, 
        n18_adj_551, n20_adj_552, n22_adj_553, n24_adj_554, n26_adj_555, 
        n27_adj_556, n28_adj_557, n30_adj_558, n31_adj_559, n32_adj_560, 
        n33_adj_561, n34_adj_562, n36_adj_563, n38_adj_564, n39_adj_565, 
        n40_adj_566, n42_adj_567, n44_adj_568, n46_adj_569, n48_adj_570, 
        n50_adj_571, n52_adj_572, n54_adj_573, n56_adj_574, n58_adj_575, 
        n60_adj_576, n62_adj_577, n64_adj_578, n14_adj_579, n42477, 
        n16_adj_580, n18_adj_581, n19_adj_582, n20_adj_583, n22_adj_584, 
        n24_adj_585, n25_adj_586, n26_adj_587, n28_adj_588, n30_adj_589, 
        n31_adj_590, n32_adj_591, n34_adj_592, n36_adj_593, n37_adj_594, 
        n38_adj_595, n40_adj_596, n42_adj_597, n44_adj_598, n46_adj_599, 
        n48_adj_600, n50_adj_601, n52_adj_602, n54_adj_603, n56_adj_604, 
        n58_adj_605, n60_adj_606, n62_adj_607, n64_adj_608, n38955, 
        n12_adj_609, n13_adj_610, n14_adj_611, n16_adj_612, n17_adj_613, 
        n18_adj_614, n20_adj_615, n22_adj_616, n23_adj_617, n24_adj_618, 
        n26_adj_619, n28_adj_620, n29_adj_621, n30_adj_622, n32_adj_623, 
        n34_adj_624, n35_adj_625, n36_adj_626, n38_adj_627, n40_adj_628, 
        n42_adj_629, n44_adj_630, n46_adj_631, n48_adj_632, n50_adj_633, 
        n52_adj_634, n54_adj_635, n56_adj_636, n58_adj_637, n60_adj_638, 
        n62_adj_639, n64_adj_640, n10_adj_641, n12_adj_642, n14_adj_643, 
        n16_adj_644, n18_adj_645, n20_adj_646, n21_adj_647, n22_adj_648, 
        n24_adj_649, n26_adj_650, n28_adj_651, n30_adj_652, n32_adj_653, 
        n33_adj_654, n34_adj_655, n36_adj_656, n38_adj_657, n40_adj_658, 
        n42_adj_659, n44_adj_660, n46_adj_661, n48_adj_662, n50_adj_663, 
        n52_adj_664, n54_adj_665, n56_adj_666, n58_adj_667, n60_adj_668, 
        n62_adj_669, n64_adj_670, n37965, n8_adj_671, n42476, n10_adj_672, 
        n12_adj_673, n13_adj_674, n14_adj_675, n16_adj_676, n18_adj_677, 
        n19_adj_678, n20_adj_679, n22_adj_680, n24_adj_681, n25_adj_682, 
        n26_adj_683, n28_adj_684, n30_adj_685, n31_adj_686, n32_adj_687, 
        n34_adj_688, n36_adj_689, n38_adj_690, n40_adj_691, n42_adj_692, 
        n44_adj_693, n46_adj_694, n48_adj_695, n50_adj_696, n52_adj_697, 
        n54_adj_698, n56_adj_699, n58_adj_700, n60_adj_701, n62_adj_702, 
        n64_adj_703, n37963, n6_adj_704, n8_adj_705, n10_adj_706, 
        n11_adj_707, n12_adj_708, n14_adj_709, n16_adj_710, n17_adj_711, 
        n18_adj_712, n20_adj_713, n21_adj_714, n22_adj_715, n24_adj_716, 
        n26_adj_717, n28_adj_718, n29_adj_719, n30_adj_720, n32_adj_721, 
        n34_adj_722, n36_adj_723, n38_adj_724, n40_adj_725, n42_adj_726, 
        n44_adj_727, n46_adj_728, n48_adj_729, n50_adj_730, n52_adj_731, 
        n54_adj_732, n56_adj_733, n58_adj_734, n60_adj_735, n62_adj_736, 
        n64_adj_737, n4_adj_738, n5_adj_739, n6_adj_740, n7_adj_741, 
        n8_adj_742, n9_adj_743, n10_adj_744, n11_adj_745, n12_adj_746, 
        n13_adj_747, n14_adj_748, n15_adj_749, n16_adj_750, n17_adj_751, 
        n18_adj_752, n19_adj_753, n20_adj_754, n21_adj_755, n22_adj_756, 
        n23_adj_757, n24_adj_758, n25_adj_759, n26_adj_760, n27_adj_761, 
        n28_adj_762, n29_adj_763, n30_adj_764, n31_adj_765, n32_adj_766, 
        n33_adj_767, n34_adj_768, n35_adj_769, n36_adj_770, n37_adj_771, 
        n38_adj_772, n39_adj_773, n40_adj_774, n42_adj_775, n43_adj_776, 
        n44_adj_777, n45_adj_778, n46_adj_779, n47_adj_780, n48_adj_781, 
        n49_adj_782, n50_adj_783, n52_adj_784, n53_adj_785, n54_adj_786, 
        n55_adj_787, n56_adj_788, n57_adj_789, n58_adj_790, n59_adj_791, 
        n60_adj_792, n61_adj_793, n62_adj_794, n37961, n37623, n42475, 
        n42474, n60_adj_795, n62_adj_796, n64_adj_797, n37616, n42473, 
        n42432, n36572, n42430, n38948, n62_adj_798, n37376, n36570, 
        n38944, n42472, n42471, n37949, n42470, n38939, n42469, 
        n64_adj_799, n37947, n37427, n38929, n38926, n37940, n38924, 
        n30962, n30878, n42468, n30881, n30884, n36562, n37932, 
        n37610, n62_adj_800, n30845, n42835, n62_adj_801, n30843, 
        n37603, n38910, n36558, n35972, n35970, n38908, n35968, 
        n37927, n42467, n37533, n35964, n37923, n38895, n37594, 
        n38892, n36556, clk_c_enable_831, n42833, n42832, n42831, 
        n42830, n38884, n42829, n42828, n42827, n37918, n42825, 
        n42824, n42823, n42822, n42821, n42820, n42819, n42818, 
        n42817, n42816, n42815, n42814, n38877, n37588, n42813, 
        n37586, n42812, n42811, n36994, n37908, n42810, n42809, 
        n42808, n42807, n42806, n42805, n36550, n36992, n42804, 
        n42803, n42802, n42801, n42800, n42799, n42798, n42797, 
        n37900, n42796, n42795, n42794, n37895, n42793, n42792, 
        n42791, n42790, n42789, n42788, n42787, n38866, n42786, 
        n42785, n42784, n36548, n42783, n42782, n42781, n37578, 
        n42780, n42779, n38862, n42778, n42777, n37576, n42776, 
        n42775, n42774, n42773, n36546, n37885, n42772, n42771, 
        n42769, n42768, n42767, n38857, n42766, n42765, n37879, 
        n42764, n37876, n42763, n42762, n42761, n42760, n42759, 
        n42758, n37446, n42757, n42756, n42755, n42754, n37571, 
        n42753, n37568, n42752, n37869, n36540, n42751, n42750, 
        n42749, n38847, n42748, n42747, n36538, n38842, n42746, 
        n38840, n42745, n37864, n42744, n37859, n42743, n42742, 
        n42466, n37854, n37455, n42465, n42741, n42464, n42740, 
        n42739, n42738, n42463, n42737, n42736, n42735, n42462, 
        n42461, n42734, n42733, n38835, n42732, n42460, n42731, 
        n42459, n39888, n42730, n42729, n42728, n42727, n42726, 
        n42725, n42724, n42458, n42723, n42722, n42721, n37845, 
        n42720, n37843, n42719, n42718, n42717, n42716, n38824, 
        n42715, n42714, n42713, n42712, n38820, n42711, n36500, 
        n42710, n38815, n42709, n42708, n42707, n42706, n42705, 
        n36498, n42704, n42703, n42702, n42701, n42700, n37558, 
        n42699, n42698, n42697, n38808, n42696, n42695, n42694, 
        n42693, n42692, n42691, n42690, n42689, n42688, n42687, 
        n36492, n36956, n42686, n42685, n42684, n37830, n38799, 
        n42683, n38797, n42682, n42681, n42680, n42679, n42678, 
        n42677, n39861, n42676, n42675, n42674, n42673, n42672, 
        n42671, n42670, n42669, n42668, n42667, n42666, n42665, 
        n37819, n42664, n42663, n42662, n42661, n42660, n42659, 
        n42658, n42657, n42656, n37812, n42655, n42654, n42653, 
        n42652, n42651, n37808, n42650, n36948, n42649, n42648, 
        n42647, n42646, n38786, n42645, n42644, n42643, n42642, 
        n36946, n38782, n42641, n42640, n42639, n42638, n42637, 
        n42636, n42635, n42634, n42633, n42632, n42631, n37795, 
        n38777, n42630, n42629, n37793, n42628, n42457, n37790, 
        n42456, n42627, n42626, n42455, n42625, n42624, n42623, 
        n42622, n42454, n42621, n42620, n42619, n42618, n42617, 
        n42616, n42615, n42614, n42453, n37781, n42613, n42452, 
        n42612, n42611, n42610, n42609, n42608, n42607, n42606, 
        n38765, n42451, n38763, n37774, n42605, n42604, n42603, 
        n37548, n42602, n37768, n42601, n42600, n42599, n39836, 
        n42598, n42597, n42596, n42450, n42595, n42594, n42449, 
        n42593, n42592, n42591, n37531, n37761, n42590, n42589, 
        n42588, n42587, n38752, n42586, n36926, n42585, n42584, 
        n42583, n42448, n42582, n42447, n38750, n42581, n42580, 
        n42579, n42578, n42577, n42576, n37752, n42575, n42574, 
        n42573, n37746, n42572, n42571, n37742, n42570, n42569, 
        n42568, n42567, n38741, n42566, n42565, n42564, n42563, 
        n42562, n42561, n42560, n42559, n42558, n42557, n42556, 
        n42555, n37738, n42554, n42553, n37733, n42552, n42551, 
        n37729, n42550, n42446, n37544, n42549, n42548, n36422, 
        n42547, n42546, n42545, n36918, n38728, n42544, n42543, 
        n42542, n38724, n36916, n42541, n37724, n38723, n42445, 
        n42540, n38721, n42539, n42444, n42538, n42537, n42536, 
        n42535, n42534, n42533, n37714, n42532, n42531, n42530, 
        n42529, n42528, n42527, n42526, n42525, n42524, n42523, 
        n42522, n42521, n42520, n37706, n42519, n42443, n42518, 
        n42517, n38711, n38709, n42516, n42515, n42514, n42513, 
        n38707, n42512, n42511, n37701, n38704, n42510, n42509, 
        n42508, n42507, n42506, n42505, n42504, n37691, n42503, 
        n42502, n42442, n35916, n35974, n42501, n42441, n42500, 
        n42499, n42498;
    
    VHI i2 (.Z(VCC_net));
    LUT4 div_4016_LessThan_2681_i29_2_lut (.A(n4093), .B(n125_adj_230), 
         .Z(n29_adj_529)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i29_2_lut.init = 16'h6666;
    FD1P3AX U_15___i508 (.D(\U[0] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i508.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1337_i48_3_lut_3_lut (.A(n2088), .B(n129), .C(n130_adj_233), 
         .Z(n48_adj_270)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1553_i51_2_lut_rep_1037 (.A(n2408), .B(n126), 
         .Z(n42736)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i51_2_lut_rep_1037.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i63_2_lut_rep_1051 (.A(n1916), .B(n123), 
         .Z(n42750)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i63_2_lut_rep_1051.init = 16'h6666;
    LUT4 i24861_3_lut (.A(\U[14] [0]), .B(\U[15] [0]), .C(i[0]), .Z(n40121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24861_3_lut.init = 16'hcaca;
    LUT4 i24860_3_lut (.A(\U[12] [0]), .B(\U[13] [0]), .C(i[0]), .Z(n40120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24860_3_lut.init = 16'hcaca;
    LUT4 i24933_3_lut (.A(\U[8] [5]), .B(\U[9] [5]), .C(i[0]), .Z(n40193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24933_3_lut.init = 16'hcaca;
    LUT4 i25176_3_lut (.A(\U[14] [21]), .B(\U[15] [21]), .C(i[0]), .Z(n40436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25176_3_lut.init = 16'hcaca;
    LUT4 i24859_3_lut (.A(\U[10] [0]), .B(\U[11] [0]), .C(i[0]), .Z(n40119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24859_3_lut.init = 16'hcaca;
    LUT4 i24858_3_lut (.A(\U[8] [0]), .B(\U[9] [0]), .C(i[0]), .Z(n40118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24858_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2762_i28_3_lut_3_lut (.A(n4200), .B(n111), .C(n123), 
         .Z(n28_adj_557)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i28_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_3206_i58_rep_18 (.BLUT(n37380), .ALUT(n37379), 
          .C0(n40074), .Z(n37378));
    LUT4 div_4016_LessThan_1226_i62_3_lut_3_lut (.A(n1916), .B(n123), .C(n60_adj_267), 
         .Z(n62_adj_268)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i62_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2841_i21_2_lut_rep_848 (.A(n4334), .B(n127_adj_231), 
         .Z(n42547)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i21_2_lut_rep_848.init = 16'h6666;
    LUT4 i24857_3_lut (.A(\U[6] [0]), .B(\U[7] [0]), .C(i[0]), .Z(n40117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24857_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_3206_i52 (.BLUT(n6_adj_740), .ALUT(n50_adj_783), 
          .C0(n40053), .Z(n52_adj_784));
    LUT4 div_4016_LessThan_1553_i48_3_lut_3_lut (.A(n2408), .B(n126), .C(n127_adj_231), 
         .Z(n48_adj_292)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25175_3_lut (.A(\U[12] [21]), .B(\U[13] [21]), .C(i[0]), .Z(n40435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25175_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i23_2_lut (.A(n4096), .B(n128_adj_232), 
         .Z(n23_adj_525)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i23_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i59_2_lut_rep_1052 (.A(n1918), .B(n125_adj_230), 
         .Z(n42751)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i59_2_lut_rep_1052.init = 16'h6666;
    LUT4 i25200_3_lut (.A(\U[2] [23]), .B(\U[3] [23]), .C(i[0]), .Z(n40460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25200_3_lut.init = 16'hcaca;
    LUT4 i24856_3_lut (.A(\U[4] [0]), .B(\U[5] [0]), .C(i[0]), .Z(n40116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24856_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1226_i56_3_lut_3_lut (.A(n1918), .B(n125_adj_230), 
         .C(n54_adj_263), .Z(n56_adj_265)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23606_3_lut_4_lut (.A(n4200), .B(n111), .C(n31_adj_559), .D(n42554), 
         .Z(n38866)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23606_3_lut_4_lut.init = 16'h0009;
    LUT4 i24855_3_lut (.A(\U[2] [0]), .B(\U[3] [0]), .C(i[0]), .Z(n40115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24855_3_lut.init = 16'hcaca;
    LUT4 i25779_3_lut_4_lut (.A(n1918), .B(n125_adj_230), .C(n55_adj_264), 
         .D(n42753), .Z(n37505)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25779_3_lut_4_lut.init = 16'hfff6;
    LUT4 i24932_3_lut (.A(\U[6] [5]), .B(\U[7] [5]), .C(i[0]), .Z(n40192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24932_3_lut.init = 16'hcaca;
    LUT4 i24854_3_lut (.A(\U[0] [0]), .B(\U[1] [0]), .C(i[0]), .Z(n40114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24854_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i32_3_lut_3_lut (.A(n4764), .B(n115_adj_223), 
         .C(n14_adj_709), .Z(n32_adj_721)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1226_i61_2_lut_rep_1053 (.A(n1917), .B(n124_adj_229), 
         .Z(n42752)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i61_2_lut_rep_1053.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i57_2_lut_rep_855 (.A(n4199), .B(n110_adj_220), 
         .Z(n42554)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i57_2_lut_rep_855.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i52_3_lut_3_lut (.A(n1917), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n52_adj_262)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24931_3_lut (.A(\U[4] [5]), .B(\U[5] [5]), .C(i[0]), .Z(n40191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24931_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_3206_i28 (.BLUT(n4_adj_738), .ALUT(n26_adj_760), 
          .C0(n39789), .Z(n28_adj_762));
    LUT4 i24930_3_lut (.A(\U[2] [5]), .B(\U[3] [5]), .C(i[0]), .Z(n40190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24930_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2762_i36_3_lut_3_lut (.A(n4199), .B(n110_adj_220), 
         .C(n28_adj_557), .Z(n36_adj_563)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i36_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 div_4016_LessThan_3137_i64 (.D0(n42_adj_726), .D1(n62_adj_736), 
            .SD(n39712), .Z(n64_adj_737));
    LUT4 div_4016_mux_5_i8_3_lut (.A(n5484), .B(n92_adj_210), .C(n5460), 
         .Z(n125_adj_230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i8_3_lut.init = 16'hcaca;
    L6MUX21 div_4016_LessThan_3137_i62 (.D0(n50_adj_730), .D1(n60_adj_735), 
            .SD(n39714), .Z(n62_adj_736));
    LUT4 i22334_3_lut_4_lut (.A(n2411), .B(n129), .C(n130_adj_233), .D(n2412), 
         .Z(n37594)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22334_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_mux_5_i19_3_lut (.A(n5473), .B(n81), .C(n5460), .Z(n114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i19_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_3137_i60 (.BLUT(n54_adj_732), .ALUT(n58_adj_734), 
          .C0(n39716), .Z(n60_adj_735));
    LUT4 i25666_4_lut_4_lut (.A(n42556), .B(n38835), .C(n46_adj_569), 
         .D(n22_adj_553), .Z(n48_adj_570)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25666_4_lut_4_lut.init = 16'hf4b0;
    PFUMX div_4016_LessThan_3137_i56 (.BLUT(n20_adj_713), .ALUT(n22_adj_715), 
          .C0(n39718), .Z(n56_adj_733));
    LUT4 i24929_3_lut (.A(\U[0] [5]), .B(\U[1] [5]), .C(i[0]), .Z(n40189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24929_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i17_3_lut (.A(n5475), .B(n83_adj_204), .C(n5460), 
         .Z(n116_adj_224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i17_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1553_i44_3_lut_3_lut (.A(n2411), .B(n129), .C(n130_adj_233), 
         .Z(n44_adj_290)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i44_3_lut_3_lut.init = 16'hd4d4;
    FD1P3AX U_15___i507 (.D(\U[0] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i507.GSR = "ENABLED";
    FD1P3AX U_15___i506 (.D(\U[0] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i506.GSR = "ENABLED";
    FD1P3AX U_15___i505 (.D(\U[0] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i505.GSR = "ENABLED";
    LUT4 i25571_4_lut_4_lut (.A(n42737), .B(n37578), .C(n58_adj_286), 
         .D(n46_adj_279), .Z(n60_adj_287)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25571_4_lut_4_lut.init = 16'hf4b0;
    FD1P3AX U_15___i504 (.D(\U[0] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i504.GSR = "ENABLED";
    FD1P3AX U_15___i503 (.D(\U[0] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i503.GSR = "ENABLED";
    L6MUX21 div_4016_LessThan_3206_i40 (.D0(n28_adj_762), .D1(n38_adj_772), 
            .SD(n39989), .Z(n40_adj_774));
    LUT4 i25787_3_lut_4_lut (.A(n4766), .B(n117), .C(n29_adj_719), .D(n42457), 
         .Z(n39602)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25787_3_lut_4_lut.init = 16'hfff6;
    LUT4 i23587_4_lut_4_lut (.A(n42556), .B(n38820), .C(n42555), .D(n42553), 
         .Z(n38847)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23587_4_lut_4_lut.init = 16'h00fb;
    PFUMX div_4016_LessThan_3206_i48 (.BLUT(n24_adj_758), .ALUT(n46_adj_779), 
          .C0(n40027), .Z(n48_adj_781));
    LUT4 i25199_3_lut (.A(\U[0] [23]), .B(\U[1] [23]), .C(i[0]), .Z(n40459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25199_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i502 (.D(\U[0] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i502.GSR = "ENABLED";
    FD1P3AX U_15___i501 (.D(\U[0] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i501.GSR = "ENABLED";
    FD1P3AX U_15___i500 (.D(\U[0] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i500.GSR = "ENABLED";
    FD1P3AX U_15___i499 (.D(\U[0] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i499.GSR = "ENABLED";
    FD1P3AX U_15___i498 (.D(\U[0] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i498.GSR = "ENABLED";
    FD1P3AX U_15___i497 (.D(\U[0] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i497.GSR = "ENABLED";
    FD1P3AX U_15___i496 (.D(\U[0] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i496.GSR = "ENABLED";
    FD1P3AX U_15___i495 (.D(\U[0] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i495.GSR = "ENABLED";
    FD1P3AX U_15___i494 (.D(\U[0] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i494.GSR = "ENABLED";
    FD1P3AX U_15___i493 (.D(\U[0] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i493.GSR = "ENABLED";
    FD1P3AX U_15___i492 (.D(\U[0] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i492.GSR = "ENABLED";
    FD1P3AX U_15___i491 (.D(\U[0] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i491.GSR = "ENABLED";
    FD1P3AX U_15___i490 (.D(\U[0] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i490.GSR = "ENABLED";
    FD1P3AX U_15___i489 (.D(\U[0] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i489.GSR = "ENABLED";
    FD1P3AX U_15___i488 (.D(\U[0] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i488.GSR = "ENABLED";
    FD1P3AX U_15___i487 (.D(\U[0] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i487.GSR = "ENABLED";
    FD1P3AX U_15___i486 (.D(\U[0] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i486.GSR = "ENABLED";
    FD1P3AX U_15___i485 (.D(\U[0] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i485.GSR = "ENABLED";
    FD1P3AX U_15___i484 (.D(\U[0] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i484.GSR = "ENABLED";
    FD1P3AX U_15___i483 (.D(\U[0] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i483.GSR = "ENABLED";
    LUT4 div_4016_mux_5_i20_3_lut (.A(n5472), .B(n80_adj_202), .C(n5460), 
         .Z(n113_adj_222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i20_3_lut.init = 16'hcaca;
    LUT4 i24921_3_lut (.A(\U[14] [4]), .B(\U[15] [4]), .C(i[0]), .Z(n40181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24921_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i482 (.D(\U[0] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i482.GSR = "ENABLED";
    LUT4 div_4016_LessThan_2762_i51_2_lut_rep_856 (.A(n4202), .B(n113_adj_222), 
         .Z(n42555)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i51_2_lut_rep_856.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i57_2_lut_rep_1054 (.A(n1919), .B(n126), 
         .Z(n42753)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i57_2_lut_rep_1054.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i54_3_lut_3_lut (.A(n1919), .B(n126), .C(n127_adj_231), 
         .Z(n54_adj_263)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1226_i51_2_lut_rep_1055 (.A(n1922), .B(n129), 
         .Z(n42754)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i51_2_lut_rep_1055.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i33_4_lut (.A(n4766), .B(n116_adj_224), 
         .C(n22256), .D(n4783), .Z(n33_adj_767)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i33_4_lut.init = 16'h663c;
    PFUMX div_4016_LessThan_3137_i50 (.BLUT(n26_adj_717), .ALUT(n48_adj_729), 
          .C0(n39678), .Z(n50_adj_730));
    LUT4 div_4016_mux_5_i21_3_lut (.A(n5471), .B(n79_adj_201), .C(n5460), 
         .Z(n112_adj_221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i21_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i481 (.D(\U[0] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i481.GSR = "ENABLED";
    FD1P3AX U_15___i480 (.D(\U[1] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i480.GSR = "ENABLED";
    FD1P3AX U_15___i479 (.D(\U[1] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i479.GSR = "ENABLED";
    FD1P3AX U_15___i478 (.D(\U[1] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i478.GSR = "ENABLED";
    FD1P3AX U_15___i477 (.D(\U[1] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i477.GSR = "ENABLED";
    FD1P3AX U_15___i476 (.D(\U[1] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i476.GSR = "ENABLED";
    FD1P3AX U_15___i475 (.D(\U[1] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i475.GSR = "ENABLED";
    FD1P3AX U_15___i474 (.D(\U[1] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i474.GSR = "ENABLED";
    FD1P3AX U_15___i473 (.D(\U[1] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i473.GSR = "ENABLED";
    FD1P3AX U_15___i472 (.D(\U[1] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i472.GSR = "ENABLED";
    FD1P3AX U_15___i471 (.D(\U[1] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i471.GSR = "ENABLED";
    FD1P3AX U_15___i470 (.D(\U[1] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i470.GSR = "ENABLED";
    FD1P3AX U_15___i469 (.D(\U[1] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i469.GSR = "ENABLED";
    FD1P3AX U_15___i468 (.D(\U[1] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i468.GSR = "ENABLED";
    FD1P3AX U_15___i467 (.D(\U[1] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i467.GSR = "ENABLED";
    FD1P3AX U_15___i466 (.D(\U[1] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i466.GSR = "ENABLED";
    FD1P3AX U_15___i465 (.D(\U[1] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i465.GSR = "ENABLED";
    FD1P3AX U_15___i464 (.D(\U[1] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i464.GSR = "ENABLED";
    FD1P3AX U_15___i463 (.D(\U[1] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i463.GSR = "ENABLED";
    FD1P3AX U_15___i462 (.D(\U[1] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i462.GSR = "ENABLED";
    FD1P3AX U_15___i461 (.D(\U[1] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i461.GSR = "ENABLED";
    FD1P3AX U_15___i460 (.D(\U[1] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i460.GSR = "ENABLED";
    FD1P3AX U_15___i459 (.D(\U[1] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i459.GSR = "ENABLED";
    FD1P3AX U_15___i458 (.D(\U[1] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i458.GSR = "ENABLED";
    FD1P3AX U_15___i457 (.D(\U[1] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i457.GSR = "ENABLED";
    FD1P3AX U_15___i456 (.D(\U[1] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i456.GSR = "ENABLED";
    FD1P3AX U_15___i455 (.D(\U[1] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i455.GSR = "ENABLED";
    FD1P3AX U_15___i454 (.D(\U[1] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i454.GSR = "ENABLED";
    FD1P3AX U_15___i453 (.D(\U[1] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i453.GSR = "ENABLED";
    FD1P3AX U_15___i452 (.D(\U[1] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i452.GSR = "ENABLED";
    FD1P3AX U_15___i451 (.D(\U[1] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i451.GSR = "ENABLED";
    FD1P3AX U_15___i450 (.D(\U[1] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i450.GSR = "ENABLED";
    FD1P3AX U_15___i449 (.D(\U[1] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[1] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i449.GSR = "ENABLED";
    FD1P3AX U_15___i448 (.D(\U[2] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i448.GSR = "ENABLED";
    FD1P3AX U_15___i447 (.D(\U[2] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i447.GSR = "ENABLED";
    FD1P3AX U_15___i446 (.D(\U[2] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i446.GSR = "ENABLED";
    FD1P3AX U_15___i445 (.D(\U[2] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i445.GSR = "ENABLED";
    FD1P3AX U_15___i444 (.D(\U[2] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i444.GSR = "ENABLED";
    FD1P3AX U_15___i443 (.D(\U[2] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i443.GSR = "ENABLED";
    FD1P3AX U_15___i442 (.D(\U[2] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i442.GSR = "ENABLED";
    FD1P3AX U_15___i441 (.D(\U[2] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i441.GSR = "ENABLED";
    FD1P3AX U_15___i440 (.D(\U[2] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i440.GSR = "ENABLED";
    FD1P3AX U_15___i439 (.D(\U[2] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i439.GSR = "ENABLED";
    FD1P3AX U_15___i438 (.D(\U[2] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i438.GSR = "ENABLED";
    FD1P3AX U_15___i437 (.D(\U[2] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i437.GSR = "ENABLED";
    FD1P3AX U_15___i436 (.D(\U[2] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i436.GSR = "ENABLED";
    FD1P3AX U_15___i435 (.D(\U[2] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i435.GSR = "ENABLED";
    FD1P3AX U_15___i434 (.D(\U[2] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i434.GSR = "ENABLED";
    FD1P3AX U_15___i433 (.D(\U[2] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i433.GSR = "ENABLED";
    FD1P3AX U_15___i432 (.D(\U[2] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i432.GSR = "ENABLED";
    FD1P3AX U_15___i431 (.D(\U[2] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i431.GSR = "ENABLED";
    FD1P3AX U_15___i430 (.D(\U[2] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i430.GSR = "ENABLED";
    FD1P3AX U_15___i429 (.D(\U[2] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i429.GSR = "ENABLED";
    FD1P3AX U_15___i428 (.D(\U[2] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i428.GSR = "ENABLED";
    FD1P3AX U_15___i427 (.D(\U[2] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i427.GSR = "ENABLED";
    FD1P3AX U_15___i426 (.D(\U[2] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i426.GSR = "ENABLED";
    FD1P3AX U_15___i425 (.D(\U[2] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i425.GSR = "ENABLED";
    FD1P3AX U_15___i424 (.D(\U[2] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i424.GSR = "ENABLED";
    FD1P3AX U_15___i423 (.D(\U[2] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i423.GSR = "ENABLED";
    FD1P3AX U_15___i422 (.D(\U[2] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i422.GSR = "ENABLED";
    FD1P3AX U_15___i421 (.D(\U[2] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i421.GSR = "ENABLED";
    FD1P3AX U_15___i420 (.D(\U[2] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i420.GSR = "ENABLED";
    FD1P3AX U_15___i419 (.D(\U[2] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i419.GSR = "ENABLED";
    FD1P3AX U_15___i418 (.D(\U[2] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i418.GSR = "ENABLED";
    FD1P3AX U_15___i417 (.D(\U[2] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[2] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i417.GSR = "ENABLED";
    FD1P3AX U_15___i416 (.D(\U[3] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i416.GSR = "ENABLED";
    FD1P3AX U_15___i415 (.D(\U[3] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i415.GSR = "ENABLED";
    FD1P3AX U_15___i414 (.D(\U[3] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i414.GSR = "ENABLED";
    FD1P3AX U_15___i413 (.D(\U[3] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i413.GSR = "ENABLED";
    FD1P3AX U_15___i412 (.D(\U[3] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i412.GSR = "ENABLED";
    FD1P3AX U_15___i411 (.D(\U[3] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i411.GSR = "ENABLED";
    FD1P3AX U_15___i410 (.D(\U[3] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i410.GSR = "ENABLED";
    FD1P3AX U_15___i409 (.D(\U[3] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i409.GSR = "ENABLED";
    FD1P3AX U_15___i408 (.D(\U[3] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i408.GSR = "ENABLED";
    FD1P3AX U_15___i407 (.D(\U[3] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i407.GSR = "ENABLED";
    FD1P3AX U_15___i406 (.D(\U[3] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i406.GSR = "ENABLED";
    FD1P3AX U_15___i405 (.D(\U[3] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i405.GSR = "ENABLED";
    FD1P3AX U_15___i404 (.D(\U[3] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i404.GSR = "ENABLED";
    LUT4 div_4016_mux_5_i6_3_lut (.A(n5486), .B(n94_adj_211), .C(n5460), 
         .Z(n127_adj_231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i6_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i403 (.D(\U[3] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i403.GSR = "ENABLED";
    FD1P3AX U_15___i402 (.D(\U[3] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i402.GSR = "ENABLED";
    IB U_in_pad_43 (.I(U_in[43]), .O(U_in_c_43));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_44 (.I(U_in[44]), .O(U_in_c_44));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_45 (.I(U_in[45]), .O(U_in_c_45));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_46 (.I(U_in[46]), .O(U_in_c_46));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i401 (.D(\U[3] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i401.GSR = "ENABLED";
    IB U_in_pad_47 (.I(U_in[47]), .O(U_in_c_47));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i400 (.D(\U[3] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i400.GSR = "ENABLED";
    IB U_in_pad_48 (.I(U_in[48]), .O(U_in_c_48));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_49 (.I(U_in[49]), .O(U_in_c_49));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_50 (.I(U_in[50]), .O(U_in_c_50));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_51 (.I(U_in[51]), .O(U_in_c_51));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_52 (.I(U_in[52]), .O(U_in_c_52));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_53 (.I(U_in[53]), .O(U_in_c_53));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_54 (.I(U_in[54]), .O(U_in_c_54));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    LUT4 div_4016_mux_5_i7_3_lut (.A(n5485), .B(n93), .C(n5460), .Z(n126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i7_3_lut.init = 16'hcaca;
    IB U_in_pad_55 (.I(U_in[55]), .O(U_in_c_55));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i399 (.D(\U[3] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i399.GSR = "ENABLED";
    FD1P3AX U_15___i398 (.D(\U[3] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i398.GSR = "ENABLED";
    FD1P3AX U_15___i397 (.D(\U[3] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i397.GSR = "ENABLED";
    FD1P3AX U_15___i396 (.D(\U[3] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i396.GSR = "ENABLED";
    FD1P3AX U_15___i395 (.D(\U[3] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i395.GSR = "ENABLED";
    FD1P3AX U_15___i394 (.D(\U[3] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i394.GSR = "ENABLED";
    FD1P3AX U_15___i393 (.D(\U[3] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i393.GSR = "ENABLED";
    FD1P3AX U_15___i392 (.D(\U[3] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i392.GSR = "ENABLED";
    FD1P3AX U_15___i391 (.D(\U[3] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i391.GSR = "ENABLED";
    FD1P3AX U_15___i390 (.D(\U[3] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i390.GSR = "ENABLED";
    FD1P3AX U_15___i389 (.D(\U[3] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i389.GSR = "ENABLED";
    FD1P3AX U_15___i388 (.D(\U[3] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i388.GSR = "ENABLED";
    FD1P3AX U_15___i387 (.D(\U[3] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i387.GSR = "ENABLED";
    FD1P3AX U_15___i386 (.D(\U[3] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i386.GSR = "ENABLED";
    FD1P3AX U_15___i385 (.D(\U[3] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[3] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i385.GSR = "ENABLED";
    FD1P3AX U_15___i384 (.D(U_0__31__N_967[383]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i384.GSR = "ENABLED";
    FD1P3AX U_15___i383 (.D(U_0__31__N_967[382]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i383.GSR = "ENABLED";
    FD1P3AX U_15___i382 (.D(U_0__31__N_967[381]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i382.GSR = "ENABLED";
    FD1P3AX U_15___i381 (.D(U_0__31__N_967[380]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i381.GSR = "ENABLED";
    FD1P3AX U_15___i380 (.D(U_0__31__N_967[379]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i380.GSR = "ENABLED";
    FD1P3AX U_15___i379 (.D(U_0__31__N_967[378]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i379.GSR = "ENABLED";
    FD1P3AX U_15___i378 (.D(U_0__31__N_967[377]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i378.GSR = "ENABLED";
    FD1P3AX U_15___i377 (.D(U_0__31__N_967[376]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i377.GSR = "ENABLED";
    FD1P3AX U_15___i376 (.D(U_0__31__N_967[375]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i376.GSR = "ENABLED";
    FD1P3AX U_15___i375 (.D(U_0__31__N_967[374]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i375.GSR = "ENABLED";
    FD1P3AX U_15___i374 (.D(U_0__31__N_967[373]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i374.GSR = "ENABLED";
    FD1P3AX U_15___i373 (.D(U_0__31__N_967[372]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i373.GSR = "ENABLED";
    FD1P3AX U_15___i372 (.D(U_0__31__N_967[371]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i372.GSR = "ENABLED";
    FD1P3AX U_15___i371 (.D(U_0__31__N_967[370]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i371.GSR = "ENABLED";
    FD1P3AX U_15___i370 (.D(U_0__31__N_967[369]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i370.GSR = "ENABLED";
    FD1P3AX U_15___i369 (.D(U_0__31__N_967[368]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i369.GSR = "ENABLED";
    FD1P3AX U_15___i368 (.D(U_0__31__N_967[367]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i368.GSR = "ENABLED";
    FD1P3AX U_15___i367 (.D(U_0__31__N_967[366]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i367.GSR = "ENABLED";
    FD1P3AX U_15___i366 (.D(U_0__31__N_967[365]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i366.GSR = "ENABLED";
    FD1P3AX U_15___i365 (.D(U_0__31__N_967[364]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i365.GSR = "ENABLED";
    FD1P3AX U_15___i364 (.D(U_0__31__N_967[363]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i364.GSR = "ENABLED";
    FD1P3AX U_15___i363 (.D(U_0__31__N_967[362]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i363.GSR = "ENABLED";
    FD1P3AX U_15___i362 (.D(U_0__31__N_967[361]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i362.GSR = "ENABLED";
    FD1P3AX U_15___i361 (.D(U_0__31__N_967[360]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i361.GSR = "ENABLED";
    FD1P3AX U_15___i360 (.D(U_0__31__N_967[359]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i360.GSR = "ENABLED";
    FD1P3AX U_15___i359 (.D(U_0__31__N_967[358]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i359.GSR = "ENABLED";
    FD1P3AX U_15___i358 (.D(U_0__31__N_967[357]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i358.GSR = "ENABLED";
    FD1P3AX U_15___i357 (.D(U_0__31__N_967[356]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i357.GSR = "ENABLED";
    FD1P3AX U_15___i356 (.D(U_0__31__N_967[355]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i356.GSR = "ENABLED";
    FD1P3AX U_15___i355 (.D(U_0__31__N_967[354]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i355.GSR = "ENABLED";
    FD1P3AX U_15___i354 (.D(U_0__31__N_967[353]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i354.GSR = "ENABLED";
    FD1P3AX U_15___i353 (.D(U_0__31__N_967[352]), .SP(clk_c_enable_831), 
            .CK(clk_c), .Q(\U[4] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i353.GSR = "ENABLED";
    FD1P3AX U_15___i352 (.D(\U[5] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i352.GSR = "ENABLED";
    FD1P3AX U_15___i351 (.D(\U[5] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i351.GSR = "ENABLED";
    FD1P3AX U_15___i350 (.D(\U[5] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i350.GSR = "ENABLED";
    FD1P3AX U_15___i349 (.D(\U[5] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i349.GSR = "ENABLED";
    FD1P3AX U_15___i348 (.D(\U[5] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i348.GSR = "ENABLED";
    FD1P3AX U_15___i347 (.D(\U[5] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i347.GSR = "ENABLED";
    FD1P3AX U_15___i346 (.D(\U[5] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i346.GSR = "ENABLED";
    FD1P3AX U_15___i345 (.D(\U[5] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i345.GSR = "ENABLED";
    FD1P3AX U_15___i344 (.D(\U[5] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i344.GSR = "ENABLED";
    FD1P3AX U_15___i343 (.D(\U[5] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i343.GSR = "ENABLED";
    FD1P3AX U_15___i342 (.D(\U[5] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i342.GSR = "ENABLED";
    FD1P3AX U_15___i341 (.D(\U[5] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i341.GSR = "ENABLED";
    FD1P3AX U_15___i340 (.D(\U[5] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i340.GSR = "ENABLED";
    FD1P3AX U_15___i339 (.D(\U[5] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i339.GSR = "ENABLED";
    FD1P3AX U_15___i338 (.D(\U[5] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i338.GSR = "ENABLED";
    FD1P3AX U_15___i337 (.D(\U[5] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i337.GSR = "ENABLED";
    FD1P3AX U_15___i336 (.D(\U[5] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i336.GSR = "ENABLED";
    FD1P3AX U_15___i335 (.D(\U[5] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i335.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1226_i50_3_lut_3_lut (.A(n1922), .B(n129), .C(n130_adj_233), 
         .Z(n50_adj_261)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3206_i13_4_lut (.A(n4776), .B(n126), .C(n22266), 
         .D(n4783), .Z(n13_adj_747)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i13_4_lut.init = 16'h663c;
    LUT4 i24920_3_lut (.A(\U[12] [4]), .B(\U[13] [4]), .C(i[0]), .Z(n40180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24920_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i334 (.D(\U[5] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i334.GSR = "ENABLED";
    FD1P3AX U_15___i333 (.D(\U[5] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i333.GSR = "ENABLED";
    FD1P3AX U_15___i332 (.D(\U[5] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i332.GSR = "ENABLED";
    FD1P3AX U_15___i331 (.D(\U[5] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i331.GSR = "ENABLED";
    FD1P3AX U_15___i330 (.D(\U[5] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i330.GSR = "ENABLED";
    FD1P3AX U_15___i329 (.D(\U[5] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i329.GSR = "ENABLED";
    FD1P3AX U_15___i328 (.D(\U[5] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i328.GSR = "ENABLED";
    FD1P3AX U_15___i327 (.D(\U[5] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i327.GSR = "ENABLED";
    FD1P3AX U_15___i326 (.D(\U[5] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i326.GSR = "ENABLED";
    FD1P3AX U_15___i325 (.D(\U[5] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i325.GSR = "ENABLED";
    FD1P3AX U_15___i324 (.D(\U[5] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i324.GSR = "ENABLED";
    FD1P3AX U_15___i323 (.D(\U[5] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i323.GSR = "ENABLED";
    FD1P3AX U_15___i322 (.D(\U[5] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i322.GSR = "ENABLED";
    FD1P3AX U_15___i321 (.D(\U[5] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[5] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i321.GSR = "ENABLED";
    FD1P3AX U_15___i320 (.D(\U[6] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i320.GSR = "ENABLED";
    FD1P3AX U_15___i319 (.D(\U[6] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i319.GSR = "ENABLED";
    FD1P3AX U_15___i318 (.D(\U[6] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i318.GSR = "ENABLED";
    FD1P3AX U_15___i317 (.D(\U[6] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i317.GSR = "ENABLED";
    FD1P3AX U_15___i316 (.D(\U[6] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i316.GSR = "ENABLED";
    FD1P3AX U_15___i315 (.D(\U[6] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i315.GSR = "ENABLED";
    FD1P3AX U_15___i314 (.D(\U[6] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i314.GSR = "ENABLED";
    FD1P3AX U_15___i313 (.D(\U[6] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i313.GSR = "ENABLED";
    FD1P3AX U_15___i312 (.D(\U[6] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i312.GSR = "ENABLED";
    FD1P3AX U_15___i311 (.D(\U[6] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i311.GSR = "ENABLED";
    FD1P3AX U_15___i310 (.D(\U[6] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i310.GSR = "ENABLED";
    FD1P3AX U_15___i309 (.D(\U[6] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i309.GSR = "ENABLED";
    FD1P3AX U_15___i308 (.D(\U[6] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i308.GSR = "ENABLED";
    FD1P3AX U_15___i307 (.D(\U[6] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i307.GSR = "ENABLED";
    FD1P3AX U_15___i306 (.D(\U[6] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i306.GSR = "ENABLED";
    FD1P3AX U_15___i305 (.D(\U[6] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i305.GSR = "ENABLED";
    FD1P3AX U_15___i304 (.D(\U[6] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i304.GSR = "ENABLED";
    FD1P3AX U_15___i303 (.D(\U[6] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i303.GSR = "ENABLED";
    FD1P3AX U_15___i302 (.D(\U[6] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i302.GSR = "ENABLED";
    FD1P3AX U_15___i301 (.D(\U[6] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i301.GSR = "ENABLED";
    FD1P3AX U_15___i300 (.D(\U[6] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i300.GSR = "ENABLED";
    FD1P3AX U_15___i299 (.D(\U[6] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i299.GSR = "ENABLED";
    FD1P3AX U_15___i298 (.D(\U[6] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i298.GSR = "ENABLED";
    FD1P3AX U_15___i297 (.D(\U[6] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i297.GSR = "ENABLED";
    FD1P3AX U_15___i296 (.D(\U[6] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i296.GSR = "ENABLED";
    FD1P3AX U_15___i295 (.D(\U[6] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i295.GSR = "ENABLED";
    FD1P3AX U_15___i294 (.D(\U[6] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i294.GSR = "ENABLED";
    FD1P3AX U_15___i293 (.D(\U[6] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i293.GSR = "ENABLED";
    FD1P3AX U_15___i292 (.D(\U[6] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i292.GSR = "ENABLED";
    FD1P3AX U_15___i291 (.D(\U[6] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i291.GSR = "ENABLED";
    FD1P3AX U_15___i290 (.D(\U[6] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i290.GSR = "ENABLED";
    FD1P3AX U_15___i289 (.D(\U[6] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[6] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i289.GSR = "ENABLED";
    FD1P3AX U_15___i288 (.D(\U[7] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i288.GSR = "ENABLED";
    FD1P3AX U_15___i287 (.D(\U[7] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i287.GSR = "ENABLED";
    FD1P3AX U_15___i286 (.D(\U[7] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i286.GSR = "ENABLED";
    FD1P3AX U_15___i285 (.D(\U[7] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i285.GSR = "ENABLED";
    FD1P3AX U_15___i284 (.D(\U[7] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i284.GSR = "ENABLED";
    FD1P3AX U_15___i283 (.D(\U[7] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i283.GSR = "ENABLED";
    FD1P3AX U_15___i282 (.D(\U[7] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i282.GSR = "ENABLED";
    FD1P3AX U_15___i281 (.D(\U[7] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i281.GSR = "ENABLED";
    FD1P3AX U_15___i280 (.D(\U[7] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i280.GSR = "ENABLED";
    FD1P3AX U_15___i279 (.D(\U[7] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i279.GSR = "ENABLED";
    FD1P3AX U_15___i278 (.D(\U[7] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i278.GSR = "ENABLED";
    FD1P3AX U_15___i277 (.D(\U[7] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i277.GSR = "ENABLED";
    FD1P3AX U_15___i276 (.D(\U[7] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i276.GSR = "ENABLED";
    FD1P3AX U_15___i275 (.D(\U[7] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i275.GSR = "ENABLED";
    FD1P3AX U_15___i274 (.D(\U[7] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i274.GSR = "ENABLED";
    FD1P3AX U_15___i273 (.D(\U[7] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i273.GSR = "ENABLED";
    FD1P3AX U_15___i272 (.D(\U[7] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i272.GSR = "ENABLED";
    IB U_in_pad_56 (.I(U_in[56]), .O(U_in_c_56));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_57 (.I(U_in[57]), .O(U_in_c_57));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_58 (.I(U_in[58]), .O(U_in_c_58));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_59 (.I(U_in[59]), .O(U_in_c_59));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_60 (.I(U_in[60]), .O(U_in_c_60));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_61 (.I(U_in[61]), .O(U_in_c_61));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_62 (.I(U_in[62]), .O(U_in_c_62));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_63 (.I(U_in[63]), .O(U_in_c_63));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_64 (.I(U_in[64]), .O(U_in_c_64));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_65 (.I(U_in[65]), .O(U_in_c_65));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_66 (.I(U_in[66]), .O(U_in_c_66));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_67 (.I(U_in[67]), .O(U_in_c_67));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_68 (.I(U_in[68]), .O(U_in_c_68));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_69 (.I(U_in[69]), .O(U_in_c_69));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_70 (.I(U_in[70]), .O(U_in_c_70));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_71 (.I(U_in[71]), .O(U_in_c_71));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    L6MUX21 div_4016_LessThan_3137_i42 (.D0(n30_adj_720), .D1(n40_adj_725), 
            .SD(n39634), .Z(n42_adj_726));
    FD1P3AX U_15___i271 (.D(\U[7] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i271.GSR = "ENABLED";
    LUT4 i24358_3_lut_4_lut (.A(n4764), .B(n115_adj_223), .C(n17_adj_711), 
         .D(n42455), .Z(n39618)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24358_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2841_i23_2_lut_rep_849 (.A(n4333), .B(n126), 
         .Z(n42548)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i23_2_lut_rep_849.init = 16'h6666;
    FD1P3AX U_15___i270 (.D(\U[7] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i270.GSR = "ENABLED";
    FD1P3AX U_15___i269 (.D(\U[7] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i269.GSR = "ENABLED";
    FD1P3AX U_15___i268 (.D(\U[7] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i268.GSR = "ENABLED";
    FD1P3AX U_15___i267 (.D(\U[7] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i267.GSR = "ENABLED";
    FD1P3AX U_15___i266 (.D(\U[7] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i266.GSR = "ENABLED";
    FD1P3AX U_15___i265 (.D(\U[7] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i265.GSR = "ENABLED";
    FD1P3AX U_15___i264 (.D(\U[7] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i264.GSR = "ENABLED";
    FD1P3AX U_15___i263 (.D(\U[7] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i263.GSR = "ENABLED";
    FD1P3AX U_15___i262 (.D(\U[7] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i262.GSR = "ENABLED";
    FD1P3AX U_15___i261 (.D(\U[7] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i261.GSR = "ENABLED";
    FD1P3AX U_15___i260 (.D(\U[7] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i260.GSR = "ENABLED";
    FD1P3AX U_15___i259 (.D(\U[7] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i259.GSR = "ENABLED";
    FD1P3AX U_15___i258 (.D(\U[7] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i258.GSR = "ENABLED";
    FD1P3AX U_15___i257 (.D(\U[7] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[7] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i257.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1446_i63_2_lut_rep_1038 (.A(n2243), .B(n121_adj_227), 
         .Z(n42737)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i63_2_lut_rep_1038.init = 16'h6666;
    FD1P3AX U_15___i256 (.D(\U[8] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i256.GSR = "ENABLED";
    LUT4 div_4016_LessThan_3206_i32_3_lut (.A(n114), .B(n113_adj_222), .C(n39_adj_773), 
         .Z(n32_adj_766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i32_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i31_2_lut_rep_758 (.A(n4767), .B(n118_adj_225), 
         .Z(n42457)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i31_2_lut_rep_758.init = 16'h6666;
    FD1P3AX U_15___i255 (.D(\U[8] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i255.GSR = "ENABLED";
    FD1P3AX U_15___i254 (.D(\U[8] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i254.GSR = "ENABLED";
    LUT4 div_4016_LessThan_3137_i16_3_lut_3_lut (.A(n4767), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n16_adj_710)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i16_3_lut_3_lut.init = 16'hd4d4;
    FD1P3AX U_15___i253 (.D(\U[8] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i253.GSR = "ENABLED";
    FD1P3AX U_15___i252 (.D(\U[8] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i252.GSR = "ENABLED";
    LUT4 i23632_2_lut_3_lut_4_lut (.A(n4333), .B(n126), .C(n127_adj_231), 
         .D(n4334), .Z(n38892)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23632_2_lut_3_lut_4_lut.init = 16'h9009;
    FD1P3AX U_15___i251 (.D(\U[8] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i251.GSR = "ENABLED";
    FD1P3AX U_15___i250 (.D(\U[8] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i250.GSR = "ENABLED";
    FD1P3AX U_15___i249 (.D(\U[8] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i249.GSR = "ENABLED";
    FD1P3AX U_15___i248 (.D(\U[8] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i248.GSR = "ENABLED";
    FD1P3AX U_15___i247 (.D(\U[8] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i247.GSR = "ENABLED";
    FD1P3AX U_15___i246 (.D(\U[8] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i246.GSR = "ENABLED";
    FD1P3AX U_15___i245 (.D(\U[8] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i245.GSR = "ENABLED";
    FD1P3AX U_15___i244 (.D(\U[8] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i244.GSR = "ENABLED";
    FD1P3AX U_15___i243 (.D(\U[8] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i243.GSR = "ENABLED";
    FD1P3AX U_15___i242 (.D(\U[8] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i242.GSR = "ENABLED";
    FD1P3AX U_15___i241 (.D(\U[8] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i241.GSR = "ENABLED";
    FD1P3AX U_15___i240 (.D(\U[8] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i240.GSR = "ENABLED";
    FD1P3AX U_15___i239 (.D(\U[8] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i239.GSR = "ENABLED";
    FD1P3AX U_15___i238 (.D(\U[8] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i238.GSR = "ENABLED";
    FD1P3AX U_15___i237 (.D(\U[8] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i237.GSR = "ENABLED";
    FD1P3AX U_15___i236 (.D(\U[8] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i236.GSR = "ENABLED";
    FD1P3AX U_15___i235 (.D(\U[8] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i235.GSR = "ENABLED";
    FD1P3AX U_15___i234 (.D(\U[8] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i234.GSR = "ENABLED";
    FD1P3AX U_15___i233 (.D(\U[8] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i233.GSR = "ENABLED";
    FD1P3AX U_15___i232 (.D(\U[8] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i232.GSR = "ENABLED";
    FD1P3AX U_15___i231 (.D(\U[8] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i231.GSR = "ENABLED";
    FD1P3AX U_15___i230 (.D(\U[8] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i230.GSR = "ENABLED";
    FD1P3AX U_15___i229 (.D(\U[8] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i229.GSR = "ENABLED";
    FD1P3AX U_15___i228 (.D(\U[8] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i228.GSR = "ENABLED";
    FD1P3AX U_15___i227 (.D(\U[8] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i227.GSR = "ENABLED";
    FD1P3AX U_15___i226 (.D(\U[8] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i226.GSR = "ENABLED";
    FD1P3AX U_15___i225 (.D(\U[8] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[8] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i225.GSR = "ENABLED";
    FD1P3AX U_15___i224 (.D(\U[9] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i224.GSR = "ENABLED";
    FD1P3AX U_15___i223 (.D(\U[9] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i223.GSR = "ENABLED";
    FD1P3AX U_15___i222 (.D(\U[9] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i222.GSR = "ENABLED";
    FD1P3AX U_15___i221 (.D(\U[9] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i221.GSR = "ENABLED";
    FD1P3AX U_15___i220 (.D(\U[9] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i220.GSR = "ENABLED";
    FD1P3AX U_15___i219 (.D(\U[9] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i219.GSR = "ENABLED";
    FD1P3AX U_15___i218 (.D(\U[9] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i218.GSR = "ENABLED";
    FD1P3AX U_15___i217 (.D(\U[9] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i217.GSR = "ENABLED";
    FD1P3AX U_15___i216 (.D(\U[9] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i216.GSR = "ENABLED";
    FD1P3AX U_15___i215 (.D(\U[9] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i215.GSR = "ENABLED";
    FD1P3AX U_15___i214 (.D(\U[9] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i214.GSR = "ENABLED";
    FD1P3AX U_15___i213 (.D(\U[9] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i213.GSR = "ENABLED";
    FD1P3AX U_15___i212 (.D(\U[9] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i212.GSR = "ENABLED";
    FD1P3AX U_15___i211 (.D(\U[9] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i211.GSR = "ENABLED";
    FD1P3AX U_15___i210 (.D(\U[9] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i210.GSR = "ENABLED";
    FD1P3AX U_15___i209 (.D(\U[9] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i209.GSR = "ENABLED";
    FD1P3AX U_15___i208 (.D(\U[9] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i208.GSR = "ENABLED";
    FD1P3AX U_15___i207 (.D(\U[9] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i207.GSR = "ENABLED";
    FD1P3AX U_15___i206 (.D(\U[9] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i206.GSR = "ENABLED";
    FD1P3AX U_15___i205 (.D(\U[9] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i205.GSR = "ENABLED";
    FD1P3AX U_15___i204 (.D(\U[9] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i204.GSR = "ENABLED";
    FD1P3AX U_15___i203 (.D(\U[9] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i203.GSR = "ENABLED";
    FD1P3AX U_15___i202 (.D(\U[9] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i202.GSR = "ENABLED";
    FD1P3AX U_15___i201 (.D(\U[9] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i201.GSR = "ENABLED";
    FD1P3AX U_15___i200 (.D(\U[9] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i200.GSR = "ENABLED";
    FD1P3AX U_15___i199 (.D(\U[9] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i199.GSR = "ENABLED";
    FD1P3AX U_15___i198 (.D(\U[9] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i198.GSR = "ENABLED";
    FD1P3AX U_15___i197 (.D(\U[9] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i197.GSR = "ENABLED";
    FD1P3AX U_15___i196 (.D(\U[9] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i196.GSR = "ENABLED";
    FD1P3AX U_15___i195 (.D(\U[9] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i195.GSR = "ENABLED";
    FD1P3AX U_15___i194 (.D(\U[9] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i194.GSR = "ENABLED";
    FD1P3AX U_15___i193 (.D(\U[9] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[9] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i193.GSR = "ENABLED";
    FD1P3AX U_15___i192 (.D(\U[10] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i192.GSR = "ENABLED";
    FD1P3AX U_15___i191 (.D(\U[10] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i191.GSR = "ENABLED";
    FD1P3AX U_15___i190 (.D(\U[10] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i190.GSR = "ENABLED";
    FD1P3AX U_15___i189 (.D(\U[10] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i189.GSR = "ENABLED";
    FD1P3AX U_15___i188 (.D(\U[10] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i188.GSR = "ENABLED";
    LUT4 div_4016_LessThan_2762_i44_3_lut_3_lut (.A(n4202), .B(n113_adj_222), 
         .C(n114), .Z(n44_adj_568)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25333_3_lut (.A(n40591), .B(n40592), .C(n9901), .Z(n5460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25333_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i1_3_lut (.A(n5491), .B(n99), .C(n5460), .Z(n132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i2_3_lut (.A(n5490), .B(n98_adj_214), .C(n5460), 
         .Z(n131_adj_234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i2_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i187 (.D(\U[10] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i187.GSR = "ENABLED";
    FD1P3AX U_15___i186 (.D(\U[10] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i186.GSR = "ENABLED";
    FD1P3AX U_15___i185 (.D(\U[10] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i185.GSR = "ENABLED";
    FD1P3AX U_15___i184 (.D(\U[10] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i184.GSR = "ENABLED";
    FD1P3AX U_15___i183 (.D(\U[10] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i183.GSR = "ENABLED";
    FD1P3AX U_15___i182 (.D(\U[10] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i182.GSR = "ENABLED";
    FD1P3AX U_15___i181 (.D(\U[10] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i181.GSR = "ENABLED";
    FD1P3AX U_15___i180 (.D(\U[10] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i180.GSR = "ENABLED";
    FD1P3AX U_15___i179 (.D(\U[10] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i179.GSR = "ENABLED";
    FD1P3AX U_15___i178 (.D(\U[10] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i178.GSR = "ENABLED";
    FD1P3AX U_15___i177 (.D(\U[10] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i177.GSR = "ENABLED";
    FD1P3AX U_15___i176 (.D(\U[10] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i176.GSR = "ENABLED";
    FD1P3AX U_15___i175 (.D(\U[10] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i175.GSR = "ENABLED";
    FD1P3AX U_15___i174 (.D(\U[10] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i174.GSR = "ENABLED";
    FD1P3AX U_15___i173 (.D(\U[10] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i173.GSR = "ENABLED";
    FD1P3AX U_15___i172 (.D(\U[10] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i172.GSR = "ENABLED";
    FD1P3AX U_15___i171 (.D(\U[10] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i171.GSR = "ENABLED";
    FD1P3AX U_15___i170 (.D(\U[10] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i170.GSR = "ENABLED";
    FD1P3AX U_15___i169 (.D(\U[10] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i169.GSR = "ENABLED";
    FD1P3AX U_15___i168 (.D(\U[10] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i168.GSR = "ENABLED";
    FD1P3AX U_15___i167 (.D(\U[10] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i167.GSR = "ENABLED";
    FD1P3AX U_15___i166 (.D(\U[10] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i166.GSR = "ENABLED";
    FD1P3AX U_15___i165 (.D(\U[10] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i165.GSR = "ENABLED";
    FD1P3AX U_15___i164 (.D(\U[10] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i164.GSR = "ENABLED";
    FD1P3AX U_15___i163 (.D(\U[10] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i163.GSR = "ENABLED";
    FD1P3AX U_15___i162 (.D(\U[10] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i162.GSR = "ENABLED";
    FD1P3AX U_15___i161 (.D(\U[10] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[10] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i161.GSR = "ENABLED";
    FD1P3AX U_15___i160 (.D(\U[11] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i160.GSR = "ENABLED";
    FD1P3AX U_15___i159 (.D(\U[11] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i159.GSR = "ENABLED";
    FD1P3AX U_15___i158 (.D(\U[11] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i158.GSR = "ENABLED";
    FD1P3AX U_15___i157 (.D(\U[11] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i157.GSR = "ENABLED";
    FD1P3AX U_15___i156 (.D(\U[11] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i156.GSR = "ENABLED";
    FD1P3AX U_15___i155 (.D(\U[11] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i155.GSR = "ENABLED";
    FD1P3AX U_15___i154 (.D(\U[11] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i154.GSR = "ENABLED";
    FD1P3AX U_15___i153 (.D(\U[11] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i153.GSR = "ENABLED";
    FD1P3AX U_15___i152 (.D(\U[11] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i152.GSR = "ENABLED";
    FD1P3AX U_15___i151 (.D(\U[11] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i151.GSR = "ENABLED";
    FD1P3AX U_15___i150 (.D(\U[11] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i150.GSR = "ENABLED";
    FD1P3AX U_15___i149 (.D(\U[11] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i149.GSR = "ENABLED";
    FD1P3AX U_15___i148 (.D(\U[11] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i148.GSR = "ENABLED";
    FD1P3AX U_15___i147 (.D(\U[11] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i147.GSR = "ENABLED";
    FD1P3AX U_15___i146 (.D(\U[11] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i146.GSR = "ENABLED";
    FD1P3AX U_15___i145 (.D(\U[11] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i145.GSR = "ENABLED";
    FD1P3AX U_15___i144 (.D(\U[11] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i144.GSR = "ENABLED";
    FD1P3AX U_15___i143 (.D(\U[11] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i143.GSR = "ENABLED";
    FD1P3AX U_15___i142 (.D(\U[11] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i142.GSR = "ENABLED";
    FD1P3AX U_15___i141 (.D(\U[11] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i141.GSR = "ENABLED";
    FD1P3AX U_15___i140 (.D(\U[11] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i140.GSR = "ENABLED";
    FD1P3AX U_15___i139 (.D(\U[11] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i139.GSR = "ENABLED";
    FD1P3AX U_15___i138 (.D(\U[11] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i138.GSR = "ENABLED";
    FD1P3AX U_15___i137 (.D(\U[11] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i137.GSR = "ENABLED";
    FD1P3AX U_15___i136 (.D(\U[11] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i136.GSR = "ENABLED";
    FD1P3AX U_15___i135 (.D(\U[11] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i135.GSR = "ENABLED";
    FD1P3AX U_15___i134 (.D(\U[11] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i134.GSR = "ENABLED";
    FD1P3AX U_15___i133 (.D(\U[11] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i133.GSR = "ENABLED";
    FD1P3AX U_15___i132 (.D(\U[11] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i132.GSR = "ENABLED";
    FD1P3AX U_15___i131 (.D(\U[11] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i131.GSR = "ENABLED";
    FD1P3AX U_15___i130 (.D(\U[11] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i130.GSR = "ENABLED";
    FD1P3AX U_15___i129 (.D(\U[11] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[11] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i129.GSR = "ENABLED";
    FD1P3AX U_15___i128 (.D(\U[12] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i128.GSR = "ENABLED";
    FD1P3AX U_15___i127 (.D(\U[12] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i127.GSR = "ENABLED";
    FD1P3AX U_15___i126 (.D(\U[12] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i126.GSR = "ENABLED";
    FD1P3AX U_15___i125 (.D(\U[12] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i125.GSR = "ENABLED";
    FD1P3IX x_3___i107 (.D(n5515), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i107.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1226_i53_2_lut_rep_1056 (.A(n1921), .B(n128_adj_232), 
         .Z(n42755)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i53_2_lut_rep_1056.init = 16'h6666;
    PFUMX div_4016_LessThan_3137_i40 (.BLUT(n32_adj_721), .ALUT(n38_adj_724), 
          .C0(n39636), .Z(n40_adj_725));
    LUT4 div_4016_LessThan_1446_i58_3_lut_3_lut (.A(n2243), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n58_adj_286)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i53_2_lut_rep_857 (.A(n4201), .B(n112_adj_221), 
         .Z(n42556)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i53_2_lut_rep_857.init = 16'h6666;
    LUT4 div_4016_LessThan_3137_i39_2_lut_rep_755 (.A(n4763), .B(n114), 
         .Z(n42454)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i39_2_lut_rep_755.init = 16'h6666;
    FD1P3AX U_15___i124 (.D(\U[12] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i124.GSR = "ENABLED";
    LUT4 div_4016_i3205_3_lut (.A(n893), .B(n22271), .C(n4783), .Z(n4883)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3205_3_lut.init = 16'hacac;
    LUT4 i25773_2_lut_3_lut_4_lut (.A(n1921), .B(n128_adj_232), .C(n124_adj_229), 
         .D(n1917), .Z(n37513)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25773_2_lut_3_lut_4_lut.init = 16'h6ff6;
    LUT4 div_4016_LessThan_3137_i25_2_lut_rep_759 (.A(n4770), .B(n121_adj_227), 
         .Z(n42458)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i25_2_lut_rep_759.init = 16'h6666;
    FD1P3AX U_15___i123 (.D(\U[12] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i123.GSR = "ENABLED";
    FD1P3AX U_15___i122 (.D(\U[12] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i122.GSR = "ENABLED";
    FD1P3AX U_15___i121 (.D(\U[12] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i121.GSR = "ENABLED";
    FD1P3AX U_15___i120 (.D(\U[12] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i120.GSR = "ENABLED";
    FD1P3AX U_15___i119 (.D(\U[12] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i119.GSR = "ENABLED";
    FD1P3AX U_15___i118 (.D(\U[12] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i118.GSR = "ENABLED";
    FD1P3AX U_15___i117 (.D(\U[12] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i117.GSR = "ENABLED";
    FD1P3AX U_15___i116 (.D(\U[12] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i116.GSR = "ENABLED";
    FD1P3AX U_15___i115 (.D(\U[12] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i115.GSR = "ENABLED";
    FD1P3AX U_15___i114 (.D(\U[12] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i114.GSR = "ENABLED";
    FD1P3AX U_15___i113 (.D(\U[12] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i113.GSR = "ENABLED";
    FD1P3AX U_15___i112 (.D(\U[12] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i112.GSR = "ENABLED";
    FD1P3AX U_15___i111 (.D(\U[12] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i111.GSR = "ENABLED";
    FD1P3AX U_15___i110 (.D(\U[12] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i110.GSR = "ENABLED";
    FD1P3AX U_15___i109 (.D(\U[12] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i109.GSR = "ENABLED";
    LUT4 i25955_4_lut (.A(n42572), .B(n42571), .C(n42573), .D(n38693), 
         .Z(n38711)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25955_4_lut.init = 16'hfffe;
    FD1P3AX U_15___i108 (.D(\U[12] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i108.GSR = "ENABLED";
    FD1P3AX U_15___i107 (.D(\U[12] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i107.GSR = "ENABLED";
    FD1P3AX U_15___i106 (.D(\U[12] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i106.GSR = "ENABLED";
    FD1P3AX U_15___i105 (.D(\U[12] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i105.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1113_i63_2_lut_rep_1057 (.A(n1748), .B(n124_adj_229), 
         .Z(n42756)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i63_2_lut_rep_1057.init = 16'h6666;
    IB U_in_pad_72 (.I(U_in[72]), .O(U_in_c_72));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_73 (.I(U_in[73]), .O(U_in_c_73));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i104 (.D(\U[12] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i104.GSR = "ENABLED";
    IB U_in_pad_74 (.I(U_in[74]), .O(U_in_c_74));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i103 (.D(\U[12] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i103.GSR = "ENABLED";
    IB U_in_pad_75 (.I(U_in[75]), .O(U_in_c_75));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_76 (.I(U_in[76]), .O(U_in_c_76));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_77 (.I(U_in[77]), .O(U_in_c_77));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i102 (.D(\U[12] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i102.GSR = "ENABLED";
    FD1P3AX U_15___i101 (.D(\U[12] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i101.GSR = "ENABLED";
    FD1P3AX U_15___i100 (.D(\U[12] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i100.GSR = "ENABLED";
    FD1P3AX U_15___i99 (.D(\U[12] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i99.GSR = "ENABLED";
    FD1P3AX U_15___i98 (.D(\U[12] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i98.GSR = "ENABLED";
    FD1P3AX U_15___i97 (.D(\U[12] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[12] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i97.GSR = "ENABLED";
    FD1P3AX U_15___i96 (.D(\U[13] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i96.GSR = "ENABLED";
    FD1P3AX U_15___i95 (.D(\U[13] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i95.GSR = "ENABLED";
    FD1P3AX U_15___i94 (.D(\U[13] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i94.GSR = "ENABLED";
    FD1P3AX U_15___i93 (.D(\U[13] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i93.GSR = "ENABLED";
    FD1P3AX U_15___i92 (.D(\U[13] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i92.GSR = "ENABLED";
    FD1P3AX U_15___i91 (.D(\U[13] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i91.GSR = "ENABLED";
    FD1P3AX U_15___i90 (.D(\U[13] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i90.GSR = "ENABLED";
    FD1P3AX U_15___i89 (.D(\U[13] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i89.GSR = "ENABLED";
    FD1P3AX U_15___i88 (.D(\U[13] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i88.GSR = "ENABLED";
    FD1P3AX U_15___i87 (.D(\U[13] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i87.GSR = "ENABLED";
    FD1P3AX U_15___i86 (.D(\U[13] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i86.GSR = "ENABLED";
    FD1P3AX U_15___i85 (.D(\U[13] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i85.GSR = "ENABLED";
    FD1P3AX U_15___i84 (.D(\U[13] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i84.GSR = "ENABLED";
    FD1P3AX U_15___i83 (.D(\U[13] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i83.GSR = "ENABLED";
    FD1P3AX U_15___i82 (.D(\U[13] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i82.GSR = "ENABLED";
    FD1P3AX U_15___i81 (.D(\U[13] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i81.GSR = "ENABLED";
    FD1P3AX U_15___i80 (.D(\U[13] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i80.GSR = "ENABLED";
    FD1P3AX U_15___i79 (.D(\U[13] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i79.GSR = "ENABLED";
    FD1P3AX U_15___i78 (.D(\U[13] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i78.GSR = "ENABLED";
    FD1P3AX U_15___i77 (.D(\U[13] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i77.GSR = "ENABLED";
    FD1P3AX U_15___i76 (.D(\U[13] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i76.GSR = "ENABLED";
    FD1P3AX U_15___i75 (.D(\U[13] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i75.GSR = "ENABLED";
    FD1P3AX U_15___i74 (.D(\U[13] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i74.GSR = "ENABLED";
    FD1P3AX U_15___i73 (.D(\U[13] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i73.GSR = "ENABLED";
    FD1P3AX U_15___i72 (.D(\U[13] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i72.GSR = "ENABLED";
    FD1P3AX U_15___i71 (.D(\U[13] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i71.GSR = "ENABLED";
    FD1P3AX U_15___i70 (.D(\U[13] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i70.GSR = "ENABLED";
    FD1P3AX U_15___i69 (.D(\U[13] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i69.GSR = "ENABLED";
    FD1P3AX U_15___i68 (.D(\U[13] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i68.GSR = "ENABLED";
    FD1P3AX U_15___i67 (.D(\U[13] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i67.GSR = "ENABLED";
    FD1P3AX U_15___i66 (.D(\U[13] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i66.GSR = "ENABLED";
    FD1P3AX U_15___i65 (.D(\U[13] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[13] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i65.GSR = "ENABLED";
    FD1P3AX U_15___i64 (.D(\U[14] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i64.GSR = "ENABLED";
    FD1P3AX U_15___i63 (.D(\U[14] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i63.GSR = "ENABLED";
    FD1P3AX U_15___i62 (.D(\U[14] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i62.GSR = "ENABLED";
    FD1P3AX U_15___i61 (.D(\U[14] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i61.GSR = "ENABLED";
    FD1P3AX U_15___i60 (.D(\U[14] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i60.GSR = "ENABLED";
    FD1P3AX U_15___i59 (.D(\U[14] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i59.GSR = "ENABLED";
    FD1P3AX U_15___i58 (.D(\U[14] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i58.GSR = "ENABLED";
    FD1P3AX U_15___i57 (.D(\U[14] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i57.GSR = "ENABLED";
    FD1P3AX U_15___i56 (.D(\U[14] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i56.GSR = "ENABLED";
    FD1P3AX U_15___i55 (.D(\U[14] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i55.GSR = "ENABLED";
    FD1P3AX U_15___i54 (.D(\U[14] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i54.GSR = "ENABLED";
    FD1P3AX U_15___i53 (.D(\U[14] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i53.GSR = "ENABLED";
    IB U_in_pad_78 (.I(U_in[78]), .O(U_in_c_78));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_79 (.I(U_in[79]), .O(U_in_c_79));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_80 (.I(U_in[80]), .O(U_in_c_80));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    FD1P3AX U_15___i52 (.D(\U[14] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i52.GSR = "ENABLED";
    IB U_in_pad_81 (.I(U_in[81]), .O(U_in_c_81));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    ALU54B lat_alu_4 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18615), .SIGNEDIB(n18688), .SIGNEDCIN(n18761), .A35(n18614), 
           .A34(n18613), .A33(n18612), .A32(n18611), .A31(n18610), .A30(n18609), 
           .A29(n18608), .A28(n18607), .A27(n18606), .A26(n18605), .A25(n18604), 
           .A24(n18603), .A23(n18602), .A22(n18601), .A21(n18600), .A20(n18599), 
           .A19(n18598), .A18(n18597), .A17(n18596), .A16(n18595), .A15(n18594), 
           .A14(n18593), .A13(n18592), .A12(n18591), .A11(n18590), .A10(n18589), 
           .A9(n18588), .A8(n18587), .A7(n18586), .A6(n18585), .A5(n18584), 
           .A4(n18583), .A3(n18582), .A2(n18581), .A1(n18580), .A0(n18579), 
           .B35(n18687), .B34(n18686), .B33(n18685), .B32(n18684), .B31(n18683), 
           .B30(n18682), .B29(n18681), .B28(n18680), .B27(n18679), .B26(n18678), 
           .B25(n18677), .B24(n18676), .B23(n18675), .B22(n18674), .B21(n18673), 
           .B20(n18672), .B19(n18671), .B18(n18670), .B17(n18669), .B16(n18668), 
           .B15(n18667), .B14(n18666), .B13(n18665), .B12(n18664), .B11(n18663), 
           .B10(n18662), .B9(n18661), .B8(n18660), .B7(n18659), .B6(n18658), 
           .B5(n18657), .B4(n18656), .B3(n18655), .B2(n18654), .B1(n18653), 
           .B0(n18652), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18651), .MA34(n18650), .MA33(n18649), .MA32(n18648), 
           .MA31(n18647), .MA30(n18646), .MA29(n18645), .MA28(n18644), 
           .MA27(n18643), .MA26(n18642), .MA25(n18641), .MA24(n18640), 
           .MA23(n18639), .MA22(n18638), .MA21(n18637), .MA20(n18636), 
           .MA19(n18635), .MA18(n18634), .MA17(n18633), .MA16(n18632), 
           .MA15(n18631), .MA14(n18630), .MA13(n18629), .MA12(n18628), 
           .MA11(n18627), .MA10(n18626), .MA9(n18625), .MA8(n18624), 
           .MA7(n18623), .MA6(n18622), .MA5(n18621), .MA4(n18620), .MA3(n18619), 
           .MA2(n18618), .MA1(n18617), .MA0(n18616), .MB35(n18724), 
           .MB34(n18723), .MB33(n18722), .MB32(n18721), .MB31(n18720), 
           .MB30(n18719), .MB29(n18718), .MB28(n18717), .MB27(n18716), 
           .MB26(n18715), .MB25(n18714), .MB24(n18713), .MB23(n18712), 
           .MB22(n18711), .MB21(n18710), .MB20(n18709), .MB19(n18708), 
           .MB18(n18707), .MB17(n18706), .MB16(n18705), .MB15(n18704), 
           .MB14(n18703), .MB13(n18702), .MB12(n18701), .MB11(n18700), 
           .MB10(n18699), .MB9(n18698), .MB8(n18697), .MB7(n18696), 
           .MB6(n18695), .MB5(n18694), .MB4(n18693), .MB3(n18692), .MB2(n18691), 
           .MB1(n18690), .MB0(n18689), .CIN53(n18760), .CIN52(n18759), 
           .CIN51(n18758), .CIN50(n18757), .CIN49(n18756), .CIN48(n18755), 
           .CIN47(n18754), .CIN46(n18753), .CIN45(n18752), .CIN44(n18751), 
           .CIN43(n18750), .CIN42(n18749), .CIN41(n18748), .CIN40(n18747), 
           .CIN39(n18746), .CIN38(n18745), .CIN37(n18744), .CIN36(n18743), 
           .CIN35(n18742), .CIN34(n18741), .CIN33(n18740), .CIN32(n18739), 
           .CIN31(n18738), .CIN30(n18737), .CIN29(n18736), .CIN28(n18735), 
           .CIN27(n18734), .CIN26(n18733), .CIN25(n18732), .CIN24(n18731), 
           .CIN23(n18730), .CIN22(n18729), .CIN21(n18728), .CIN20(n18727), 
           .CIN19(n18726), .CIN18(n18725), .CIN17(n177_adj_134), .CIN16(n178), 
           .CIN15(n179_adj_131), .CIN14(n180_adj_130), .CIN13(n181_adj_129), 
           .CIN12(n182_adj_128), .CIN11(n183), .CIN10(n184_adj_125), .CIN9(n185_adj_124), 
           .CIN8(n186_adj_123), .CIN7(n187_adj_122), .CIN6(n188), .CIN5(n189_adj_119), 
           .CIN4(n190_adj_118), .CIN3(n191_adj_117), .CIN2(n192_adj_116), 
           .CIN1(n193), .CIN0(n194_adj_114), .OP10(GND_net), .OP9(VCC_net), 
           .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), 
           .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), 
           .OP0(VCC_net), .R13(n163), .R12(n164_adj_149), .R11(n165_adj_148), 
           .R10(n166_adj_147), .R9(n167_adj_146), .R8(n168), .R7(n169_adj_143), 
           .R6(n170_adj_142), .R5(n171_adj_141), .R4(n172_adj_140), .R3(n173), 
           .R2(n174_adj_137), .R1(n175_adj_136), .R0(n176_adj_135));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[16:35])
    defparam lat_alu_4.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_4.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_4.REG_FLAG_CLK = "NONE";
    defparam lat_alu_4.REG_FLAG_CE = "CE0";
    defparam lat_alu_4.REG_FLAG_RST = "RST0";
    defparam lat_alu_4.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASK01 = "0x00000000000000";
    defparam lat_alu_4.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_4.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_4.CLK0_DIV = "ENABLED";
    defparam lat_alu_4.CLK1_DIV = "ENABLED";
    defparam lat_alu_4.CLK2_DIV = "ENABLED";
    defparam lat_alu_4.CLK3_DIV = "ENABLED";
    defparam lat_alu_4.MCPAT = "0x00000000000000";
    defparam lat_alu_4.MASKPAT = "0x00000000000000";
    defparam lat_alu_4.RNDPAT = "0x00000000000000";
    defparam lat_alu_4.GSR = "ENABLED";
    defparam lat_alu_4.RESETMODE = "SYNC";
    defparam lat_alu_4.MULT9_MODE = "DISABLED";
    defparam lat_alu_4.LEGACY = "DISABLED";
    FD1P3AX U_15___i51 (.D(\U[14] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i51.GSR = "ENABLED";
    FD1P3AX U_15___i50 (.D(\U[14] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i50.GSR = "ENABLED";
    FD1P3AX U_15___i49 (.D(\U[14] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i49.GSR = "ENABLED";
    FD1P3AX U_15___i48 (.D(\U[14] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i48.GSR = "ENABLED";
    FD1P3AX U_15___i47 (.D(\U[14] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i47.GSR = "ENABLED";
    FD1P3AX U_15___i46 (.D(\U[14] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i46.GSR = "ENABLED";
    LUT4 div_4016_LessThan_2841_i20_3_lut_3_lut (.A(n4333), .B(n126), .C(n127_adj_231), 
         .Z(n20_adj_583)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_3_i1_3_lut (.A(n5356), .B(n33_adj_193), .C(n5325), 
         .Z(n708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_4010_i1_4_lut (.A(n163_adj_11), .B(n36644), .C(n15805), .D(i[1]), 
         .Z(n5356)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i1_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut (.A(i[0]), .B(\y[3] [0]), .Z(n36644)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i24919_3_lut (.A(\U[10] [4]), .B(\U[11] [4]), .C(i[0]), .Z(n40179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24919_3_lut.init = 16'hcaca;
    FD1P3AX U_15___i45 (.D(\U[14] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i45.GSR = "ENABLED";
    FD1P3AX U_15___i44 (.D(\U[14] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i44.GSR = "ENABLED";
    FD1P3AX U_15___i43 (.D(\U[14] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i43.GSR = "ENABLED";
    FD1P3AX U_15___i42 (.D(\U[14] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i42.GSR = "ENABLED";
    FD1P3AX U_15___i41 (.D(\U[14] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i41.GSR = "ENABLED";
    FD1P3AX U_15___i40 (.D(\U[14] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i40.GSR = "ENABLED";
    FD1P3AX U_15___i39 (.D(\U[14] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i39.GSR = "ENABLED";
    FD1P3AX U_15___i38 (.D(\U[14] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i38.GSR = "ENABLED";
    FD1P3AX U_15___i37 (.D(\U[14] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i37.GSR = "ENABLED";
    FD1P3AX U_15___i36 (.D(\U[14] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i36.GSR = "ENABLED";
    FD1P3AX U_15___i35 (.D(\U[14] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i35.GSR = "ENABLED";
    FD1P3AX U_15___i34 (.D(\U[14] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i34.GSR = "ENABLED";
    FD1P3AX U_15___i33 (.D(\U[14] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[14] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i33.GSR = "ENABLED";
    FD1P3AX U_15___i32 (.D(\U[15] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i32.GSR = "ENABLED";
    FD1P3AX U_15___i31 (.D(\U[15] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i31.GSR = "ENABLED";
    FD1P3AX U_15___i30 (.D(\U[15] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i30.GSR = "ENABLED";
    FD1P3AX U_15___i29 (.D(\U[15] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i29.GSR = "ENABLED";
    FD1P3AX U_15___i28 (.D(\U[15] [27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i28.GSR = "ENABLED";
    FD1P3AX U_15___i27 (.D(\U[15] [26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i27.GSR = "ENABLED";
    FD1P3AX U_15___i26 (.D(\U[15] [25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i26.GSR = "ENABLED";
    FD1P3AX U_15___i25 (.D(\U[15] [24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i25.GSR = "ENABLED";
    FD1P3AX U_15___i24 (.D(\U[15] [23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i24.GSR = "ENABLED";
    FD1P3AX U_15___i23 (.D(\U[15] [22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i23.GSR = "ENABLED";
    FD1P3AX U_15___i22 (.D(\U[15] [21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i22.GSR = "ENABLED";
    FD1P3AX U_15___i21 (.D(\U[15] [20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i21.GSR = "ENABLED";
    FD1P3AX U_15___i20 (.D(\U[15] [19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i20.GSR = "ENABLED";
    FD1P3AX U_15___i19 (.D(\U[15] [18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i19.GSR = "ENABLED";
    FD1P3AX U_15___i18 (.D(\U[15] [17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i18.GSR = "ENABLED";
    FD1P3AX U_15___i17 (.D(\U[15] [16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i17.GSR = "ENABLED";
    FD1P3AX U_15___i16 (.D(\U[15] [15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i16.GSR = "ENABLED";
    FD1P3AX U_15___i15 (.D(\U[15] [14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i15.GSR = "ENABLED";
    FD1P3AX U_15___i14 (.D(\U[15] [13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i14.GSR = "ENABLED";
    FD1P3AX U_15___i13 (.D(\U[15] [12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i13.GSR = "ENABLED";
    FD1P3AX U_15___i12 (.D(\U[15] [11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i12.GSR = "ENABLED";
    FD1P3AX U_15___i11 (.D(\U[15] [10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i11.GSR = "ENABLED";
    FD1P3AX U_15___i10 (.D(\U[15] [9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i10.GSR = "ENABLED";
    FD1P3AX U_15___i9 (.D(\U[15] [8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i9.GSR = "ENABLED";
    FD1P3AX U_15___i8 (.D(\U[15] [7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i8.GSR = "ENABLED";
    FD1P3AX U_15___i7 (.D(\U[15] [6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i7.GSR = "ENABLED";
    FD1P3AX U_15___i6 (.D(\U[15] [5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i6.GSR = "ENABLED";
    FD1P3AX U_15___i5 (.D(\U[15] [4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i5.GSR = "ENABLED";
    FD1P3AX U_15___i4 (.D(\U[15] [3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i4.GSR = "ENABLED";
    FD1P3AX U_15___i3 (.D(\U[15] [2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i3.GSR = "ENABLED";
    FD1P3AX U_15___i2 (.D(\U[15] [1]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i2.GSR = "ENABLED";
    FD1P3AX y_3___i32 (.D(y_in_c_127), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i32.GSR = "ENABLED";
    LUT4 mux_4010_i32_4_lut (.A(n70_adj_87), .B(n36700), .C(n15805), .D(i[1]), 
         .Z(n5325)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i32_4_lut.init = 16'hca0a;
    LUT4 i24918_3_lut (.A(\U[8] [4]), .B(\U[9] [4]), .C(i[0]), .Z(n40178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24918_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i17_2_lut_rep_850 (.A(n4336), .B(n129), 
         .Z(n42549)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i17_2_lut_rep_850.init = 16'h6666;
    IB U_in_pad_82 (.I(U_in[82]), .O(U_in_c_82));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_83 (.I(U_in[83]), .O(U_in_c_83));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_84 (.I(U_in[84]), .O(U_in_c_84));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_85 (.I(U_in[85]), .O(U_in_c_85));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_86 (.I(U_in[86]), .O(U_in_c_86));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_87 (.I(U_in[87]), .O(U_in_c_87));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_88 (.I(U_in[88]), .O(U_in_c_88));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_89 (.I(U_in[89]), .O(U_in_c_89));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_90 (.I(U_in[90]), .O(U_in_c_90));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_91 (.I(U_in[91]), .O(U_in_c_91));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_92 (.I(U_in[92]), .O(U_in_c_92));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_93 (.I(U_in[93]), .O(U_in_c_93));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_94 (.I(U_in[94]), .O(U_in_c_94));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_95 (.I(U_in[95]), .O(U_in_c_95));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_96 (.I(U_in[96]), .O(U_in_c_96));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_97 (.I(U_in[97]), .O(U_in_c_97));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_98 (.I(U_in[98]), .O(U_in_c_98));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_99 (.I(U_in[99]), .O(U_in_c_99));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_100 (.I(U_in[100]), .O(U_in_c_100));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_101 (.I(U_in[101]), .O(U_in_c_101));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    LUT4 div_4016_LessThan_3137_i20_3_lut_3_lut (.A(n4770), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n20_adj_713)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i46_3_lut_3_lut (.A(n4201), .B(n112_adj_221), 
         .C(n44_adj_568), .Z(n46_adj_569)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2841_i16_3_lut_3_lut (.A(n4336), .B(n129), .C(n130_adj_233), 
         .Z(n16_adj_580)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_3_i8_3_lut (.A(n5349), .B(n26_adj_186), .C(n5325), 
         .Z(n887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i27_2_lut_rep_760 (.A(n4769), .B(n120), 
         .Z(n42459)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i27_2_lut_rep_760.init = 16'h6666;
    FD1P3IX x_3___i108 (.D(n5514), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i108.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_1 (.A(i[0]), .B(\y[3] [31]), .Z(n36700)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_1.init = 16'h8888;
    LUT4 div_4016_LessThan_1113_i62_3_lut_3_lut (.A(n1748), .B(n124_adj_229), 
         .C(n54_adj_254), .Z(n62_adj_259)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i62_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i49_2_lut_rep_858 (.A(n4203), .B(n114), 
         .Z(n42557)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i49_2_lut_rep_858.init = 16'h6666;
    LUT4 i23575_2_lut_3_lut_4_lut (.A(n4203), .B(n114), .C(n113_adj_222), 
         .D(n4202), .Z(n38835)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23575_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i24917_3_lut (.A(\U[6] [4]), .B(\U[7] [4]), .C(i[0]), .Z(n40177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24917_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1113_i61_2_lut_rep_1058 (.A(n1749), .B(n125_adj_230), 
         .Z(n42757)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i61_2_lut_rep_1058.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i47_2_lut_rep_859 (.A(n4204), .B(n115_adj_223), 
         .Z(n42558)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i47_2_lut_rep_859.init = 16'h6666;
    LUT4 i25191_3_lut (.A(\U[14] [22]), .B(\U[15] [22]), .C(i[0]), .Z(n40451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25191_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1113_i58_3_lut_3_lut (.A(n1749), .B(n125_adj_230), 
         .C(n56_adj_255), .Z(n58_adj_257)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i42_3_lut_3_lut (.A(n4204), .B(n115_adj_223), 
         .C(n24_adj_554), .Z(n42_adj_567)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25798_3_lut_4_lut (.A(n1749), .B(n125_adj_230), .C(n57_adj_256), 
         .D(n42758), .Z(n37482)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25798_3_lut_4_lut.init = 16'hfff6;
    PFUMX div_4016_LessThan_3137_i30 (.BLUT(n6_adj_704), .ALUT(n28_adj_718), 
          .C0(n39602), .Z(n30_adj_720));
    LUT4 i1_4_lut (.A(n36562), .B(n36572), .C(n36570), .D(i[3]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i23564_3_lut_4_lut (.A(n4204), .B(n115_adj_223), .C(n27_adj_556), 
         .D(n42560), .Z(n38824)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23564_3_lut_4_lut.init = 16'h0009;
    LUT4 i1_2_lut_adj_2 (.A(i[16]), .B(i[12]), .Z(n36562)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_2_lut_adj_2.init = 16'heeee;
    CCU2C equal_22116_32 (.A0(n5480), .B0(n5477), .C0(n5468), .D0(n5467), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n37339), 
          .S1(n37334));
    defparam equal_22116_32.INIT0 = 16'h0001;
    defparam equal_22116_32.INIT1 = 16'h0000;
    defparam equal_22116_32.INJECT1_0 = "YES";
    defparam equal_22116_32.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(i[1]), .B(i[0]), .C(i[3]), .D(i[2]), .Z(n9901)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[29:36])
    defparam i2_4_lut.init = 16'h965a;
    CCU2C equal_22116_31 (.A0(n5491), .B0(n5474), .C0(n5483), .D0(n5465), 
          .A1(n5490), .B1(n5475), .C1(n5485), .D1(n5471), .CIN(n37338), 
          .COUT(n37339));
    defparam equal_22116_31.INIT0 = 16'h0001;
    defparam equal_22116_31.INIT1 = 16'h0001;
    defparam equal_22116_31.INJECT1_0 = "YES";
    defparam equal_22116_31.INJECT1_1 = "YES";
    LUT4 div_4016_LessThan_1113_i59_2_lut_rep_1059 (.A(n1750), .B(n126), 
         .Z(n42758)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i59_2_lut_rep_1059.init = 16'h6666;
    LUT4 i1_4_lut_adj_3 (.A(i[31]), .B(n36556), .C(n36558), .D(i[18]), 
         .Z(n36572)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut_adj_3.init = 16'hfffe;
    LUT4 div_4016_LessThan_2762_i43_2_lut_rep_860 (.A(n4206), .B(n117), 
         .Z(n42559)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i43_2_lut_rep_860.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i38_3_lut_3_lut (.A(n4206), .B(n117), .C(n26_adj_555), 
         .Z(n38_adj_564)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1113_i56_3_lut_3_lut (.A(n1750), .B(n126), .C(n127_adj_231), 
         .Z(n56_adj_255)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25935_3_lut_4_lut (.A(n4206), .B(n117), .C(n39_adj_565), .D(n42561), 
         .Z(n38808)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25935_3_lut_4_lut.init = 16'hfff6;
    CCU2C equal_22116_29 (.A0(n5473), .B0(n5489), .C0(n5462), .D0(n5482), 
          .A1(n5478), .B1(n5487), .C1(n5461), .D1(n5476), .CIN(n37337), 
          .COUT(n37338));
    defparam equal_22116_29.INIT0 = 16'h0001;
    defparam equal_22116_29.INIT1 = 16'h0001;
    defparam equal_22116_29.INJECT1_0 = "YES";
    defparam equal_22116_29.INJECT1_1 = "YES";
    LUT4 i25876_4_lut (.A(n42568), .B(n38723), .C(n42569), .D(n38728), 
         .Z(n40104)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25876_4_lut.init = 16'hbfbb;
    LUT4 i1_4_lut_adj_4 (.A(i[20]), .B(i[10]), .C(i[23]), .D(i[8]), 
         .Z(n36570)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut_adj_4.init = 16'hfffe;
    LUT4 div_4016_LessThan_1446_i59_2_lut_rep_1039 (.A(n2245), .B(n123), 
         .Z(n42738)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i59_2_lut_rep_1039.init = 16'h6666;
    L6MUX21 div_4016_LessThan_3066_i62 (.D0(n52_adj_697), .D1(n60_adj_701), 
            .SD(n39525), .Z(n62_adj_702));
    CCU2C equal_22116_27 (.A0(n5470), .B0(n5481), .C0(n5484), .D0(n5486), 
          .A1(n5466), .B1(n5469), .C1(n5464), .D1(n5463), .CIN(n37336), 
          .COUT(n37337));
    defparam equal_22116_27.INIT0 = 16'h0001;
    defparam equal_22116_27.INIT1 = 16'h0001;
    defparam equal_22116_27.INJECT1_0 = "YES";
    defparam equal_22116_27.INJECT1_1 = "YES";
    LUT4 i25190_3_lut (.A(\U[12] [22]), .B(\U[13] [22]), .C(i[0]), .Z(n40450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25190_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_3066_i60 (.BLUT(n56_adj_699), .ALUT(n58_adj_700), 
          .C0(n39531), .Z(n60_adj_701));
    IB U_in_pad_102 (.I(U_in[102]), .O(U_in_c_102));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_103 (.I(U_in[103]), .O(U_in_c_103));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_104 (.I(U_in[104]), .O(U_in_c_104));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_105 (.I(U_in[105]), .O(U_in_c_105));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_106 (.I(U_in[106]), .O(U_in_c_106));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_107 (.I(U_in[107]), .O(U_in_c_107));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_108 (.I(U_in[108]), .O(U_in_c_108));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_109 (.I(U_in[109]), .O(U_in_c_109));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_110 (.I(U_in[110]), .O(U_in_c_110));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_111 (.I(U_in[111]), .O(U_in_c_111));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_112 (.I(U_in[112]), .O(U_in_c_112));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_113 (.I(U_in[113]), .O(U_in_c_113));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_114 (.I(U_in[114]), .O(U_in_c_114));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_115 (.I(U_in[115]), .O(U_in_c_115));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_116 (.I(U_in[116]), .O(U_in_c_116));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_117 (.I(U_in[117]), .O(U_in_c_117));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_118 (.I(U_in[118]), .O(U_in_c_118));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_119 (.I(U_in[119]), .O(U_in_c_119));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_120 (.I(U_in[120]), .O(U_in_c_120));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_121 (.I(U_in[121]), .O(U_in_c_121));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_122 (.I(U_in[122]), .O(U_in_c_122));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_123 (.I(U_in[123]), .O(U_in_c_123));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_124 (.I(U_in[124]), .O(U_in_c_124));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_125 (.I(U_in[125]), .O(U_in_c_125));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_126 (.I(U_in[126]), .O(U_in_c_126));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_127 (.I(U_in[127]), .O(U_in_c_127));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_128 (.I(U_in[128]), .O(U_in_c_128));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_129 (.I(U_in[129]), .O(U_in_c_129));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_130 (.I(U_in[130]), .O(U_in_c_130));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_131 (.I(U_in[131]), .O(U_in_c_131));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_132 (.I(U_in[132]), .O(U_in_c_132));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C equal_22116_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n5460), .B1(n5479), .C1(n5488), .D1(n5472), .COUT(n37336));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(115[14:29])
    defparam equal_22116_0.INIT0 = 16'h000F;
    defparam equal_22116_0.INIT1 = 16'h0001;
    defparam equal_22116_0.INJECT1_0 = "NO";
    defparam equal_22116_0.INJECT1_1 = "YES";
    LUT4 div_4016_LessThan_3206_i20_3_lut (.A(n120), .B(n103_adj_215), .C(n59_adj_791), 
         .Z(n20_adj_754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i20_3_lut.init = 16'hcaca;
    LUT4 i24916_3_lut (.A(\U[4] [4]), .B(\U[5] [4]), .C(i[0]), .Z(n40176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24916_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_5 (.A(i[15]), .B(i[17]), .Z(n36556)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_2_lut_adj_5.init = 16'heeee;
    FD1P3IX x_3___i109 (.D(n5513), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i109.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1446_i56_3_lut_3_lut (.A(n2245), .B(n123), .C(n48_adj_280), 
         .Z(n56_adj_285)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_6 (.A(i[24]), .B(i[4]), .Z(n36558)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_2_lut_adj_6.init = 16'heeee;
    LUT4 div_4016_LessThan_2762_i45_2_lut_rep_861 (.A(n4205), .B(n116_adj_224), 
         .Z(n42560)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i45_2_lut_rep_861.init = 16'h6666;
    LUT4 div_4016_LessThan_1113_i53_2_lut_rep_1060 (.A(n1753), .B(n129), 
         .Z(n42759)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i53_2_lut_rep_1060.init = 16'h6666;
    LUT4 div_4016_LessThan_1113_i52_3_lut_3_lut (.A(n1753), .B(n129), .C(n130_adj_233), 
         .Z(n52_adj_253)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3206_i17_4_lut (.A(n4774), .B(n124_adj_229), 
         .C(n22264), .D(n4783), .Z(n17_adj_751)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i17_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_3206_i42_3_lut (.A(n109_adj_219), .B(n108), .C(n49_adj_782), 
         .Z(n42_adj_775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i42_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_3066_i52 (.BLUT(n28_adj_684), .ALUT(n50_adj_696), 
          .C0(n39500), .Z(n52_adj_697));
    LUT4 div_4016_LessThan_1113_i55_2_lut_rep_1061 (.A(n1752), .B(n128_adj_232), 
         .Z(n42760)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i55_2_lut_rep_1061.init = 16'h6666;
    LUT4 i1_4_lut_adj_7 (.A(n36538), .B(n36550), .C(n36548), .D(n36532), 
         .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut_adj_7.init = 16'hfffe;
    LUT4 i1_2_lut_adj_8 (.A(i[28]), .B(i[19]), .Z(n36538)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_2_lut_adj_8.init = 16'heeee;
    LUT4 i24915_3_lut (.A(\U[2] [4]), .B(\U[3] [4]), .C(i[0]), .Z(n40175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24915_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1446_i55_2_lut_rep_1040 (.A(n2247), .B(n125_adj_230), 
         .Z(n42739)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i55_2_lut_rep_1040.init = 16'h6666;
    IB U_in_pad_133 (.I(U_in[133]), .O(U_in_c_133));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    ALU54B lat_alu_3 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18469), .SIGNEDIB(n18542), .SIGNEDCIN(GND_net), 
           .A35(n18468), .A34(n18467), .A33(n18466), .A32(n18465), .A31(n18464), 
           .A30(n18463), .A29(n18462), .A28(n18461), .A27(n18460), .A26(n18459), 
           .A25(n18458), .A24(n18457), .A23(n18456), .A22(n18455), .A21(n18454), 
           .A20(n18453), .A19(n18452), .A18(n18451), .A17(n18450), .A16(n18449), 
           .A15(n18448), .A14(n18447), .A13(n18446), .A12(n18445), .A11(n18444), 
           .A10(n18443), .A9(n18442), .A8(n18441), .A7(n18440), .A6(n18439), 
           .A5(n18438), .A4(n18437), .A3(n18436), .A2(n18435), .A1(n18434), 
           .A0(n18433), .B35(n18541), .B34(n18540), .B33(n18539), .B32(n18538), 
           .B31(n18537), .B30(n18536), .B29(n18535), .B28(n18534), .B27(n18533), 
           .B26(n18532), .B25(n18531), .B24(n18530), .B23(n18529), .B22(n18528), 
           .B21(n18527), .B20(n18526), .B19(n18525), .B18(n18524), .B17(n18523), 
           .B16(n18522), .B15(n18521), .B14(n18520), .B13(n18519), .B12(n18518), 
           .B11(n18517), .B10(n18516), .B9(n18515), .B8(n18514), .B7(n18513), 
           .B6(n18512), .B5(n18511), .B4(n18510), .B3(n18509), .B2(n18508), 
           .B1(n18507), .B0(n18506), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18505), .MA34(n18504), .MA33(n18503), .MA32(n18502), 
           .MA31(n18501), .MA30(n18500), .MA29(n18499), .MA28(n18498), 
           .MA27(n18497), .MA26(n18496), .MA25(n18495), .MA24(n18494), 
           .MA23(n18493), .MA22(n18492), .MA21(n18491), .MA20(n18490), 
           .MA19(n18489), .MA18(n18488), .MA17(n18487), .MA16(n18486), 
           .MA15(n18485), .MA14(n18484), .MA13(n18483), .MA12(n18482), 
           .MA11(n18481), .MA10(n18480), .MA9(n18479), .MA8(n18478), 
           .MA7(n18477), .MA6(n18476), .MA5(n18475), .MA4(n18474), .MA3(n18473), 
           .MA2(n18472), .MA1(n18471), .MA0(n18470), .MB35(n18578), 
           .MB34(n18577), .MB33(n18576), .MB32(n18575), .MB31(n18574), 
           .MB30(n18573), .MB29(n18572), .MB28(n18571), .MB27(n18570), 
           .MB26(n18569), .MB25(n18568), .MB24(n18567), .MB23(n18566), 
           .MB22(n18565), .MB21(n18564), .MB20(n18563), .MB19(n18562), 
           .MB18(n18561), .MB17(n18560), .MB16(n18559), .MB15(n18558), 
           .MB14(n18557), .MB13(n18556), .MB12(n18555), .MB11(n18554), 
           .MB10(n18553), .MB9(n18552), .MB8(n18551), .MB7(n18550), 
           .MB6(n18549), .MB5(n18548), .MB4(n18547), .MB3(n18546), .MB2(n18545), 
           .MB1(n18544), .MB0(n18543), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n18760), 
           .R52(n18759), .R51(n18758), .R50(n18757), .R49(n18756), .R48(n18755), 
           .R47(n18754), .R46(n18753), .R45(n18752), .R44(n18751), .R43(n18750), 
           .R42(n18749), .R41(n18748), .R40(n18747), .R39(n18746), .R38(n18745), 
           .R37(n18744), .R36(n18743), .R35(n18742), .R34(n18741), .R33(n18740), 
           .R32(n18739), .R31(n18738), .R30(n18737), .R29(n18736), .R28(n18735), 
           .R27(n18734), .R26(n18733), .R25(n18732), .R24(n18731), .R23(n18730), 
           .R22(n18729), .R21(n18728), .R20(n18727), .R19(n18726), .R18(n18725), 
           .R17(n177_adj_134), .R16(n178), .R15(n179_adj_131), .R14(n180_adj_130), 
           .R13(n181_adj_129), .R12(n182_adj_128), .R11(n183), .R10(n184_adj_125), 
           .R9(n185_adj_124), .R8(n186_adj_123), .R7(n187_adj_122), .R6(n188), 
           .R5(n189_adj_119), .R4(n190_adj_118), .R3(n191_adj_117), .R2(n192_adj_116), 
           .R1(n193), .R0(n194_adj_114), .SIGNEDR(n18761));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[16:35])
    defparam lat_alu_3.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_3.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_3.REG_FLAG_CLK = "NONE";
    defparam lat_alu_3.REG_FLAG_CE = "CE0";
    defparam lat_alu_3.REG_FLAG_RST = "RST0";
    defparam lat_alu_3.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASK01 = "0x00000000000000";
    defparam lat_alu_3.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_3.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_3.CLK0_DIV = "ENABLED";
    defparam lat_alu_3.CLK1_DIV = "ENABLED";
    defparam lat_alu_3.CLK2_DIV = "ENABLED";
    defparam lat_alu_3.CLK3_DIV = "ENABLED";
    defparam lat_alu_3.MCPAT = "0x00000000000000";
    defparam lat_alu_3.MASKPAT = "0x00000000000000";
    defparam lat_alu_3.RNDPAT = "0x00000000000000";
    defparam lat_alu_3.GSR = "ENABLED";
    defparam lat_alu_3.RESETMODE = "SYNC";
    defparam lat_alu_3.MULT9_MODE = "DISABLED";
    defparam lat_alu_3.LEGACY = "DISABLED";
    IB U_in_pad_134 (.I(U_in[134]), .O(U_in_c_134));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_135 (.I(U_in[135]), .O(U_in_c_135));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_136 (.I(U_in[136]), .O(U_in_c_136));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_137 (.I(U_in[137]), .O(U_in_c_137));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_138 (.I(U_in[138]), .O(U_in_c_138));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_139 (.I(U_in[139]), .O(U_in_c_139));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_140 (.I(U_in[140]), .O(U_in_c_140));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_141 (.I(U_in[141]), .O(U_in_c_141));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_142 (.I(U_in[142]), .O(U_in_c_142));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_143 (.I(U_in[143]), .O(U_in_c_143));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_144 (.I(U_in[144]), .O(U_in_c_144));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_145 (.I(U_in[145]), .O(U_in_c_145));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_146 (.I(U_in[146]), .O(U_in_c_146));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_147 (.I(U_in[147]), .O(U_in_c_147));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_148 (.I(U_in[148]), .O(U_in_c_148));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    L6MUX21 div_4016_LessThan_3066_i44 (.D0(n32_adj_687), .D1(n42_adj_692), 
            .SD(n39456), .Z(n44_adj_693));
    LUT4 i1_4_lut_adj_9 (.A(i[7]), .B(n36546), .C(n36540), .D(i[29]), 
         .Z(n36550)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut_adj_9.init = 16'hfffe;
    IB U_in_pad_149 (.I(U_in[149]), .O(U_in_c_149));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_150 (.I(U_in[150]), .O(U_in_c_150));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_151 (.I(U_in[151]), .O(U_in_c_151));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_152 (.I(U_in[152]), .O(U_in_c_152));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_153 (.I(U_in[153]), .O(U_in_c_153));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_154 (.I(U_in[154]), .O(U_in_c_154));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_155 (.I(U_in[155]), .O(U_in_c_155));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_156 (.I(U_in[156]), .O(U_in_c_156));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_157 (.I(U_in[157]), .O(U_in_c_157));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_158 (.I(U_in[158]), .O(U_in_c_158));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_159 (.I(U_in[159]), .O(U_in_c_159));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_160 (.I(U_in[160]), .O(U_in_c_160));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_161 (.I(U_in[161]), .O(U_in_c_161));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_162 (.I(U_in[162]), .O(U_in_c_162));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_163 (.I(U_in[163]), .O(U_in_c_163));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_164 (.I(U_in[164]), .O(U_in_c_164));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    LUT4 i1_4_lut_adj_10 (.A(i[13]), .B(i[26]), .C(i[25]), .D(i[27]), 
         .Z(n36548)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut_adj_10.init = 16'hfffe;
    LUT4 i1_2_lut_adj_11 (.A(i[30]), .B(i[14]), .Z(n36532)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_2_lut_adj_11.init = 16'heeee;
    LUT4 div_4016_LessThan_1113_i54_3_lut_3_lut (.A(n1752), .B(n128_adj_232), 
         .C(n52_adj_253), .Z(n54_adj_254)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i54_3_lut_3_lut.init = 16'hd4d4;
    IB U_in_pad_42 (.I(U_in[42]), .O(U_in_c_42));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    OB x_out_pad_122 (.I(x_out_c_122), .O(x_out[122]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    LUT4 div_4016_LessThan_2762_i24_3_lut_3_lut (.A(n4205), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n24_adj_554)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i41_2_lut_rep_862 (.A(n4207), .B(n118_adj_225), 
         .Z(n42561)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i41_2_lut_rep_862.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i26_3_lut_3_lut (.A(n4207), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n26_adj_555)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i26_3_lut_3_lut.init = 16'hd4d4;
    FD1P3IX x_3___i110 (.D(n5512), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i110.GSR = "ENABLED";
    LUT4 i24914_3_lut (.A(\U[0] [4]), .B(\U[1] [4]), .C(i[0]), .Z(n40174)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24914_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_12 (.A(i[22]), .B(i[5]), .C(i[9]), .D(i[6]), .Z(n36546)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_4_lut_adj_12.init = 16'hfffe;
    LUT4 div_4016_LessThan_1446_i52_3_lut_3_lut (.A(n2247), .B(n125_adj_230), 
         .C(n50_adj_281), .Z(n52_adj_283)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_998_i63_2_lut_rep_1062 (.A(n1577), .B(n125_adj_230), 
         .Z(n42761)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i63_2_lut_rep_1062.init = 16'h6666;
    LUT4 div_4016_LessThan_998_i60_3_lut_3_lut (.A(n1577), .B(n125_adj_230), 
         .C(n58_adj_249), .Z(n60_adj_250)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25670_4_lut_4_lut (.A(n42550), .B(n38877), .C(n56_adj_574), 
         .D(n20_adj_552), .Z(n58_adj_575)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25670_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2762_i64_4_lut_4_lut (.A(n42550), .B(n38862), 
         .C(n62_adj_577), .D(n52_adj_572), .Z(n64_adj_578)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i64_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25764_2_lut_3_lut_4_lut (.A(n4769), .B(n120), .C(n103_adj_215), 
         .D(n4752), .Z(n39718)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25764_2_lut_3_lut_4_lut.init = 16'h6ff6;
    LUT4 i25946_3_lut_4_lut (.A(n2247), .B(n125_adj_230), .C(n51_adj_282), 
         .D(n42741), .Z(n37568)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25946_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_2762_i35_2_lut_rep_863 (.A(n4210), .B(n121_adj_227), 
         .Z(n42562)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i35_2_lut_rep_863.init = 16'h6666;
    PFUMX div_4016_LessThan_3066_i42 (.BLUT(n34_adj_688), .ALUT(n40_adj_691), 
          .C0(n39458), .Z(n42_adj_692));
    MULT18X18D lat_mult_11 (.A17(\U[6] [17]), .A16(\U[6] [16]), .A15(\U[6] [15]), 
            .A14(\U[6] [14]), .A13(\U[6] [13]), .A12(\U[6] [12]), .A11(\U[6] [11]), 
            .A10(\U[6] [10]), .A9(\U[6] [9]), .A8(\U[6] [8]), .A7(\U[6] [7]), 
            .A6(\U[6] [6]), .A5(\U[6] [5]), .A4(\U[6] [4]), .A3(\U[6] [3]), 
            .A2(\U[6] [2]), .A1(\U[6] [1]), .A0(\U[6] [0]), .B17(\x[2] [31]), 
            .B16(\x[2] [31]), .B15(\x[2] [31]), .B14(\x[2] [31]), .B13(\x[2] [31]), 
            .B12(\x[2] [30]), .B11(\x[2] [29]), .B10(\x[2] [28]), .B9(\x[2] [27]), 
            .B8(\x[2] [26]), .B7(\x[2] [25]), .B6(\x[2] [24]), .B5(\x[2] [23]), 
            .B4(\x[2] [22]), .B3(\x[2] [21]), .B2(\x[2] [20]), .B1(\x[2] [19]), 
            .B0(\x[2] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19318), 
            .ROA16(n19317), .ROA15(n19316), .ROA14(n19315), .ROA13(n19314), 
            .ROA12(n19313), .ROA11(n19312), .ROA10(n19311), .ROA9(n19310), 
            .ROA8(n19309), .ROA7(n19308), .ROA6(n19307), .ROA5(n19306), 
            .ROA4(n19305), .ROA3(n19304), .ROA2(n19303), .ROA1(n19302), 
            .ROA0(n19301), .ROB17(n19336), .ROB16(n19335), .ROB15(n19334), 
            .ROB14(n19333), .ROB13(n19332), .ROB12(n19331), .ROB11(n19330), 
            .ROB10(n19329), .ROB9(n19328), .ROB8(n19327), .ROB7(n19326), 
            .ROB6(n19325), .ROB5(n19324), .ROB4(n19323), .ROB3(n19322), 
            .ROB2(n19321), .ROB1(n19320), .ROB0(n19319), .P35(n19373), 
            .P34(n19372), .P33(n19371), .P32(n19370), .P31(n19369), 
            .P30(n19368), .P29(n19367), .P28(n19366), .P27(n19365), 
            .P26(n19364), .P25(n19363), .P24(n19362), .P23(n19361), 
            .P22(n19360), .P21(n19359), .P20(n19358), .P19(n19357), 
            .P18(n19356), .P17(n19355), .P16(n19354), .P15(n19353), 
            .P14(n19352), .P13(n19351), .P12(n19350), .P11(n19349), 
            .P10(n19348), .P9(n19347), .P8(n19346), .P7(n19345), .P6(n19344), 
            .P5(n19343), .P4(n19342), .P3(n19341), .P2(n19340), .P1(n19339), 
            .P0(n19338), .SIGNEDP(n19337));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[19:38])
    defparam lat_mult_11.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTA_CE = "CE0";
    defparam lat_mult_11.REG_INPUTA_RST = "RST0";
    defparam lat_mult_11.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTB_CE = "CE0";
    defparam lat_mult_11.REG_INPUTB_RST = "RST0";
    defparam lat_mult_11.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTC_CE = "CE0";
    defparam lat_mult_11.REG_INPUTC_RST = "RST0";
    defparam lat_mult_11.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_11.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_11.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_11.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_11.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_11.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_11.CLK0_DIV = "ENABLED";
    defparam lat_mult_11.CLK1_DIV = "ENABLED";
    defparam lat_mult_11.CLK2_DIV = "ENABLED";
    defparam lat_mult_11.CLK3_DIV = "ENABLED";
    defparam lat_mult_11.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_11.GSR = "ENABLED";
    defparam lat_mult_11.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_11.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_11.MULT_BYPASS = "DISABLED";
    defparam lat_mult_11.RESETMODE = "SYNC";
    LUT4 i1_2_lut_adj_13 (.A(i[11]), .B(i[21]), .Z(n36540)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i1_2_lut_adj_13.init = 16'heeee;
    LUT4 div_4016_LessThan_2762_i30_3_lut_3_lut (.A(n4210), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n30_adj_558)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25831_3_lut_4_lut (.A(n1577), .B(n125_adj_230), .C(n59), .D(n42762), 
         .Z(n37462)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25831_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_mux_3_i2_3_lut (.A(n5355), .B(n32_adj_192), .C(n5325), 
         .Z(n893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i25189_3_lut (.A(\U[10] [22]), .B(\U[11] [22]), .C(i[0]), .Z(n40449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25189_3_lut.init = 16'hcaca;
    LUT4 i24906_3_lut (.A(\U[14] [3]), .B(\U[15] [3]), .C(i[0]), .Z(n40166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24906_3_lut.init = 16'hcaca;
    LUT4 i24905_3_lut (.A(\U[12] [3]), .B(\U[13] [3]), .C(i[0]), .Z(n40165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24905_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_998_i61_2_lut_rep_1063 (.A(n1578), .B(n126), 
         .Z(n42762)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i61_2_lut_rep_1063.init = 16'h6666;
    LUT4 div_4016_LessThan_998_i58_3_lut_3_lut (.A(n1578), .B(n126), .C(n127_adj_231), 
         .Z(n58_adj_249)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24904_3_lut (.A(\U[10] [3]), .B(\U[11] [3]), .C(i[0]), .Z(n40164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24904_3_lut.init = 16'hcaca;
    LUT4 mux_4010_i2_4_lut (.A(n160), .B(n36642), .C(n15805), .D(i[1]), 
         .Z(n5355)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i2_4_lut.init = 16'hca0a;
    FD1P3IX x_3___i111 (.D(n5511), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i111.GSR = "ENABLED";
    LUT4 i24369_2_lut_3_lut_4_lut (.A(n4763), .B(n114), .C(n113_adj_222), 
         .D(n4762), .Z(n39629)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24369_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_998_i57_2_lut_rep_1064 (.A(n1580), .B(n128_adj_232), 
         .Z(n42763)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i57_2_lut_rep_1064.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i63_2_lut_rep_851 (.A(n4196), .B(n107_adj_218), 
         .Z(n42550)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i63_2_lut_rep_851.init = 16'h6666;
    LUT4 div_4016_LessThan_1446_i57_2_lut_rep_1041 (.A(n2246), .B(n124_adj_229), 
         .Z(n42740)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i57_2_lut_rep_1041.init = 16'h6666;
    PFUMX div_4016_LessThan_3066_i32 (.BLUT(n8_adj_671), .ALUT(n30_adj_685), 
          .C0(n39424), .Z(n32_adj_687));
    LUT4 div_4016_LessThan_998_i56_3_lut_3_lut (.A(n1580), .B(n128_adj_232), 
         .C(n54_adj_247), .Z(n56_adj_248)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_14 (.A(i[0]), .B(\y[3] [1]), .Z(n36642)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_14.init = 16'h8888;
    FD1P3IX x_3___i112 (.D(n5510), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i112.GSR = "ENABLED";
    LUT4 i25937_3_lut_4_lut (.A(n4210), .B(n121_adj_227), .C(n33_adj_561), 
         .D(n42563), .Z(n38786)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25937_3_lut_4_lut.init = 16'hfff6;
    LUT4 i24903_3_lut (.A(\U[8] [3]), .B(\U[9] [3]), .C(i[0]), .Z(n40163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24903_3_lut.init = 16'hcaca;
    LUT4 i25188_3_lut (.A(\U[8] [22]), .B(\U[9] [22]), .C(i[0]), .Z(n40448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25188_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_998_i54_3_lut_3_lut (.A(n1581), .B(n129), .C(n130_adj_233), 
         .Z(n54_adj_247)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i37_2_lut_rep_864 (.A(n4209), .B(n120), 
         .Z(n42563)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i37_2_lut_rep_864.init = 16'h6666;
    LUT4 i22186_3_lut_4_lut (.A(n1581), .B(n129), .C(n130_adj_233), .D(n1582), 
         .Z(n37446)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22186_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_1446_i48_3_lut_3_lut (.A(n2246), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n48_adj_280)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_5_i31_3_lut (.A(n5461), .B(n69), .C(n5460), .Z(n102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i31_3_lut.init = 16'hcaca;
    FD1P3IX x_3___i113 (.D(n5509), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i113.GSR = "ENABLED";
    LUT4 i24902_3_lut (.A(\U[6] [3]), .B(\U[7] [3]), .C(i[0]), .Z(n40162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24902_3_lut.init = 16'hcaca;
    LUT4 i25561_4_lut_4_lut (.A(n42764), .B(n61), .C(n60_adj_244), .D(n54), 
         .Z(n62_adj_245)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25561_4_lut_4_lut.init = 16'hf4b0;
    PFUMX div_4016_LessThan_2993_i62 (.BLUT(n54_adj_665), .ALUT(n60_adj_668), 
          .C0(n39349), .Z(n62_adj_669));
    LUT4 i25883_4_lut (.A(n42585), .B(n42587), .C(n42586), .D(n38531), 
         .Z(n40096)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25883_4_lut.init = 16'hfffe;
    LUT4 i24901_3_lut (.A(\U[4] [3]), .B(\U[5] [3]), .C(i[0]), .Z(n40161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24901_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2762_i56_3_lut_3_lut (.A(n4196), .B(n107_adj_218), 
         .C(n54_adj_573), .Z(n56_adj_574)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3137_i35_2_lut_rep_756 (.A(n4765), .B(n116_adj_224), 
         .Z(n42455)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i35_2_lut_rep_756.init = 16'h6666;
    LUT4 i23271_4_lut (.A(n42596), .B(n42595), .C(n37_adj_505), .D(n38517), 
         .Z(n38531)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23271_4_lut.init = 16'h0001;
    LUT4 i24900_3_lut (.A(\U[2] [3]), .B(\U[3] [3]), .C(i[0]), .Z(n40160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24900_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2762_i59_2_lut_rep_852 (.A(n4198), .B(n109_adj_219), 
         .Z(n42551)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i59_2_lut_rep_852.init = 16'h6666;
    LUT4 i24899_3_lut (.A(\U[0] [3]), .B(\U[1] [3]), .C(i[0]), .Z(n40159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24899_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i14_3_lut_3_lut (.A(n4765), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n14_adj_709)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i14_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_2993_i58 (.BLUT(n26_adj_650), .ALUT(n56_adj_666), 
          .C0(n39351), .Z(n58_adj_667));
    LUT4 div_4016_LessThan_1446_i53_2_lut_rep_1042 (.A(n2248), .B(n126), 
         .Z(n42741)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i53_2_lut_rep_1042.init = 16'h6666;
    LUT4 div_4016_LessThan_881_i63_2_lut_rep_1065 (.A(n1403), .B(n126), 
         .Z(n42764)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i63_2_lut_rep_1065.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i32_3_lut_3_lut (.A(n4209), .B(n120), .C(n30_adj_558), 
         .Z(n32_adj_560)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_881_i60_3_lut_3_lut (.A(n1403), .B(n126), .C(n127_adj_231), 
         .Z(n60_adj_244)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i29_2_lut_rep_865 (.A(n4213), .B(n124_adj_229), 
         .Z(n42564)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i29_2_lut_rep_865.init = 16'h6666;
    LUT4 div_4016_LessThan_3137_i23_2_lut_rep_761 (.A(n4771), .B(n122_adj_228), 
         .Z(n42460)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i23_2_lut_rep_761.init = 16'h6666;
    LUT4 div_4016_LessThan_1446_i50_3_lut_3_lut (.A(n2248), .B(n126), .C(n127_adj_231), 
         .Z(n50_adj_281)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24313_2_lut_3_lut_4_lut (.A(n4771), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n4770), .Z(n39573)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24313_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2762_i20_3_lut_3_lut (.A(n4213), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n20_adj_552)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24891_3_lut (.A(\U[14] [2]), .B(\U[15] [2]), .C(i[0]), .Z(n40151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24891_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i33_2_lut_rep_757 (.A(n4766), .B(n117), 
         .Z(n42456)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i33_2_lut_rep_757.init = 16'h6666;
    LUT4 div_4016_LessThan_881_i56_3_lut_3_lut (.A(n1406), .B(n129), .C(n130_adj_233), 
         .Z(n56_adj_242)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22171_3_lut_4_lut (.A(n1406), .B(n129), .C(n130_adj_233), .D(n1407), 
         .Z(n37431)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22171_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_1446_i47_2_lut_rep_1043 (.A(n2251), .B(n129), 
         .Z(n42742)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i47_2_lut_rep_1043.init = 16'h6666;
    LUT4 div_4016_LessThan_881_i59_2_lut_rep_1066 (.A(n1405), .B(n128_adj_232), 
         .Z(n42765)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i59_2_lut_rep_1066.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i23_2_lut_rep_866 (.A(n4216), .B(n127_adj_231), 
         .Z(n42565)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i23_2_lut_rep_866.init = 16'h6666;
    LUT4 div_4016_LessThan_881_i58_3_lut_3_lut (.A(n1405), .B(n128_adj_232), 
         .C(n56_adj_242), .Z(n58_adj_243)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3206_i14_3_lut (.A(n119_adj_226), .B(n118_adj_225), 
         .C(n29_adj_763), .Z(n14_adj_748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i14_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i16_3_lut (.A(n5476), .B(n84), .C(n5460), .Z(n117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i16_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_762_i63_2_lut_rep_1067 (.A(n35972), .B(n127_adj_231), 
         .Z(n42766)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i63_2_lut_rep_1067.init = 16'h6666;
    FD1P3IX x_3___i114 (.D(n5508), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i114.GSR = "ENABLED";
    FD1P3JX i_i0_i0 (.D(n30843), .SP(clk_c_enable_831), .PD(clk_c_enable_708), 
            .CK(clk_c), .Q(i[0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i0.GSR = "ENABLED";
    LUT4 i24890_3_lut (.A(\U[12] [2]), .B(\U[13] [2]), .C(i[0]), .Z(n40150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24890_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1446_i46_3_lut_3_lut (.A(n2251), .B(n129), .C(n130_adj_233), 
         .Z(n46_adj_279)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_762_i62_3_lut_3_lut (.A(n35972), .B(n127_adj_231), 
         .C(n56_adj_237), .Z(n62_adj_240)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i62_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25187_3_lut (.A(\U[6] [22]), .B(\U[7] [22]), .C(i[0]), .Z(n40447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25187_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i28_3_lut_3_lut (.A(n4766), .B(n117), .C(n16_adj_710), 
         .Z(n28_adj_718)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_762_i59_2_lut_rep_1068 (.A(n1228), .B(n129), 
         .Z(n42767)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i59_2_lut_rep_1068.init = 16'h6666;
    LUT4 i24889_3_lut (.A(\U[10] [2]), .B(\U[11] [2]), .C(i[0]), .Z(n40149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24889_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i31_4_lut (.A(n4767), .B(n117), .C(n22257), 
         .D(n4783), .Z(n31_adj_765)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i31_4_lut.init = 16'h663c;
    LUT4 i25957_4_lut (.A(n42572), .B(n42571), .C(n42573), .D(n38684), 
         .Z(n38709)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25957_4_lut.init = 16'hfeff;
    L6MUX21 div_4016_LessThan_2993_i46 (.D0(n34_adj_655), .D1(n44_adj_660), 
            .SD(n39289), .Z(n46_adj_661));
    LUT4 div_4016_LessThan_2762_i25_2_lut_rep_867 (.A(n4215), .B(n126), 
         .Z(n42566)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i25_2_lut_rep_867.init = 16'h6666;
    LUT4 i24888_3_lut (.A(\U[8] [2]), .B(\U[9] [2]), .C(i[0]), .Z(n40148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24888_3_lut.init = 16'hcaca;
    LUT4 i23492_2_lut_3_lut_4_lut (.A(n4215), .B(n126), .C(n127_adj_231), 
         .D(n4216), .Z(n38752)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23492_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i24887_3_lut (.A(\U[6] [2]), .B(\U[7] [2]), .C(i[0]), .Z(n40147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24887_3_lut.init = 16'hcaca;
    LUT4 i23424_4_lut (.A(n42574), .B(n42576), .C(n42575), .D(n38668), 
         .Z(n38684)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23424_4_lut.init = 16'h1011;
    LUT4 i23408_4_lut (.A(n42577), .B(n41_adj_537), .C(n29_adj_529), .D(n38621), 
         .Z(n38668)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23408_4_lut.init = 16'h1011;
    FD1P3IX x_3___i115 (.D(n5507), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i115.GSR = "ENABLED";
    LUT4 div_4016_LessThan_762_i58_3_lut_3_lut (.A(n1228), .B(n129), .C(n130_adj_233), 
         .Z(n58_adj_238)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2598_i25_2_lut (.A(n3972), .B(n128_adj_232), 
         .Z(n25_adj_497)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i25_2_lut.init = 16'h6666;
    PFUMX div_4016_LessThan_2993_i44 (.BLUT(n36_adj_656), .ALUT(n42_adj_659), 
          .C0(n39291), .Z(n44_adj_660));
    LUT4 div_4016_LessThan_762_i61_2_lut_rep_1069 (.A(n1227), .B(n128_adj_232), 
         .Z(n42768)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i61_2_lut_rep_1069.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i22_3_lut_3_lut (.A(n4215), .B(n126), .C(n127_adj_231), 
         .Z(n22_adj_553)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24886_3_lut (.A(\U[4] [2]), .B(\U[5] [2]), .C(i[0]), .Z(n40146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24886_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_762_i60_3_lut_3_lut (.A(n1227), .B(n128_adj_232), 
         .C(n58_adj_238), .Z(n60_adj_239)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2762_i21_2_lut_rep_868 (.A(n4217), .B(n128_adj_232), 
         .Z(n42567)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i21_2_lut_rep_868.init = 16'h6666;
    LUT4 i25186_3_lut (.A(\U[4] [22]), .B(\U[5] [22]), .C(i[0]), .Z(n40446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25186_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2762_i61_2_lut_rep_853 (.A(n4197), .B(n108), 
         .Z(n42552)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i61_2_lut_rep_853.init = 16'h6666;
    LUT4 i24286_2_lut_3_lut_4_lut (.A(n4775), .B(n126), .C(n127_adj_231), 
         .D(n4776), .Z(n39546)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24286_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i23505_2_lut_3_lut_4_lut (.A(n4217), .B(n128_adj_232), .C(n124_adj_229), 
         .D(n4213), .Z(n38765)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23505_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_1446_i49_2_lut_rep_1044 (.A(n2250), .B(n128_adj_232), 
         .Z(n42743)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i49_2_lut_rep_1044.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i61_4_lut (.A(n4752), .B(n102), .C(n22242), 
         .D(n4783), .Z(n61_adj_793)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i61_4_lut.init = 16'h663c;
    LUT4 i22316_2_lut_3_lut_4_lut (.A(n2250), .B(n128_adj_232), .C(n124_adj_229), 
         .D(n2246), .Z(n37576)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22316_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i23481_3_lut_4_lut (.A(n4218), .B(n129), .C(n130_adj_233), .D(n4219), 
         .Z(n38741)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23481_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_3137_i19_2_lut_rep_762 (.A(n4773), .B(n124_adj_229), 
         .Z(n42461)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i19_2_lut_rep_762.init = 16'h6666;
    PFUMX div_4016_LessThan_2993_i34 (.BLUT(n10_adj_641), .ALUT(n32_adj_653), 
          .C0(n39257), .Z(n34_adj_655));
    LUT4 div_4016_mux_5_i14_3_lut (.A(n5478), .B(n86_adj_206), .C(n5460), 
         .Z(n119_adj_226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i14_3_lut.init = 16'hcaca;
    LUT4 i24885_3_lut (.A(\U[2] [2]), .B(\U[3] [2]), .C(i[0]), .Z(n40145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24885_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i15_3_lut (.A(n5477), .B(n85_adj_205), .C(n5460), 
         .Z(n118_adj_225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2762_i18_3_lut_3_lut (.A(n4218), .B(n129), .C(n130_adj_233), 
         .Z(n18_adj_551)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2598_i37_2_lut (.A(n3966), .B(n122_adj_228), 
         .Z(n37_adj_505)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i37_2_lut.init = 16'h6666;
    PFUMX div_4016_LessThan_2918_i62 (.BLUT(n56_adj_636), .ALUT(n60_adj_638), 
          .C0(n39184), .Z(n62_adj_639));
    LUT4 i25660_4_lut_4_lut (.A(n42568), .B(n38723), .C(n56_adj_545), 
         .D(n22_adj_524), .Z(n58_adj_546)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25660_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_i733_4_lut_4_lut (.A(n1048), .B(n130_adj_233), .C(n42835), 
         .D(n1078), .Z(n1228)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam div_4016_i733_4_lut_4_lut.init = 16'haa69;
    LUT4 div_4016_LessThan_1337_i63_2_lut_rep_1045 (.A(n2081), .B(n122_adj_228), 
         .Z(n42744)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i63_2_lut_rep_1045.init = 16'h6666;
    LUT4 i25878_3_lut_4_lut (.A(n1048), .B(n130_adj_233), .C(n42771), 
         .D(n42772), .Z(n37417)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;
    defparam i25878_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_641_i61_2_lut_rep_1072 (.A(n1047), .B(n129), 
         .Z(n42771)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_641_i61_2_lut_rep_1072.init = 16'h6666;
    LUT4 div_4016_LessThan_2681_i64_4_lut_4_lut (.A(n42568), .B(n38724), 
         .C(n62_adj_548), .D(n54_adj_544), .Z(n64_adj_549)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i64_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_3206_i29_4_lut (.A(n4768), .B(n118_adj_225), 
         .C(n22258), .D(n4783), .Z(n29_adj_763)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i29_4_lut.init = 16'h663c;
    LUT4 i24884_3_lut (.A(\U[0] [2]), .B(\U[1] [2]), .C(i[0]), .Z(n40144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24884_3_lut.init = 16'hcaca;
    LUT4 i24725_2_lut (.A(n39_adj_773), .B(n37_adj_771), .Z(n39985)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24725_2_lut.init = 16'h1111;
    LUT4 div_4016_LessThan_2681_i63_2_lut_rep_869 (.A(n4076), .B(n108), 
         .Z(n42568)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i63_2_lut_rep_869.init = 16'h6666;
    LUT4 div_4016_LessThan_2681_i56_3_lut_3_lut (.A(n4076), .B(n108), .C(n109_adj_219), 
         .Z(n56_adj_545)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1337_i60_3_lut_3_lut (.A(n2081), .B(n122_adj_228), 
         .C(n48_adj_270), .Z(n60_adj_276)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25755_3_lut (.A(n31_adj_765), .B(n29_adj_763), .C(n27_adj_761), 
         .Z(n39789)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25755_3_lut.init = 16'hfefe;
    LUT4 div_4016_LessThan_1337_i61_2_lut_rep_1046 (.A(n2082), .B(n123), 
         .Z(n42745)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i61_2_lut_rep_1046.init = 16'h6666;
    L6MUX21 div_4016_LessThan_2918_i48 (.D0(n36_adj_626), .D1(n46_adj_631), 
            .SD(n39131), .Z(n48_adj_632));
    LUT4 div_4016_i732_4_lut_4_lut (.A(n1047), .B(n129), .C(n60), .D(n1078), 
         .Z(n1227)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i732_4_lut_4_lut.init = 16'haa69;
    PFUMX div_4016_LessThan_2918_i58 (.BLUT(n28_adj_620), .ALUT(n30_adj_622), 
          .C0(n39186), .Z(n58_adj_637));
    LUT4 i23617_2_lut_3_lut_4_lut (.A(n4197), .B(n108), .C(n109_adj_219), 
         .D(n4198), .Z(n38877)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23617_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_641_i60_3_lut_3_lut (.A(n1047), .B(n129), .C(n130_adj_233), 
         .Z(n60_adj_236)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_641_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25656_4_lut_4_lut (.A(n42572), .B(n38704), .C(n48_adj_541), 
         .D(n24_adj_526), .Z(n50_adj_542)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25656_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_3137_i10_3_lut_3_lut (.A(n4773), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n10_adj_706)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1337_i58_3_lut_3_lut (.A(n2082), .B(n123), .C(n50_adj_271), 
         .Z(n58_adj_275)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1337_i57_2_lut_rep_1047 (.A(n2084), .B(n125_adj_230), 
         .Z(n42746)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i57_2_lut_rep_1047.init = 16'h6666;
    LUT4 div_4016_LessThan_641_i63_2_lut_rep_1073 (.A(n35970), .B(n128_adj_232), 
         .Z(n42772)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_641_i63_2_lut_rep_1073.init = 16'h9999;
    LUT4 div_4016_LessThan_3206_i27_4_lut (.A(n4769), .B(n119_adj_226), 
         .C(n22259), .D(n4783), .Z(n27_adj_761)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i27_4_lut.init = 16'h663c;
    LUT4 i23447_4_lut_4_lut (.A(n42572), .B(n38682), .C(n42573), .D(n42571), 
         .Z(n38707)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23447_4_lut_4_lut.init = 16'h0004;
    LUT4 i24876_3_lut (.A(\U[14] [1]), .B(\U[15] [1]), .C(i[0]), .Z(n40136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24876_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i13_3_lut (.A(n5479), .B(n87), .C(n5460), .Z(n120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i13_3_lut.init = 16'hcaca;
    LUT4 div_4016_i731_4_lut_4_lut (.A(n35970), .B(n128_adj_232), .C(n42432), 
         .D(n1078), .Z(n35972)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i731_4_lut_4_lut.init = 16'h5596;
    LUT4 div_4016_LessThan_641_i62_3_lut_3_lut (.A(n35970), .B(n128_adj_232), 
         .C(n60_adj_236), .Z(n62)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_641_i62_3_lut_3_lut.init = 16'he8e8;
    PFUMX div_4016_LessThan_2918_i46 (.BLUT(n38_adj_627), .ALUT(n44_adj_630), 
          .C0(n39133), .Z(n46_adj_631));
    LUT4 div_4016_LessThan_3137_i12_3_lut_3_lut (.A(n4775), .B(n126), .C(n127_adj_231), 
         .Z(n12_adj_708)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1337_i54_3_lut_3_lut (.A(n2084), .B(n125_adj_230), 
         .C(n52_adj_272), .Z(n54_adj_273)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i54_3_lut_3_lut.init = 16'hd4d4;
    FD1P3AX y_3___i31 (.D(y_in_c_126), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i31.GSR = "ENABLED";
    FD1P3AX y_3___i30 (.D(y_in_c_125), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i30.GSR = "ENABLED";
    FD1P3AX y_3___i29 (.D(y_in_c_124), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i29.GSR = "ENABLED";
    FD1P3AX y_3___i28 (.D(y_in_c_123), .SP(clk_c_enable_541), .CK(clk_c), 
            .Q(\y[3] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i28.GSR = "ENABLED";
    FD1P3AX y_3___i27 (.D(y_in_c_122), .SP(clk_c_enable_541), .CK(clk_c), 
            .Q(\y[3] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i27.GSR = "ENABLED";
    FD1P3AX y_3___i26 (.D(y_in_c_121), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i26.GSR = "ENABLED";
    FD1P3AX y_3___i25 (.D(y_in_c_120), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i25.GSR = "ENABLED";
    LUT4 i24875_3_lut (.A(\U[12] [1]), .B(\U[13] [1]), .C(i[0]), .Z(n40135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24875_3_lut.init = 16'hcaca;
    FD1P3AX y_3___i24 (.D(y_in_c_119), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i24.GSR = "ENABLED";
    FD1P3AX y_3___i23 (.D(y_in_c_118), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i23.GSR = "ENABLED";
    FD1P3AX y_3___i22 (.D(y_in_c_117), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i22.GSR = "ENABLED";
    FD1P3AX y_3___i21 (.D(y_in_c_116), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i21.GSR = "ENABLED";
    FD1P3AX y_3___i20 (.D(y_in_c_115), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i20.GSR = "ENABLED";
    FD1P3AX y_3___i19 (.D(y_in_c_114), .SP(clk_c_enable_541), .CK(clk_c), 
            .Q(\y[3] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i19.GSR = "ENABLED";
    FD1P3AX y_3___i18 (.D(y_in_c_113), .SP(clk_c_enable_541), .CK(clk_c), 
            .Q(\y[3] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i18.GSR = "ENABLED";
    FD1P3AX y_3___i17 (.D(y_in_c_112), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i17.GSR = "ENABLED";
    FD1P3AX y_3___i16 (.D(y_in_c_111), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i16.GSR = "ENABLED";
    FD1P3AX y_3___i15 (.D(y_in_c_110), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i15.GSR = "ENABLED";
    FD1P3AX y_3___i14 (.D(y_in_c_109), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i14.GSR = "ENABLED";
    FD1P3AX y_3___i13 (.D(y_in_c_108), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i13.GSR = "ENABLED";
    FD1P3AX y_3___i12 (.D(y_in_c_107), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i12.GSR = "ENABLED";
    FD1P3AX y_3___i11 (.D(y_in_c_106), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i11.GSR = "ENABLED";
    FD1P3AX y_3___i10 (.D(y_in_c_105), .SP(clk_c_enable_541), .CK(clk_c), 
            .Q(\y[3] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i10.GSR = "ENABLED";
    FD1P3AX y_3___i9 (.D(y_in_c_104), .SP(clk_c_enable_541), .CK(clk_c), 
            .Q(\y[3] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i9.GSR = "ENABLED";
    FD1P3AX y_3___i8 (.D(y_in_c_103), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i8.GSR = "ENABLED";
    FD1P3AX y_3___i7 (.D(y_in_c_102), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i7.GSR = "ENABLED";
    FD1P3AX y_3___i6 (.D(y_in_c_101), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i6.GSR = "ENABLED";
    FD1P3AX y_3___i5 (.D(y_in_c_100), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i5.GSR = "ENABLED";
    FD1P3AX y_3___i4 (.D(y_in_c_99), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i4.GSR = "ENABLED";
    FD1P3AX y_3___i3 (.D(y_in_c_98), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i3.GSR = "ENABLED";
    FD1P3AX y_3___i2 (.D(y_in_c_97), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i2.GSR = "ENABLED";
    FD1P3IX x_3___i116 (.D(n5506), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i116.GSR = "ENABLED";
    LUT4 div_4016_i610_4_lut_4_lut (.A(n35968), .B(n129), .C(n42430), 
         .D(n36422), .Z(n35970)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i610_4_lut_4_lut.init = 16'haa69;
    LUT4 div_4016_LessThan_2681_i59_2_lut_rep_870 (.A(n4078), .B(n110_adj_220), 
         .Z(n42569)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i59_2_lut_rep_870.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i45_4_lut (.A(n4760), .B(n110_adj_220), 
         .C(n22250), .D(n4783), .Z(n45_adj_778)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i45_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_518_i62_3_lut_3_lut (.A(n35968), .B(n129), .C(n130_adj_233), 
         .Z(n62_adj_796)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_518_i62_3_lut_3_lut.init = 16'he8e8;
    LUT4 i25185_3_lut (.A(\U[2] [22]), .B(\U[3] [22]), .C(i[0]), .Z(n40445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25185_3_lut.init = 16'hcaca;
    LUT4 i24275_3_lut_4_lut (.A(n4778), .B(n129), .C(n130_adj_233), .D(n4779), 
         .Z(n39535)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24275_3_lut_4_lut.init = 16'h9009;
    LUT4 i25184_3_lut (.A(\U[0] [22]), .B(\U[1] [22]), .C(i[0]), .Z(n40444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25184_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i43_4_lut (.A(n4761), .B(n111), .C(n22251), 
         .D(n4783), .Z(n43_adj_776)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i43_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_3137_i8_3_lut_3_lut (.A(n4778), .B(n129), .C(n130_adj_233), 
         .Z(n8_adj_705)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2681_i38_3_lut_3_lut (.A(n4078), .B(n110_adj_220), 
         .C(n30_adj_530), .Z(n38_adj_535)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25766_4_lut (.A(n42589), .B(n42588), .C(n42590), .D(n38562), 
         .Z(n38587)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25766_4_lut.init = 16'hfeff;
    LUT4 i25894_2_lut_3_lut_4_lut (.A(n864), .B(n130_adj_233), .C(n129), 
         .D(n35968), .Z(n40078)) /* synthesis lut_function=(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25894_2_lut_3_lut_4_lut.init = 16'hf66f;
    LUT4 i24874_3_lut (.A(\U[10] [1]), .B(\U[11] [1]), .C(i[0]), .Z(n40134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24874_3_lut.init = 16'hcaca;
    LUT4 div_4016_i611_4_lut_4_lut (.A(n864), .B(n130_adj_233), .C(n60_adj_162), 
         .D(n36422), .Z(n1047)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i611_4_lut_4_lut.init = 16'haa69;
    PFUMX div_4016_LessThan_2918_i36 (.BLUT(n12_adj_609), .ALUT(n34_adj_624), 
          .C0(n39099), .Z(n36_adj_626));
    LUT4 i25759_3_lut_4_lut (.A(n2084), .B(n125_adj_230), .C(n53), .D(n42748), 
         .Z(n37533)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25759_3_lut_4_lut.init = 16'hfff6;
    MULT18X18D lat_mult_10 (.A17(\U[6] [31]), .A16(\U[6] [31]), .A15(\U[6] [31]), 
            .A14(\U[6] [31]), .A13(\U[6] [31]), .A12(\U[6] [30]), .A11(\U[6] [29]), 
            .A10(\U[6] [28]), .A9(\U[6] [27]), .A8(\U[6] [26]), .A7(\U[6] [25]), 
            .A6(\U[6] [24]), .A5(\U[6] [23]), .A4(\U[6] [22]), .A3(\U[6] [21]), 
            .A2(\U[6] [20]), .A1(\U[6] [19]), .A0(\U[6] [18]), .B17(\x[2] [17]), 
            .B16(\x[2] [16]), .B15(\x[2] [15]), .B14(\x[2] [14]), .B13(\x[2] [13]), 
            .B12(\x[2] [12]), .B11(\x[2] [11]), .B10(\x[2] [10]), .B9(\x[2] [9]), 
            .B8(\x[2] [8]), .B7(\x[2] [7]), .B6(\x[2] [6]), .B5(\x[2] [5]), 
            .B4(\x[2] [4]), .B3(\x[2] [3]), .B2(\x[2] [2]), .B1(\x[2] [1]), 
            .B0(\x[2] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19245), 
            .ROA16(n19244), .ROA15(n19243), .ROA14(n19242), .ROA13(n19241), 
            .ROA12(n19240), .ROA11(n19239), .ROA10(n19238), .ROA9(n19237), 
            .ROA8(n19236), .ROA7(n19235), .ROA6(n19234), .ROA5(n19233), 
            .ROA4(n19232), .ROA3(n19231), .ROA2(n19230), .ROA1(n19229), 
            .ROA0(n19228), .ROB17(n19263), .ROB16(n19262), .ROB15(n19261), 
            .ROB14(n19260), .ROB13(n19259), .ROB12(n19258), .ROB11(n19257), 
            .ROB10(n19256), .ROB9(n19255), .ROB8(n19254), .ROB7(n19253), 
            .ROB6(n19252), .ROB5(n19251), .ROB4(n19250), .ROB3(n19249), 
            .ROB2(n19248), .ROB1(n19247), .ROB0(n19246), .P35(n19300), 
            .P34(n19299), .P33(n19298), .P32(n19297), .P31(n19296), 
            .P30(n19295), .P29(n19294), .P28(n19293), .P27(n19292), 
            .P26(n19291), .P25(n19290), .P24(n19289), .P23(n19288), 
            .P22(n19287), .P21(n19286), .P20(n19285), .P19(n19284), 
            .P18(n19283), .P17(n19282), .P16(n19281), .P15(n19280), 
            .P14(n19279), .P13(n19278), .P12(n19277), .P11(n19276), 
            .P10(n19275), .P9(n19274), .P8(n19273), .P7(n19272), .P6(n19271), 
            .P5(n19270), .P4(n19269), .P3(n19268), .P2(n19267), .P1(n19266), 
            .P0(n19265), .SIGNEDP(n19264));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[19:38])
    defparam lat_mult_10.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTA_CE = "CE0";
    defparam lat_mult_10.REG_INPUTA_RST = "RST0";
    defparam lat_mult_10.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTB_CE = "CE0";
    defparam lat_mult_10.REG_INPUTB_RST = "RST0";
    defparam lat_mult_10.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTC_CE = "CE0";
    defparam lat_mult_10.REG_INPUTC_RST = "RST0";
    defparam lat_mult_10.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_10.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_10.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_10.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_10.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_10.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_10.CLK0_DIV = "ENABLED";
    defparam lat_mult_10.CLK1_DIV = "ENABLED";
    defparam lat_mult_10.CLK2_DIV = "ENABLED";
    defparam lat_mult_10.CLK3_DIV = "ENABLED";
    defparam lat_mult_10.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_10.GSR = "ENABLED";
    defparam lat_mult_10.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_10.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_10.MULT_BYPASS = "DISABLED";
    defparam lat_mult_10.RESETMODE = "SYNC";
    MULT18X18D mult_4003_mult_2 (.A17(\U[6] [17]), .A16(\U[6] [16]), .A15(\U[6] [15]), 
            .A14(\U[6] [14]), .A13(\U[6] [13]), .A12(\U[6] [12]), .A11(\U[6] [11]), 
            .A10(\U[6] [10]), .A9(\U[6] [9]), .A8(\U[6] [8]), .A7(\U[6] [7]), 
            .A6(\U[6] [6]), .A5(\U[6] [5]), .A4(\U[6] [4]), .A3(\U[6] [3]), 
            .A2(\U[6] [2]), .A1(\U[6] [1]), .A0(\U[6] [0]), .B17(\x[2] [17]), 
            .B16(\x[2] [16]), .B15(\x[2] [15]), .B14(\x[2] [14]), .B13(\x[2] [13]), 
            .B12(\x[2] [12]), .B11(\x[2] [11]), .B10(\x[2] [10]), .B9(\x[2] [9]), 
            .B8(\x[2] [8]), .B7(\x[2] [7]), .B6(\x[2] [6]), .B5(\x[2] [5]), 
            .B4(\x[2] [4]), .B3(\x[2] [3]), .B2(\x[2] [2]), .B1(\x[2] [1]), 
            .B0(\x[2] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19172), 
            .ROA16(n19171), .ROA15(n19170), .ROA14(n19169), .ROA13(n19168), 
            .ROA12(n19167), .ROA11(n19166), .ROA10(n19165), .ROA9(n19164), 
            .ROA8(n19163), .ROA7(n19162), .ROA6(n19161), .ROA5(n19160), 
            .ROA4(n19159), .ROA3(n19158), .ROA2(n19157), .ROA1(n19156), 
            .ROA0(n19155), .ROB17(n19190), .ROB16(n19189), .ROB15(n19188), 
            .ROB14(n19187), .ROB13(n19186), .ROB12(n19185), .ROB11(n19184), 
            .ROB10(n19183), .ROB9(n19182), .ROB8(n19181), .ROB7(n19180), 
            .ROB6(n19179), .ROB5(n19178), .ROB4(n19177), .ROB3(n19176), 
            .ROB2(n19175), .ROB1(n19174), .ROB0(n19173), .P35(n19227), 
            .P34(n19226), .P33(n19225), .P32(n19224), .P31(n19223), 
            .P30(n19222), .P29(n19221), .P28(n19220), .P27(n19219), 
            .P26(n19218), .P25(n19217), .P24(n19216), .P23(n19215), 
            .P22(n19214), .P21(n19213), .P20(n19212), .P19(n19211), 
            .P18(n19210), .P17(n19209), .P16(n19208), .P15(n19207), 
            .P14(n19206), .P13(n19205), .P12(n19204), .P11(n19203), 
            .P10(n19202), .P9(n19201), .P8(n19200), .P7(n19199), .P6(n19198), 
            .P5(n19197), .P4(n19196), .P3(n19195), .P2(n19194), .P1(n19193), 
            .P0(n19192), .SIGNEDP(n19191));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[19:38])
    defparam mult_4003_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_4003_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_4003_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_4003_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_4003_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_4003_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_4003_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_4003_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_4003_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_4003_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_4003_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_4003_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_4003_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_4003_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_4003_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_4003_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_4003_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_4003_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_4003_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_4003_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_4003_mult_2.GSR = "ENABLED";
    defparam mult_4003_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_4003_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_4003_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_4003_mult_2.RESETMODE = "SYNC";
    ALU54B lat_alu_9 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18976), .SIGNEDIB(n19049), .SIGNEDCIN(n19122), .A35(n18975), 
           .A34(n18974), .A33(n18973), .A32(n18972), .A31(n18971), .A30(n18970), 
           .A29(n18969), .A28(n18968), .A27(n18967), .A26(n18966), .A25(n18965), 
           .A24(n18964), .A23(n18963), .A22(n18962), .A21(n18961), .A20(n18960), 
           .A19(n18959), .A18(n18958), .A17(n18957), .A16(n18956), .A15(n18955), 
           .A14(n18954), .A13(n18953), .A12(n18952), .A11(n18951), .A10(n18950), 
           .A9(n18949), .A8(n18948), .A7(n18947), .A6(n18946), .A5(n18945), 
           .A4(n18944), .A3(n18943), .A2(n18942), .A1(n18941), .A0(n18940), 
           .B35(n19048), .B34(n19047), .B33(n19046), .B32(n19045), .B31(n19044), 
           .B30(n19043), .B29(n19042), .B28(n19041), .B27(n19040), .B26(n19039), 
           .B25(n19038), .B24(n19037), .B23(n19036), .B22(n19035), .B21(n19034), 
           .B20(n19033), .B19(n19032), .B18(n19031), .B17(n19030), .B16(n19029), 
           .B15(n19028), .B14(n19027), .B13(n19026), .B12(n19025), .B11(n19024), 
           .B10(n19023), .B9(n19022), .B8(n19021), .B7(n19020), .B6(n19019), 
           .B5(n19018), .B4(n19017), .B3(n19016), .B2(n19015), .B1(n19014), 
           .B0(n19013), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n19012), .MA34(n19011), .MA33(n19010), .MA32(n19009), 
           .MA31(n19008), .MA30(n19007), .MA29(n19006), .MA28(n19005), 
           .MA27(n19004), .MA26(n19003), .MA25(n19002), .MA24(n19001), 
           .MA23(n19000), .MA22(n18999), .MA21(n18998), .MA20(n18997), 
           .MA19(n18996), .MA18(n18995), .MA17(n18994), .MA16(n18993), 
           .MA15(n18992), .MA14(n18991), .MA13(n18990), .MA12(n18989), 
           .MA11(n18988), .MA10(n18987), .MA9(n18986), .MA8(n18985), 
           .MA7(n18984), .MA6(n18983), .MA5(n18982), .MA4(n18981), .MA3(n18980), 
           .MA2(n18979), .MA1(n18978), .MA0(n18977), .MB35(n19085), 
           .MB34(n19084), .MB33(n19083), .MB32(n19082), .MB31(n19081), 
           .MB30(n19080), .MB29(n19079), .MB28(n19078), .MB27(n19077), 
           .MB26(n19076), .MB25(n19075), .MB24(n19074), .MB23(n19073), 
           .MB22(n19072), .MB21(n19071), .MB20(n19070), .MB19(n19069), 
           .MB18(n19068), .MB17(n19067), .MB16(n19066), .MB15(n19065), 
           .MB14(n19064), .MB13(n19063), .MB12(n19062), .MB11(n19061), 
           .MB10(n19060), .MB9(n19059), .MB8(n19058), .MB7(n19057), 
           .MB6(n19056), .MB5(n19055), .MB4(n19054), .MB3(n19053), .MB2(n19052), 
           .MB1(n19051), .MB0(n19050), .CIN53(n19121), .CIN52(n19120), 
           .CIN51(n19119), .CIN50(n19118), .CIN49(n19117), .CIN48(n19116), 
           .CIN47(n19115), .CIN46(n19114), .CIN45(n19113), .CIN44(n19112), 
           .CIN43(n19111), .CIN42(n19110), .CIN41(n19109), .CIN40(n19108), 
           .CIN39(n19107), .CIN38(n19106), .CIN37(n19105), .CIN36(n19104), 
           .CIN35(n19103), .CIN34(n19102), .CIN33(n19101), .CIN32(n19100), 
           .CIN31(n19099), .CIN30(n19098), .CIN29(n19097), .CIN28(n19096), 
           .CIN27(n19095), .CIN26(n19094), .CIN25(n19093), .CIN24(n19092), 
           .CIN23(n19091), .CIN22(n19090), .CIN21(n19089), .CIN20(n19088), 
           .CIN19(n19087), .CIN18(n19086), .CIN17(n177), .CIN16(n178_adj_5), 
           .CIN15(n179), .CIN14(n180), .CIN13(n181), .CIN12(n182), .CIN11(n183_adj_3), 
           .CIN10(n184), .CIN9(n185), .CIN8(n186), .CIN7(n187), .CIN6(n188_adj_2), 
           .CIN5(n189), .CIN4(n190), .CIN3(n191), .CIN2(n192), .CIN1(n193_adj_1), 
           .CIN0(n194), .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), 
           .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), 
           .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), 
           .R13(n163_adj_12), .R12(n164), .R11(n165), .R10(n166), .R9(n167), 
           .R8(n168_adj_10), .R7(n169), .R6(n170), .R5(n171), .R4(n172_adj_8), 
           .R3(n173_adj_9), .R2(n174), .R1(n175), .R0(n176));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(102[16:35])
    defparam lat_alu_9.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_9.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_9.REG_FLAG_CLK = "NONE";
    defparam lat_alu_9.REG_FLAG_CE = "CE0";
    defparam lat_alu_9.REG_FLAG_RST = "RST0";
    defparam lat_alu_9.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASK01 = "0x00000000000000";
    defparam lat_alu_9.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_9.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_9.CLK0_DIV = "ENABLED";
    defparam lat_alu_9.CLK1_DIV = "ENABLED";
    defparam lat_alu_9.CLK2_DIV = "ENABLED";
    defparam lat_alu_9.CLK3_DIV = "ENABLED";
    defparam lat_alu_9.MCPAT = "0x00000000000000";
    defparam lat_alu_9.MASKPAT = "0x00000000000000";
    defparam lat_alu_9.RNDPAT = "0x00000000000000";
    defparam lat_alu_9.GSR = "ENABLED";
    defparam lat_alu_9.RESETMODE = "SYNC";
    defparam lat_alu_9.MULT9_MODE = "DISABLED";
    defparam lat_alu_9.LEGACY = "DISABLED";
    ALU54B lat_alu_8 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18830), .SIGNEDIB(n18903), .SIGNEDCIN(GND_net), 
           .A35(n18829), .A34(n18828), .A33(n18827), .A32(n18826), .A31(n18825), 
           .A30(n18824), .A29(n18823), .A28(n18822), .A27(n18821), .A26(n18820), 
           .A25(n18819), .A24(n18818), .A23(n18817), .A22(n18816), .A21(n18815), 
           .A20(n18814), .A19(n18813), .A18(n18812), .A17(n18811), .A16(n18810), 
           .A15(n18809), .A14(n18808), .A13(n18807), .A12(n18806), .A11(n18805), 
           .A10(n18804), .A9(n18803), .A8(n18802), .A7(n18801), .A6(n18800), 
           .A5(n18799), .A4(n18798), .A3(n18797), .A2(n18796), .A1(n18795), 
           .A0(n18794), .B35(n18902), .B34(n18901), .B33(n18900), .B32(n18899), 
           .B31(n18898), .B30(n18897), .B29(n18896), .B28(n18895), .B27(n18894), 
           .B26(n18893), .B25(n18892), .B24(n18891), .B23(n18890), .B22(n18889), 
           .B21(n18888), .B20(n18887), .B19(n18886), .B18(n18885), .B17(n18884), 
           .B16(n18883), .B15(n18882), .B14(n18881), .B13(n18880), .B12(n18879), 
           .B11(n18878), .B10(n18877), .B9(n18876), .B8(n18875), .B7(n18874), 
           .B6(n18873), .B5(n18872), .B4(n18871), .B3(n18870), .B2(n18869), 
           .B1(n18868), .B0(n18867), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18866), .MA34(n18865), .MA33(n18864), .MA32(n18863), 
           .MA31(n18862), .MA30(n18861), .MA29(n18860), .MA28(n18859), 
           .MA27(n18858), .MA26(n18857), .MA25(n18856), .MA24(n18855), 
           .MA23(n18854), .MA22(n18853), .MA21(n18852), .MA20(n18851), 
           .MA19(n18850), .MA18(n18849), .MA17(n18848), .MA16(n18847), 
           .MA15(n18846), .MA14(n18845), .MA13(n18844), .MA12(n18843), 
           .MA11(n18842), .MA10(n18841), .MA9(n18840), .MA8(n18839), 
           .MA7(n18838), .MA6(n18837), .MA5(n18836), .MA4(n18835), .MA3(n18834), 
           .MA2(n18833), .MA1(n18832), .MA0(n18831), .MB35(n18939), 
           .MB34(n18938), .MB33(n18937), .MB32(n18936), .MB31(n18935), 
           .MB30(n18934), .MB29(n18933), .MB28(n18932), .MB27(n18931), 
           .MB26(n18930), .MB25(n18929), .MB24(n18928), .MB23(n18927), 
           .MB22(n18926), .MB21(n18925), .MB20(n18924), .MB19(n18923), 
           .MB18(n18922), .MB17(n18921), .MB16(n18920), .MB15(n18919), 
           .MB14(n18918), .MB13(n18917), .MB12(n18916), .MB11(n18915), 
           .MB10(n18914), .MB9(n18913), .MB8(n18912), .MB7(n18911), 
           .MB6(n18910), .MB5(n18909), .MB4(n18908), .MB3(n18907), .MB2(n18906), 
           .MB1(n18905), .MB0(n18904), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n19121), 
           .R52(n19120), .R51(n19119), .R50(n19118), .R49(n19117), .R48(n19116), 
           .R47(n19115), .R46(n19114), .R45(n19113), .R44(n19112), .R43(n19111), 
           .R42(n19110), .R41(n19109), .R40(n19108), .R39(n19107), .R38(n19106), 
           .R37(n19105), .R36(n19104), .R35(n19103), .R34(n19102), .R33(n19101), 
           .R32(n19100), .R31(n19099), .R30(n19098), .R29(n19097), .R28(n19096), 
           .R27(n19095), .R26(n19094), .R25(n19093), .R24(n19092), .R23(n19091), 
           .R22(n19090), .R21(n19089), .R20(n19088), .R19(n19087), .R18(n19086), 
           .R17(n177), .R16(n178_adj_5), .R15(n179), .R14(n180), .R13(n181), 
           .R12(n182), .R11(n183_adj_3), .R10(n184), .R9(n185), .R8(n186), 
           .R7(n187), .R6(n188_adj_2), .R5(n189), .R4(n190), .R3(n191), 
           .R2(n192), .R1(n193_adj_1), .R0(n194), .SIGNEDR(n19122));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(102[16:35])
    defparam lat_alu_8.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_8.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_8.REG_FLAG_CLK = "NONE";
    defparam lat_alu_8.REG_FLAG_CE = "CE0";
    defparam lat_alu_8.REG_FLAG_RST = "RST0";
    defparam lat_alu_8.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASK01 = "0x00000000000000";
    defparam lat_alu_8.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_8.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_8.CLK0_DIV = "ENABLED";
    defparam lat_alu_8.CLK1_DIV = "ENABLED";
    defparam lat_alu_8.CLK2_DIV = "ENABLED";
    defparam lat_alu_8.CLK3_DIV = "ENABLED";
    defparam lat_alu_8.MCPAT = "0x00000000000000";
    defparam lat_alu_8.MASKPAT = "0x00000000000000";
    defparam lat_alu_8.RNDPAT = "0x00000000000000";
    defparam lat_alu_8.GSR = "ENABLED";
    defparam lat_alu_8.RESETMODE = "SYNC";
    defparam lat_alu_8.MULT9_MODE = "DISABLED";
    defparam lat_alu_8.LEGACY = "DISABLED";
    OB x_out_pad_123 (.I(x_out_c_123), .O(x_out[123]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    MULT18X18D lat_mult_7 (.A17(\U[3] [31]), .A16(\U[3] [31]), .A15(\U[3] [31]), 
            .A14(\U[3] [31]), .A13(\U[3] [31]), .A12(\U[3] [30]), .A11(\U[3] [29]), 
            .A10(\U[3] [28]), .A9(\U[3] [27]), .A8(\U[3] [26]), .A7(\U[3] [25]), 
            .A6(\U[3] [24]), .A5(\U[3] [23]), .A4(\U[3] [22]), .A3(\U[3] [21]), 
            .A2(\U[3] [20]), .A1(\U[3] [19]), .A0(\U[3] [18]), .B17(\x[3] [31]), 
            .B16(\x[3] [31]), .B15(\x[3] [31]), .B14(\x[3] [31]), .B13(\x[3] [31]), 
            .B12(\x[3] [30]), .B11(\x[3] [29]), .B10(\x[3] [28]), .B9(\x[3] [27]), 
            .B8(\x[3] [26]), .B7(\x[3] [25]), .B6(\x[3] [24]), .B5(\x[3] [23]), 
            .B4(\x[3] [22]), .B3(\x[3] [21]), .B2(\x[3] [20]), .B1(\x[3] [19]), 
            .B0(\x[3] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19030), 
            .ROA16(n19029), .ROA15(n19028), .ROA14(n19027), .ROA13(n19026), 
            .ROA12(n19025), .ROA11(n19024), .ROA10(n19023), .ROA9(n19022), 
            .ROA8(n19021), .ROA7(n19020), .ROA6(n19019), .ROA5(n19018), 
            .ROA4(n19017), .ROA3(n19016), .ROA2(n19015), .ROA1(n19014), 
            .ROA0(n19013), .ROB17(n19048), .ROB16(n19047), .ROB15(n19046), 
            .ROB14(n19045), .ROB13(n19044), .ROB12(n19043), .ROB11(n19042), 
            .ROB10(n19041), .ROB9(n19040), .ROB8(n19039), .ROB7(n19038), 
            .ROB6(n19037), .ROB5(n19036), .ROB4(n19035), .ROB3(n19034), 
            .ROB2(n19033), .ROB1(n19032), .ROB0(n19031), .P35(n19085), 
            .P34(n19084), .P33(n19083), .P32(n19082), .P31(n19081), 
            .P30(n19080), .P29(n19079), .P28(n19078), .P27(n19077), 
            .P26(n19076), .P25(n19075), .P24(n19074), .P23(n19073), 
            .P22(n19072), .P21(n19071), .P20(n19070), .P19(n19069), 
            .P18(n19068), .P17(n19067), .P16(n19066), .P15(n19065), 
            .P14(n19064), .P13(n19063), .P12(n19062), .P11(n19061), 
            .P10(n19060), .P9(n19059), .P8(n19058), .P7(n19057), .P6(n19056), 
            .P5(n19055), .P4(n19054), .P3(n19053), .P2(n19052), .P1(n19051), 
            .P0(n19050), .SIGNEDP(n19049));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(102[16:35])
    defparam lat_mult_7.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTA_CE = "CE0";
    defparam lat_mult_7.REG_INPUTA_RST = "RST0";
    defparam lat_mult_7.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTB_CE = "CE0";
    defparam lat_mult_7.REG_INPUTB_RST = "RST0";
    defparam lat_mult_7.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTC_CE = "CE0";
    defparam lat_mult_7.REG_INPUTC_RST = "RST0";
    defparam lat_mult_7.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_7.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_7.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_7.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_7.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_7.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_7.CLK0_DIV = "ENABLED";
    defparam lat_mult_7.CLK1_DIV = "ENABLED";
    defparam lat_mult_7.CLK2_DIV = "ENABLED";
    defparam lat_mult_7.CLK3_DIV = "ENABLED";
    defparam lat_mult_7.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_7.GSR = "ENABLED";
    defparam lat_mult_7.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_7.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_7.MULT_BYPASS = "DISABLED";
    defparam lat_mult_7.RESETMODE = "SYNC";
    LUT4 i25717_4_lut_4_lut (.A(n42466), .B(n39520), .C(n54_adj_698), 
         .D(n10_adj_672), .Z(n56_adj_699)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25717_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i24873_3_lut (.A(\U[8] [1]), .B(\U[9] [1]), .C(i[0]), .Z(n40133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24873_3_lut.init = 16'hcaca;
    LUT4 i23302_4_lut (.A(n42591), .B(n42593), .C(n42592), .D(n38546), 
         .Z(n38562)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23302_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_1337_i59_2_lut_rep_1048 (.A(n2083), .B(n124_adj_229), 
         .Z(n42747)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i59_2_lut_rep_1048.init = 16'h6666;
    FD1P3AX x_out_i0_i1 (.D(\x[0] [0]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_0));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i1.GSR = "ENABLED";
    FD1P3IX state_FSM_i1 (.D(n37411), .SP(done_N_1932), .CD(rst_c), .CK(clk_c), 
            .Q(done_N_1934));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 i25910_4_lut (.A(n42439), .B(n49_adj_782), .C(n47_adj_780), .D(n40011), 
         .Z(n40027)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25910_4_lut.init = 16'hfffe;
    MULT18X18D lat_mult_6 (.A17(\U[3] [17]), .A16(\U[3] [16]), .A15(\U[3] [15]), 
            .A14(\U[3] [14]), .A13(\U[3] [13]), .A12(\U[3] [12]), .A11(\U[3] [11]), 
            .A10(\U[3] [10]), .A9(\U[3] [9]), .A8(\U[3] [8]), .A7(\U[3] [7]), 
            .A6(\U[3] [6]), .A5(\U[3] [5]), .A4(\U[3] [4]), .A3(\U[3] [3]), 
            .A2(\U[3] [2]), .A1(\U[3] [1]), .A0(\U[3] [0]), .B17(\x[3] [31]), 
            .B16(\x[3] [31]), .B15(\x[3] [31]), .B14(\x[3] [31]), .B13(\x[3] [31]), 
            .B12(\x[3] [30]), .B11(\x[3] [29]), .B10(\x[3] [28]), .B9(\x[3] [27]), 
            .B8(\x[3] [26]), .B7(\x[3] [25]), .B6(\x[3] [24]), .B5(\x[3] [23]), 
            .B4(\x[3] [22]), .B3(\x[3] [21]), .B2(\x[3] [20]), .B1(\x[3] [19]), 
            .B0(\x[3] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18957), 
            .ROA16(n18956), .ROA15(n18955), .ROA14(n18954), .ROA13(n18953), 
            .ROA12(n18952), .ROA11(n18951), .ROA10(n18950), .ROA9(n18949), 
            .ROA8(n18948), .ROA7(n18947), .ROA6(n18946), .ROA5(n18945), 
            .ROA4(n18944), .ROA3(n18943), .ROA2(n18942), .ROA1(n18941), 
            .ROA0(n18940), .ROB17(n18975), .ROB16(n18974), .ROB15(n18973), 
            .ROB14(n18972), .ROB13(n18971), .ROB12(n18970), .ROB11(n18969), 
            .ROB10(n18968), .ROB9(n18967), .ROB8(n18966), .ROB7(n18965), 
            .ROB6(n18964), .ROB5(n18963), .ROB4(n18962), .ROB3(n18961), 
            .ROB2(n18960), .ROB1(n18959), .ROB0(n18958), .P35(n19012), 
            .P34(n19011), .P33(n19010), .P32(n19009), .P31(n19008), 
            .P30(n19007), .P29(n19006), .P28(n19005), .P27(n19004), 
            .P26(n19003), .P25(n19002), .P24(n19001), .P23(n19000), 
            .P22(n18999), .P21(n18998), .P20(n18997), .P19(n18996), 
            .P18(n18995), .P17(n18994), .P16(n18993), .P15(n18992), 
            .P14(n18991), .P13(n18990), .P12(n18989), .P11(n18988), 
            .P10(n18987), .P9(n18986), .P8(n18985), .P7(n18984), .P6(n18983), 
            .P5(n18982), .P4(n18981), .P3(n18980), .P2(n18979), .P1(n18978), 
            .P0(n18977), .SIGNEDP(n18976));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(102[16:35])
    defparam lat_mult_6.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTA_CE = "CE0";
    defparam lat_mult_6.REG_INPUTA_RST = "RST0";
    defparam lat_mult_6.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTB_CE = "CE0";
    defparam lat_mult_6.REG_INPUTB_RST = "RST0";
    defparam lat_mult_6.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTC_CE = "CE0";
    defparam lat_mult_6.REG_INPUTC_RST = "RST0";
    defparam lat_mult_6.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_6.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_6.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_6.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_6.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_6.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_6.CLK0_DIV = "ENABLED";
    defparam lat_mult_6.CLK1_DIV = "ENABLED";
    defparam lat_mult_6.CLK2_DIV = "ENABLED";
    defparam lat_mult_6.CLK3_DIV = "ENABLED";
    defparam lat_mult_6.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_6.GSR = "ENABLED";
    defparam lat_mult_6.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_6.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_6.MULT_BYPASS = "DISABLED";
    defparam lat_mult_6.RESETMODE = "SYNC";
    MULT18X18D lat_mult_12 (.A17(\U[6] [31]), .A16(\U[6] [31]), .A15(\U[6] [31]), 
            .A14(\U[6] [31]), .A13(\U[6] [31]), .A12(\U[6] [30]), .A11(\U[6] [29]), 
            .A10(\U[6] [28]), .A9(\U[6] [27]), .A8(\U[6] [26]), .A7(\U[6] [25]), 
            .A6(\U[6] [24]), .A5(\U[6] [23]), .A4(\U[6] [22]), .A3(\U[6] [21]), 
            .A2(\U[6] [20]), .A1(\U[6] [19]), .A0(\U[6] [18]), .B17(\x[2] [31]), 
            .B16(\x[2] [31]), .B15(\x[2] [31]), .B14(\x[2] [31]), .B13(\x[2] [31]), 
            .B12(\x[2] [30]), .B11(\x[2] [29]), .B10(\x[2] [28]), .B9(\x[2] [27]), 
            .B8(\x[2] [26]), .B7(\x[2] [25]), .B6(\x[2] [24]), .B5(\x[2] [23]), 
            .B4(\x[2] [22]), .B3(\x[2] [21]), .B2(\x[2] [20]), .B1(\x[2] [19]), 
            .B0(\x[2] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19391), 
            .ROA16(n19390), .ROA15(n19389), .ROA14(n19388), .ROA13(n19387), 
            .ROA12(n19386), .ROA11(n19385), .ROA10(n19384), .ROA9(n19383), 
            .ROA8(n19382), .ROA7(n19381), .ROA6(n19380), .ROA5(n19379), 
            .ROA4(n19378), .ROA3(n19377), .ROA2(n19376), .ROA1(n19375), 
            .ROA0(n19374), .ROB17(n19409), .ROB16(n19408), .ROB15(n19407), 
            .ROB14(n19406), .ROB13(n19405), .ROB12(n19404), .ROB11(n19403), 
            .ROB10(n19402), .ROB9(n19401), .ROB8(n19400), .ROB7(n19399), 
            .ROB6(n19398), .ROB5(n19397), .ROB4(n19396), .ROB3(n19395), 
            .ROB2(n19394), .ROB1(n19393), .ROB0(n19392), .P35(n19446), 
            .P34(n19445), .P33(n19444), .P32(n19443), .P31(n19442), 
            .P30(n19441), .P29(n19440), .P28(n19439), .P27(n19438), 
            .P26(n19437), .P25(n19436), .P24(n19435), .P23(n19434), 
            .P22(n19433), .P21(n19432), .P20(n19431), .P19(n19430), 
            .P18(n19429), .P17(n19428), .P16(n19427), .P15(n19426), 
            .P14(n19425), .P13(n19424), .P12(n19423), .P11(n19422), 
            .P10(n19421), .P9(n19420), .P8(n19419), .P7(n19418), .P6(n19417), 
            .P5(n19416), .P4(n19415), .P3(n19414), .P2(n19413), .P1(n19412), 
            .P0(n19411), .SIGNEDP(n19410));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[19:38])
    defparam lat_mult_12.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTA_CE = "CE0";
    defparam lat_mult_12.REG_INPUTA_RST = "RST0";
    defparam lat_mult_12.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTB_CE = "CE0";
    defparam lat_mult_12.REG_INPUTB_RST = "RST0";
    defparam lat_mult_12.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTC_CE = "CE0";
    defparam lat_mult_12.REG_INPUTC_RST = "RST0";
    defparam lat_mult_12.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_12.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_12.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_12.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_12.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_12.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_12.CLK0_DIV = "ENABLED";
    defparam lat_mult_12.CLK1_DIV = "ENABLED";
    defparam lat_mult_12.CLK2_DIV = "ENABLED";
    defparam lat_mult_12.CLK3_DIV = "ENABLED";
    defparam lat_mult_12.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_12.GSR = "ENABLED";
    defparam lat_mult_12.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_12.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_12.MULT_BYPASS = "DISABLED";
    defparam lat_mult_12.RESETMODE = "SYNC";
    MULT18X18D lat_mult_20 (.A17(\U[7] [31]), .A16(\U[7] [31]), .A15(\U[7] [31]), 
            .A14(\U[7] [31]), .A13(\U[7] [31]), .A12(\U[7] [30]), .A11(\U[7] [29]), 
            .A10(\U[7] [28]), .A9(\U[7] [27]), .A8(\U[7] [26]), .A7(\U[7] [25]), 
            .A6(\U[7] [24]), .A5(\U[7] [23]), .A4(\U[7] [22]), .A3(\U[7] [21]), 
            .A2(\U[7] [20]), .A1(\U[7] [19]), .A0(\U[7] [18]), .B17(\x[3] [17]), 
            .B16(\x[3] [16]), .B15(\x[3] [15]), .B14(\x[3] [14]), .B13(\x[3] [13]), 
            .B12(\x[3] [12]), .B11(\x[3] [11]), .B10(\x[3] [10]), .B9(\x[3] [9]), 
            .B8(\x[3] [8]), .B7(\x[3] [7]), .B6(\x[3] [6]), .B5(\x[3] [5]), 
            .B4(\x[3] [4]), .B3(\x[3] [3]), .B2(\x[3] [2]), .B1(\x[3] [1]), 
            .B0(\x[3] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19967), 
            .ROA16(n19966), .ROA15(n19965), .ROA14(n19964), .ROA13(n19963), 
            .ROA12(n19962), .ROA11(n19961), .ROA10(n19960), .ROA9(n19959), 
            .ROA8(n19958), .ROA7(n19957), .ROA6(n19956), .ROA5(n19955), 
            .ROA4(n19954), .ROA3(n19953), .ROA2(n19952), .ROA1(n19951), 
            .ROA0(n19950), .ROB17(n19985), .ROB16(n19984), .ROB15(n19983), 
            .ROB14(n19982), .ROB13(n19981), .ROB12(n19980), .ROB11(n19979), 
            .ROB10(n19978), .ROB9(n19977), .ROB8(n19976), .ROB7(n19975), 
            .ROB6(n19974), .ROB5(n19973), .ROB4(n19972), .ROB3(n19971), 
            .ROB2(n19970), .ROB1(n19969), .ROB0(n19968), .P35(n20022), 
            .P34(n20021), .P33(n20020), .P32(n20019), .P31(n20018), 
            .P30(n20017), .P29(n20016), .P28(n20015), .P27(n20014), 
            .P26(n20013), .P25(n20012), .P24(n20011), .P23(n20010), 
            .P22(n20009), .P21(n20008), .P20(n20007), .P19(n20006), 
            .P18(n20005), .P17(n20004), .P16(n20003), .P15(n20002), 
            .P14(n20001), .P13(n20000), .P12(n19999), .P11(n19998), 
            .P10(n19997), .P9(n19996), .P8(n19995), .P7(n19994), .P6(n19993), 
            .P5(n19992), .P4(n19991), .P3(n19990), .P2(n19989), .P1(n19988), 
            .P0(n19987), .SIGNEDP(n19986));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(106[16:35])
    defparam lat_mult_20.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_20.REG_INPUTA_CE = "CE0";
    defparam lat_mult_20.REG_INPUTA_RST = "RST0";
    defparam lat_mult_20.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_20.REG_INPUTB_CE = "CE0";
    defparam lat_mult_20.REG_INPUTB_RST = "RST0";
    defparam lat_mult_20.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_20.REG_INPUTC_CE = "CE0";
    defparam lat_mult_20.REG_INPUTC_RST = "RST0";
    defparam lat_mult_20.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_20.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_20.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_20.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_20.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_20.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_20.CLK0_DIV = "ENABLED";
    defparam lat_mult_20.CLK1_DIV = "ENABLED";
    defparam lat_mult_20.CLK2_DIV = "ENABLED";
    defparam lat_mult_20.CLK3_DIV = "ENABLED";
    defparam lat_mult_20.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_20.GSR = "ENABLED";
    defparam lat_mult_20.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_20.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_20.MULT_BYPASS = "DISABLED";
    defparam lat_mult_20.RESETMODE = "SYNC";
    FD1S3JX state_FSM_i4 (.D(n27528), .CK(clk_c), .PD(rst_c), .Q(done_N_1929));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam state_FSM_i4.GSR = "ENABLED";
    MULT18X18D lat_mult_21 (.A17(\U[7] [17]), .A16(\U[7] [16]), .A15(\U[7] [15]), 
            .A14(\U[7] [14]), .A13(\U[7] [13]), .A12(\U[7] [12]), .A11(\U[7] [11]), 
            .A10(\U[7] [10]), .A9(\U[7] [9]), .A8(\U[7] [8]), .A7(\U[7] [7]), 
            .A6(\U[7] [6]), .A5(\U[7] [5]), .A4(\U[7] [4]), .A3(\U[7] [3]), 
            .A2(\U[7] [2]), .A1(\U[7] [1]), .A0(\U[7] [0]), .B17(\x[3] [31]), 
            .B16(\x[3] [31]), .B15(\x[3] [31]), .B14(\x[3] [31]), .B13(\x[3] [31]), 
            .B12(\x[3] [30]), .B11(\x[3] [29]), .B10(\x[3] [28]), .B9(\x[3] [27]), 
            .B8(\x[3] [26]), .B7(\x[3] [25]), .B6(\x[3] [24]), .B5(\x[3] [23]), 
            .B4(\x[3] [22]), .B3(\x[3] [21]), .B2(\x[3] [20]), .B1(\x[3] [19]), 
            .B0(\x[3] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n20040), 
            .ROA16(n20039), .ROA15(n20038), .ROA14(n20037), .ROA13(n20036), 
            .ROA12(n20035), .ROA11(n20034), .ROA10(n20033), .ROA9(n20032), 
            .ROA8(n20031), .ROA7(n20030), .ROA6(n20029), .ROA5(n20028), 
            .ROA4(n20027), .ROA3(n20026), .ROA2(n20025), .ROA1(n20024), 
            .ROA0(n20023), .ROB17(n20058), .ROB16(n20057), .ROB15(n20056), 
            .ROB14(n20055), .ROB13(n20054), .ROB12(n20053), .ROB11(n20052), 
            .ROB10(n20051), .ROB9(n20050), .ROB8(n20049), .ROB7(n20048), 
            .ROB6(n20047), .ROB5(n20046), .ROB4(n20045), .ROB3(n20044), 
            .ROB2(n20043), .ROB1(n20042), .ROB0(n20041), .P35(n20095), 
            .P34(n20094), .P33(n20093), .P32(n20092), .P31(n20091), 
            .P30(n20090), .P29(n20089), .P28(n20088), .P27(n20087), 
            .P26(n20086), .P25(n20085), .P24(n20084), .P23(n20083), 
            .P22(n20082), .P21(n20081), .P20(n20080), .P19(n20079), 
            .P18(n20078), .P17(n20077), .P16(n20076), .P15(n20075), 
            .P14(n20074), .P13(n20073), .P12(n20072), .P11(n20071), 
            .P10(n20070), .P9(n20069), .P8(n20068), .P7(n20067), .P6(n20066), 
            .P5(n20065), .P4(n20064), .P3(n20063), .P2(n20062), .P1(n20061), 
            .P0(n20060), .SIGNEDP(n20059));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(106[16:35])
    defparam lat_mult_21.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_21.REG_INPUTA_CE = "CE0";
    defparam lat_mult_21.REG_INPUTA_RST = "RST0";
    defparam lat_mult_21.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_21.REG_INPUTB_CE = "CE0";
    defparam lat_mult_21.REG_INPUTB_RST = "RST0";
    defparam lat_mult_21.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_21.REG_INPUTC_CE = "CE0";
    defparam lat_mult_21.REG_INPUTC_RST = "RST0";
    defparam lat_mult_21.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_21.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_21.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_21.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_21.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_21.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_21.CLK0_DIV = "ENABLED";
    defparam lat_mult_21.CLK1_DIV = "ENABLED";
    defparam lat_mult_21.CLK2_DIV = "ENABLED";
    defparam lat_mult_21.CLK3_DIV = "ENABLED";
    defparam lat_mult_21.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_21.GSR = "ENABLED";
    defparam lat_mult_21.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_21.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_21.MULT_BYPASS = "DISABLED";
    defparam lat_mult_21.RESETMODE = "SYNC";
    PFUMX div_4016_LessThan_2841_i62 (.BLUT(n58_adj_605), .ALUT(n60_adj_606), 
          .C0(n39028), .Z(n62_adj_607));
    LUT4 div_4016_LessThan_2681_i57_2_lut_rep_871 (.A(n4079), .B(n111), 
         .Z(n42570)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i57_2_lut_rep_871.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i54_3_lut_3_lut (.A(n4197), .B(n108), .C(n109_adj_219), 
         .Z(n54_adj_573)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23286_4_lut (.A(n42594), .B(n43_adj_509), .C(n31_adj_501), .D(n38499), 
         .Z(n38546)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23286_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_1337_i50_3_lut_3_lut (.A(n2083), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n50_adj_271)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24751_3_lut (.A(n45_adj_778), .B(n43_adj_776), .C(n19_adj_753), 
         .Z(n40011)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24751_3_lut.init = 16'h0101;
    LUT4 i25794_4_lut_4_lut (.A(n42466), .B(n39511), .C(n42465), .D(n42464), 
         .Z(n39531)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25794_4_lut_4_lut.init = 16'hff04;
    LUT4 div_4016_LessThan_1337_i55_2_lut_rep_1049 (.A(n2085), .B(n126), 
         .Z(n42748)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i55_2_lut_rep_1049.init = 16'h6666;
    LUT4 div_4016_i489_3_lut_4_lut (.A(n42776), .B(n30965), .C(n132), 
         .D(n42784), .Z(n865)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam div_4016_i489_3_lut_4_lut.init = 16'hef10;
    LUT4 div_4016_LessThan_3206_i39_4_lut (.A(n4763), .B(n113_adj_222), 
         .C(n22253), .D(n4783), .Z(n39_adj_773)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i39_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_3206_i19_4_lut (.A(n4773), .B(n123), .C(n22263), 
         .D(n4783), .Z(n19_adj_753)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i19_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2681_i30_3_lut_3_lut (.A(n4079), .B(n111), .C(n123), 
         .Z(n30_adj_530)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i3313_3_lut_4_lut (.A(n42776), .B(n30965), .C(n42786), 
         .D(n22277), .Z(n5496)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam div_4016_i3313_3_lut_4_lut.init = 16'hf101;
    LUT4 div_4016_LessThan_2598_i43_2_lut (.A(n3963), .B(n119_adj_226), 
         .Z(n43_adj_509)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i43_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2681_i53_2_lut_rep_872 (.A(n4081), .B(n113_adj_222), 
         .Z(n42571)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i53_2_lut_rep_872.init = 16'h6666;
    LUT4 i25775_4_lut (.A(n42445), .B(n42448), .C(n42447), .D(n39660), 
         .Z(n39678)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25775_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2598_i31_2_lut (.A(n3969), .B(n125_adj_230), 
         .Z(n31_adj_501)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i31_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_1076_4_lut_4_lut (.A(n35964), .B(n130_adj_233), .C(n30965), 
         .D(n62_adj_798), .Z(n42775)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (C+(D))+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i1_2_lut_rep_1076_4_lut_4_lut.init = 16'hfef8;
    LUT4 div_4016_LessThan_1337_i52_3_lut_3_lut (.A(n2085), .B(n126), .C(n127_adj_231), 
         .Z(n52_adj_272)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3137_i13_2_lut_rep_763 (.A(n4776), .B(n127_adj_231), 
         .Z(n42462)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i13_2_lut_rep_763.init = 16'h6666;
    L6MUX21 div_4016_LessThan_2841_i50 (.D0(n38_adj_595), .D1(n48_adj_600), 
            .SD(n38980), .Z(n50_adj_601));
    LUT4 i24254_4_lut_4_lut (.A(n42466), .B(n39487), .C(n42468), .D(n42465), 
         .Z(n39514)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24254_4_lut_4_lut.init = 16'h0004;
    LUT4 div_4016_LessThan_3206_i37_4_lut (.A(n4764), .B(n114), .C(n22254), 
         .D(n4783), .Z(n37_adj_771)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i37_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_393_i64_3_lut_rep_1077_3_lut (.A(n35964), .B(n130_adj_233), 
         .C(n62_adj_798), .Z(n42776)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_393_i64_3_lut_rep_1077_3_lut.init = 16'he8e8;
    LUT4 div_4016_LessThan_2681_i46_3_lut_3_lut (.A(n4081), .B(n113_adj_222), 
         .C(n114), .Z(n46_adj_540)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i14088_3_lut (.A(U_in_c_159), .B(\U[4] [31]), .C(done_N_1931), 
         .Z(U_0__31__N_967[383])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14088_3_lut.init = 16'hacac;
    LUT4 div_4016_LessThan_2762_i55_2_lut_rep_854 (.A(n4200), .B(n111), 
         .Z(n42553)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i55_2_lut_rep_854.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i63_2_lut_rep_765 (.A(n4646), .B(n103_adj_215), 
         .Z(n42464)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i63_2_lut_rep_765.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i58_3_lut_3_lut (.A(n4646), .B(n103_adj_215), 
         .C(n24_adj_681), .Z(n58_adj_700)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24872_3_lut (.A(\U[6] [1]), .B(\U[7] [1]), .C(i[0]), .Z(n40132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24872_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i55_2_lut_rep_873 (.A(n4080), .B(n112_adj_221), 
         .Z(n42572)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i55_2_lut_rep_873.init = 16'h6666;
    LUT4 div_4016_LessThan_1337_i49_2_lut_rep_1050 (.A(n2088), .B(n129), 
         .Z(n42749)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i49_2_lut_rep_1050.init = 16'h6666;
    LUT4 div_4016_i487_4_lut_4_lut (.A(n35964), .B(n130_adj_233), .C(n62_adj_801), 
         .D(n42775), .Z(n35968)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i487_4_lut_4_lut.init = 16'haa69;
    PFUMX div_4016_LessThan_2841_i48 (.BLUT(n40_adj_596), .ALUT(n46_adj_599), 
          .C0(n38982), .Z(n48_adj_600));
    LUT4 i14090_3_lut (.A(U_in_c_158), .B(\U[4] [30]), .C(done_N_1931), 
         .Z(U_0__31__N_967[382])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14090_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_1078 (.A(n64_adj_799), .B(n35916), .Z(n42777)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1078.init = 16'heeee;
    LUT4 i14092_3_lut (.A(U_in_c_157), .B(\U[4] [29]), .C(done_N_1931), 
         .Z(U_0__31__N_967[381])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14092_3_lut.init = 16'hacac;
    LUT4 i25714_4_lut_4_lut (.A(n42467), .B(n39493), .C(n48_adj_695), 
         .D(n12_adj_673), .Z(n50_adj_696)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25714_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2681_i48_3_lut_3_lut (.A(n4080), .B(n112_adj_221), 
         .C(n46_adj_540), .Z(n48_adj_541)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i14094_3_lut (.A(U_in_c_156), .B(\U[4] [28]), .C(done_N_1931), 
         .Z(U_0__31__N_967[380])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14094_3_lut.init = 16'hacac;
    LUT4 div_4016_i363_3_lut_4_lut (.A(n64_adj_799), .B(n35916), .C(n132), 
         .D(n42785), .Z(n678)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam div_4016_i363_3_lut_4_lut.init = 16'hef10;
    LUT4 i24227_4_lut_4_lut (.A(n42467), .B(n39466), .C(n42470), .D(n42469), 
         .Z(n39487)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24227_4_lut_4_lut.init = 16'h0004;
    LUT4 i24871_3_lut (.A(\U[4] [1]), .B(\U[5] [1]), .C(i[0]), .Z(n40131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24871_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i51_2_lut_rep_874 (.A(n4082), .B(n114), 
         .Z(n42573)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i51_2_lut_rep_874.init = 16'h6666;
    LUT4 i23444_2_lut_3_lut_4_lut (.A(n4082), .B(n114), .C(n113_adj_222), 
         .D(n4081), .Z(n38704)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23444_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_i3312_3_lut_4_lut (.A(n64_adj_799), .B(n35916), .C(n42786), 
         .D(n22276), .Z(n5495)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam div_4016_i3312_3_lut_4_lut.init = 16'hf101;
    LUT4 i24870_3_lut (.A(\U[2] [1]), .B(\U[3] [1]), .C(i[0]), .Z(n40130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24870_3_lut.init = 16'hcaca;
    LUT4 i24869_3_lut (.A(\U[0] [1]), .B(\U[1] [1]), .C(i[0]), .Z(n40129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24869_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i49_2_lut_rep_875 (.A(n4083), .B(n115_adj_223), 
         .Z(n42574)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i49_2_lut_rep_875.init = 16'h6666;
    LUT4 i14096_3_lut (.A(U_in_c_155), .B(\U[4] [27]), .C(done_N_1931), 
         .Z(U_0__31__N_967[379])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14096_3_lut.init = 16'hacac;
    LUT4 div_4016_i3322_4_lut (.A(n37186), .B(n22286), .C(n42786), .D(n64_adj_289), 
         .Z(n5505)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3322_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_2681_i41_2_lut (.A(n4087), .B(n119_adj_226), 
         .Z(n41_adj_537)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i41_2_lut.init = 16'h6666;
    FD1S3IX state_FSM_i3 (.D(n10098), .CK(clk_c), .CD(rst_c), .Q(done_N_1931));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i2 (.D(n27533), .CK(clk_c), .CD(rst_c), .Q(done_N_1932));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1P3AX x_out_i0_i128 (.D(\x[3] [31]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_127));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i128.GSR = "ENABLED";
    LUT4 i10575_2_lut_rep_1081 (.A(n2), .B(n5325), .Z(n42780)) /* synthesis lut_function=(A (B)) */ ;
    defparam i10575_2_lut_rep_1081.init = 16'h8888;
    LUT4 div_4016_LessThan_2681_i44_3_lut_3_lut (.A(n4083), .B(n115_adj_223), 
         .C(n26_adj_527), .Z(n44_adj_539)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3066_i59_2_lut_rep_766 (.A(n4648), .B(n105), 
         .Z(n42465)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i59_2_lut_rep_766.init = 16'h6666;
    LUT4 i23433_3_lut_4_lut (.A(n4083), .B(n115_adj_223), .C(n29_adj_529), 
         .D(n42576), .Z(n38693)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23433_3_lut_4_lut.init = 16'h0009;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n2), .B(n5325), .C(n131_adj_234), .D(n132), 
         .Z(n4_adj_235)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf7f0;
    LUT4 i14098_3_lut (.A(U_in_c_154), .B(\U[4] [26]), .C(done_N_1931), 
         .Z(U_0__31__N_967[378])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14098_3_lut.init = 16'hacac;
    FD1P3AX x_out_i0_i127 (.D(\x[3] [30]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_126));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i127.GSR = "ENABLED";
    FD1P3AX x_out_i0_i126 (.D(\x[3] [29]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_125));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i126.GSR = "ENABLED";
    FD1P3AX x_out_i0_i125 (.D(\x[3] [28]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_124));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i125.GSR = "ENABLED";
    FD1P3AX x_out_i0_i124 (.D(\x[3] [27]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_123));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i124.GSR = "ENABLED";
    FD1P3AX x_out_i0_i123 (.D(\x[3] [26]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_122));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i123.GSR = "ENABLED";
    FD1P3AX x_out_i0_i122 (.D(\x[3] [25]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_121));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i122.GSR = "ENABLED";
    FD1P3AX x_out_i0_i121 (.D(\x[3] [24]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_120));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i121.GSR = "ENABLED";
    FD1P3AX x_out_i0_i120 (.D(\x[3] [23]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_119));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i120.GSR = "ENABLED";
    FD1P3AX x_out_i0_i119 (.D(\x[3] [22]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_118));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i119.GSR = "ENABLED";
    FD1P3AX x_out_i0_i118 (.D(\x[3] [21]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_117));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i118.GSR = "ENABLED";
    FD1P3AX x_out_i0_i117 (.D(\x[3] [20]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_116));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i117.GSR = "ENABLED";
    FD1P3AX x_out_i0_i116 (.D(\x[3] [19]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_115));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i116.GSR = "ENABLED";
    FD1P3AX x_out_i0_i115 (.D(\x[3] [18]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_114));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i115.GSR = "ENABLED";
    FD1P3AX x_out_i0_i114 (.D(\x[3] [17]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_113));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i114.GSR = "ENABLED";
    LUT4 i16452_2_lut_rep_1079_3_lut (.A(n2), .B(n5325), .C(n132), .Z(n42778)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i16452_2_lut_rep_1079_3_lut.init = 16'h7070;
    LUT4 i14189_3_lut (.A(U_in_c_153), .B(\U[4] [25]), .C(done_N_1931), 
         .Z(U_0__31__N_967[377])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14189_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_15 (.A(n37178), .B(n35961), .C(n37180), .D(n37176), 
         .Z(n37186)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_15.init = 16'hfffe;
    FD1P3AX x_out_i0_i113 (.D(\x[3] [16]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_112));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i113.GSR = "ENABLED";
    FD1P3AX x_out_i0_i112 (.D(\x[3] [15]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_111));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i112.GSR = "ENABLED";
    FD1P3AX x_out_i0_i111 (.D(\x[3] [14]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_110));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i111.GSR = "ENABLED";
    FD1P3AX x_out_i0_i110 (.D(\x[3] [13]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_109));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i110.GSR = "ENABLED";
    FD1P3AX x_out_i0_i109 (.D(\x[3] [12]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_108));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i109.GSR = "ENABLED";
    FD1P3AX x_out_i0_i108 (.D(\x[3] [11]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_107));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i108.GSR = "ENABLED";
    FD1P3AX x_out_i0_i107 (.D(\x[3] [10]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_106));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i107.GSR = "ENABLED";
    FD1P3AX x_out_i0_i106 (.D(\x[3] [9]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_105));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i106.GSR = "ENABLED";
    FD1P3AX x_out_i0_i105 (.D(\x[3] [8]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_104));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i105.GSR = "ENABLED";
    FD1P3AX x_out_i0_i104 (.D(\x[3] [7]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_103));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i104.GSR = "ENABLED";
    FD1P3AX x_out_i0_i103 (.D(\x[3] [6]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_102));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i103.GSR = "ENABLED";
    FD1P3AX x_out_i0_i102 (.D(\x[3] [5]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_101));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i102.GSR = "ENABLED";
    FD1P3AX x_out_i0_i101 (.D(\x[3] [4]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_100));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i101.GSR = "ENABLED";
    FD1P3AX x_out_i0_i100 (.D(\x[3] [3]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_99));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i100.GSR = "ENABLED";
    FD1P3AX x_out_i0_i99 (.D(\x[3] [2]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_98));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i99.GSR = "ENABLED";
    FD1P3AX x_out_i0_i98 (.D(\x[3] [1]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_97));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i98.GSR = "ENABLED";
    FD1P3AX x_out_i0_i97 (.D(\x[3] [0]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_96));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i97.GSR = "ENABLED";
    FD1P3AX x_out_i0_i96 (.D(\x[2] [31]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_95));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i96.GSR = "ENABLED";
    FD1P3AX x_out_i0_i95 (.D(\x[2] [30]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_94));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i95.GSR = "ENABLED";
    FD1P3AX x_out_i0_i94 (.D(\x[2] [29]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_93));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i94.GSR = "ENABLED";
    FD1P3AX x_out_i0_i93 (.D(\x[2] [28]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_92));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i93.GSR = "ENABLED";
    FD1P3AX x_out_i0_i92 (.D(\x[2] [27]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_91));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i92.GSR = "ENABLED";
    FD1P3AX x_out_i0_i91 (.D(\x[2] [26]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_90));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i91.GSR = "ENABLED";
    FD1P3AX x_out_i0_i90 (.D(\x[2] [25]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_89));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i90.GSR = "ENABLED";
    FD1P3AX x_out_i0_i89 (.D(\x[2] [24]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_88));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i89.GSR = "ENABLED";
    FD1P3AX x_out_i0_i88 (.D(\x[2] [23]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_87));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i88.GSR = "ENABLED";
    FD1P3AX x_out_i0_i87 (.D(\x[2] [22]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_86));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i87.GSR = "ENABLED";
    FD1P3AX x_out_i0_i86 (.D(\x[2] [21]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_85));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i86.GSR = "ENABLED";
    FD1P3AX x_out_i0_i85 (.D(\x[2] [20]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_84));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i85.GSR = "ENABLED";
    FD1P3AX x_out_i0_i84 (.D(\x[2] [19]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_83));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i84.GSR = "ENABLED";
    FD1P3AX x_out_i0_i83 (.D(\x[2] [18]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_82));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i83.GSR = "ENABLED";
    FD1P3AX x_out_i0_i82 (.D(\x[2] [17]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_81));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i82.GSR = "ENABLED";
    FD1P3AX x_out_i0_i81 (.D(\x[2] [16]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_80));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i81.GSR = "ENABLED";
    FD1P3AX x_out_i0_i80 (.D(\x[2] [15]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_79));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i80.GSR = "ENABLED";
    FD1P3AX x_out_i0_i79 (.D(\x[2] [14]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_78));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i79.GSR = "ENABLED";
    FD1P3AX x_out_i0_i78 (.D(\x[2] [13]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_77));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i78.GSR = "ENABLED";
    FD1P3AX x_out_i0_i77 (.D(\x[2] [12]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_76));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i77.GSR = "ENABLED";
    FD1P3AX x_out_i0_i76 (.D(\x[2] [11]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_75));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i76.GSR = "ENABLED";
    FD1P3AX x_out_i0_i75 (.D(\x[2] [10]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_74));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i75.GSR = "ENABLED";
    FD1P3AX x_out_i0_i74 (.D(\x[2] [9]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_73));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i74.GSR = "ENABLED";
    FD1P3AX x_out_i0_i73 (.D(\x[2] [8]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_72));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i73.GSR = "ENABLED";
    FD1P3AX x_out_i0_i72 (.D(\x[2] [7]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_71));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i72.GSR = "ENABLED";
    FD1P3AX x_out_i0_i71 (.D(\x[2] [6]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_70));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i71.GSR = "ENABLED";
    FD1P3AX x_out_i0_i70 (.D(\x[2] [5]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_69));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i70.GSR = "ENABLED";
    FD1P3AX x_out_i0_i69 (.D(\x[2] [4]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_68));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i69.GSR = "ENABLED";
    FD1P3AX x_out_i0_i68 (.D(\x[2] [3]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_67));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i68.GSR = "ENABLED";
    FD1P3AX x_out_i0_i67 (.D(\x[2] [2]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_66));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i67.GSR = "ENABLED";
    FD1P3AX x_out_i0_i66 (.D(\x[2] [1]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_65));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i66.GSR = "ENABLED";
    FD1P3AX x_out_i0_i65 (.D(\x[2] [0]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_64));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i65.GSR = "ENABLED";
    FD1P3AX x_out_i0_i64 (.D(\x[1] [31]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_63));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i64.GSR = "ENABLED";
    FD1P3AX x_out_i0_i63 (.D(\x[1] [30]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_62));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i63.GSR = "ENABLED";
    FD1P3AX x_out_i0_i62 (.D(\x[1] [29]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_61));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i62.GSR = "ENABLED";
    FD1P3AX x_out_i0_i61 (.D(\x[1] [28]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_60));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i61.GSR = "ENABLED";
    FD1P3AX x_out_i0_i60 (.D(\x[1] [27]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_59));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i60.GSR = "ENABLED";
    FD1P3AX x_out_i0_i59 (.D(\x[1] [26]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_58));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i59.GSR = "ENABLED";
    FD1P3AX x_out_i0_i58 (.D(\x[1] [25]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_57));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i58.GSR = "ENABLED";
    FD1P3AX x_out_i0_i57 (.D(\x[1] [24]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_56));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i57.GSR = "ENABLED";
    FD1P3AX x_out_i0_i56 (.D(\x[1] [23]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_55));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i56.GSR = "ENABLED";
    FD1P3AX x_out_i0_i55 (.D(\x[1] [22]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_54));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i55.GSR = "ENABLED";
    FD1P3AX x_out_i0_i54 (.D(\x[1] [21]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_53));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i54.GSR = "ENABLED";
    FD1P3AX x_out_i0_i53 (.D(\x[1] [20]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_52));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i53.GSR = "ENABLED";
    FD1P3AX x_out_i0_i52 (.D(\x[1] [19]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_51));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i52.GSR = "ENABLED";
    FD1P3AX x_out_i0_i51 (.D(\x[1] [18]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_50));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i51.GSR = "ENABLED";
    FD1P3AX x_out_i0_i50 (.D(\x[1] [17]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_49));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i50.GSR = "ENABLED";
    FD1P3AX x_out_i0_i49 (.D(\x[1] [16]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_48));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i49.GSR = "ENABLED";
    FD1P3AX x_out_i0_i48 (.D(\x[1] [15]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_47));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i48.GSR = "ENABLED";
    FD1P3AX x_out_i0_i47 (.D(\x[1] [14]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_46));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i47.GSR = "ENABLED";
    FD1P3AX x_out_i0_i46 (.D(\x[1] [13]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_45));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i46.GSR = "ENABLED";
    FD1P3AX x_out_i0_i45 (.D(\x[1] [12]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_44));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i45.GSR = "ENABLED";
    FD1P3AX x_out_i0_i44 (.D(\x[1] [11]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_43));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i44.GSR = "ENABLED";
    FD1P3AX x_out_i0_i43 (.D(\x[1] [10]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_42));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i43.GSR = "ENABLED";
    FD1P3AX x_out_i0_i42 (.D(\x[1] [9]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_41));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i42.GSR = "ENABLED";
    FD1P3AX x_out_i0_i41 (.D(\x[1] [8]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_40));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i41.GSR = "ENABLED";
    FD1P3AX x_out_i0_i40 (.D(\x[1] [7]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_39));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i40.GSR = "ENABLED";
    FD1P3AX x_out_i0_i39 (.D(\x[1] [6]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_38));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i39.GSR = "ENABLED";
    FD1P3AX x_out_i0_i38 (.D(\x[1] [5]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_37));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i38.GSR = "ENABLED";
    FD1P3AX x_out_i0_i37 (.D(\x[1] [4]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_36));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i37.GSR = "ENABLED";
    FD1P3AX x_out_i0_i36 (.D(\x[1] [3]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_35));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i36.GSR = "ENABLED";
    FD1P3AX x_out_i0_i35 (.D(\x[1] [2]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_34));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i35.GSR = "ENABLED";
    FD1P3AX x_out_i0_i34 (.D(\x[1] [1]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_33));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i34.GSR = "ENABLED";
    FD1P3AX x_out_i0_i33 (.D(\x[1] [0]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_32));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i33.GSR = "ENABLED";
    FD1P3AX x_out_i0_i32 (.D(\x[0] [31]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_31));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i32.GSR = "ENABLED";
    FD1P3AX x_out_i0_i31 (.D(\x[0] [30]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_30));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i31.GSR = "ENABLED";
    FD1P3AX x_out_i0_i30 (.D(\x[0] [29]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_29));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i30.GSR = "ENABLED";
    FD1P3AX x_out_i0_i29 (.D(\x[0] [28]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_28));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i29.GSR = "ENABLED";
    FD1P3AX x_out_i0_i28 (.D(\x[0] [27]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_27));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i28.GSR = "ENABLED";
    FD1P3AX x_out_i0_i27 (.D(\x[0] [26]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_26));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i27.GSR = "ENABLED";
    FD1P3AX x_out_i0_i26 (.D(\x[0] [25]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_25));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i26.GSR = "ENABLED";
    FD1P3AX x_out_i0_i25 (.D(\x[0] [24]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_24));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i25.GSR = "ENABLED";
    FD1P3AX x_out_i0_i24 (.D(\x[0] [23]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_23));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i24.GSR = "ENABLED";
    FD1P3AX x_out_i0_i23 (.D(\x[0] [22]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_22));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i23.GSR = "ENABLED";
    FD1P3AX x_out_i0_i22 (.D(\x[0] [21]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_21));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i22.GSR = "ENABLED";
    FD1P3AX x_out_i0_i21 (.D(\x[0] [20]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_20));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i21.GSR = "ENABLED";
    FD1P3AX x_out_i0_i20 (.D(\x[0] [19]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_19));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i20.GSR = "ENABLED";
    FD1P3AX x_out_i0_i19 (.D(\x[0] [18]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_18));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i19.GSR = "ENABLED";
    FD1P3AX x_out_i0_i18 (.D(\x[0] [17]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_17));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i18.GSR = "ENABLED";
    FD1P3AX x_out_i0_i17 (.D(\x[0] [16]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_16));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i17.GSR = "ENABLED";
    FD1P3AX x_out_i0_i16 (.D(\x[0] [15]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_15));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i16.GSR = "ENABLED";
    FD1P3AX x_out_i0_i15 (.D(\x[0] [14]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_14));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i15.GSR = "ENABLED";
    FD1P3AX x_out_i0_i14 (.D(\x[0] [13]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_13));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i14.GSR = "ENABLED";
    FD1P3AX x_out_i0_i13 (.D(\x[0] [12]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_12));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i13.GSR = "ENABLED";
    FD1P3AX x_out_i0_i12 (.D(\x[0] [11]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_11));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i12.GSR = "ENABLED";
    FD1P3AX x_out_i0_i11 (.D(\x[0] [10]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_10));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i11.GSR = "ENABLED";
    FD1P3AX x_out_i0_i10 (.D(\x[0] [9]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_9));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i10.GSR = "ENABLED";
    FD1P3AX x_out_i0_i9 (.D(\x[0] [8]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_8));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i9.GSR = "ENABLED";
    FD1P3AX x_out_i0_i8 (.D(\x[0] [7]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_7));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i8.GSR = "ENABLED";
    FD1P3AX x_out_i0_i7 (.D(\x[0] [6]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_6));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i7.GSR = "ENABLED";
    FD1P3AX x_out_i0_i6 (.D(\x[0] [5]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_5));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i6.GSR = "ENABLED";
    FD1P3AX x_out_i0_i5 (.D(\x[0] [4]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_4));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i5.GSR = "ENABLED";
    FD1P3AX x_out_i0_i4 (.D(\x[0] [3]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_3));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i4.GSR = "ENABLED";
    FD1P3AX x_out_i0_i3 (.D(\x[0] [2]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_2));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i3.GSR = "ENABLED";
    FD1P3AX x_out_i0_i2 (.D(\x[0] [1]), .SP(clk_c_enable_677), .CK(clk_c), 
            .Q(x_out_c_1));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_out_i0_i2.GSR = "ENABLED";
    PFUMX div_4016_LessThan_2841_i38 (.BLUT(n14_adj_579), .ALUT(n36_adj_593), 
          .C0(n38948), .Z(n38_adj_595));
    LUT4 i14892_3_lut (.A(U_in_c_152), .B(\U[4] [24]), .C(done_N_1931), 
         .Z(U_0__31__N_967[376])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14892_3_lut.init = 16'hacac;
    PFUMX div_4016_LessThan_2841_i32 (.BLUT(n16_adj_580), .ALUT(n30_adj_589), 
          .C0(n38926), .Z(n32_adj_591));
    LUT4 i1_4_lut_adj_16 (.A(n42812), .B(n37172), .C(n115_adj_223), .D(n117), 
         .Z(n37180)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_16.init = 16'hfffe;
    LUT4 div_4016_LessThan_2681_i45_2_lut_rep_876 (.A(n4085), .B(n117), 
         .Z(n42575)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i45_2_lut_rep_876.init = 16'h6666;
    LUT4 i14890_3_lut (.A(U_in_c_151), .B(\U[4] [23]), .C(done_N_1931), 
         .Z(U_0__31__N_967[375])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14890_3_lut.init = 16'hacac;
    LUT4 div_4016_LessThan_2681_i40_3_lut_3_lut (.A(n4085), .B(n117), .C(n28_adj_528), 
         .Z(n40_adj_536)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_518_i60_4_lut (.A(n132), .B(n131_adj_234), .C(n865), 
         .D(n42787), .Z(n60_adj_795)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_518_i60_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_3066_i26_3_lut_3_lut (.A(n4648), .B(n105), .C(n106_adj_217), 
         .Z(n26_adj_683)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25757_3_lut_4_lut (.A(n4085), .B(n117), .C(n41_adj_537), .D(n42577), 
         .Z(n38677)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25757_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_2681_i47_2_lut_rep_877 (.A(n4084), .B(n116_adj_224), 
         .Z(n42576)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i47_2_lut_rep_877.init = 16'h6666;
    LUT4 i14888_3_lut (.A(U_in_c_150), .B(\U[4] [22]), .C(done_N_1931), 
         .Z(U_0__31__N_967[374])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14888_3_lut.init = 16'hacac;
    LUT4 i14886_3_lut (.A(U_in_c_149), .B(\U[4] [21]), .C(done_N_1931), 
         .Z(U_0__31__N_967[373])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14886_3_lut.init = 16'hacac;
    LUT4 div_4016_LessThan_2681_i26_3_lut_3_lut (.A(n4084), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n26_adj_527)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2681_i43_2_lut_rep_878 (.A(n4086), .B(n118_adj_225), 
         .Z(n42577)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i43_2_lut_rep_878.init = 16'h6666;
    LUT4 div_4016_LessThan_641_i58_4_lut (.A(n132), .B(n131_adj_234), .C(n1049), 
         .D(n42788), .Z(n58)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_641_i58_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2681_i28_3_lut_3_lut (.A(n4086), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n28_adj_528)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i14884_3_lut (.A(U_in_c_148), .B(\U[4] [20]), .C(done_N_1931), 
         .Z(U_0__31__N_967[372])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14884_3_lut.init = 16'hacac;
    LUT4 div_4016_mux_3_i30_3_lut_rep_1085 (.A(n5327), .B(n4_adj_164), .C(n5325), 
         .Z(n42784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i30_3_lut_rep_1085.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i37_2_lut_rep_879 (.A(n4089), .B(n121_adj_227), 
         .Z(n42578)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i37_2_lut_rep_879.init = 16'h6666;
    FD1P3AX i_i0_i31 (.D(i_31__N_1607[31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i31.GSR = "ENABLED";
    FD1P3AX i_i0_i30 (.D(i_31__N_1607[30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i30.GSR = "ENABLED";
    FD1P3AX i_i0_i29 (.D(i_31__N_1607[29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i29.GSR = "ENABLED";
    FD1P3AX i_i0_i28 (.D(i_31__N_1607[28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i28.GSR = "ENABLED";
    FD1P3AX i_i0_i27 (.D(i_31__N_1607[27]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i27.GSR = "ENABLED";
    FD1P3AX i_i0_i26 (.D(i_31__N_1607[26]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i26.GSR = "ENABLED";
    FD1P3AX i_i0_i25 (.D(i_31__N_1607[25]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i25.GSR = "ENABLED";
    FD1P3AX i_i0_i24 (.D(i_31__N_1607[24]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i24.GSR = "ENABLED";
    FD1P3AX i_i0_i23 (.D(i_31__N_1607[23]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i23.GSR = "ENABLED";
    FD1P3AX i_i0_i22 (.D(i_31__N_1607[22]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i22.GSR = "ENABLED";
    FD1P3AX i_i0_i21 (.D(i_31__N_1607[21]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i21.GSR = "ENABLED";
    FD1P3AX i_i0_i20 (.D(i_31__N_1607[20]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i20.GSR = "ENABLED";
    FD1P3AX i_i0_i19 (.D(i_31__N_1607[19]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i19.GSR = "ENABLED";
    FD1P3AX i_i0_i18 (.D(i_31__N_1607[18]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i18.GSR = "ENABLED";
    FD1P3AX i_i0_i17 (.D(i_31__N_1607[17]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i17.GSR = "ENABLED";
    FD1P3AX i_i0_i16 (.D(i_31__N_1607[16]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i16.GSR = "ENABLED";
    FD1P3AX i_i0_i15 (.D(i_31__N_1607[15]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i15.GSR = "ENABLED";
    FD1P3AX i_i0_i14 (.D(i_31__N_1607[14]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i14.GSR = "ENABLED";
    FD1P3AX i_i0_i13 (.D(i_31__N_1607[13]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i13.GSR = "ENABLED";
    FD1P3AX i_i0_i12 (.D(i_31__N_1607[12]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i12.GSR = "ENABLED";
    FD1P3AX i_i0_i11 (.D(i_31__N_1607[11]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i11.GSR = "ENABLED";
    FD1P3AX i_i0_i10 (.D(i_31__N_1607[10]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i10.GSR = "ENABLED";
    FD1P3AX i_i0_i9 (.D(i_31__N_1607[9]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i9.GSR = "ENABLED";
    FD1P3AX i_i0_i8 (.D(i_31__N_1607[8]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i8.GSR = "ENABLED";
    FD1P3AX i_i0_i7 (.D(i_31__N_1607[7]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i7.GSR = "ENABLED";
    FD1P3AX i_i0_i6 (.D(i_31__N_1607[6]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i6.GSR = "ENABLED";
    FD1P3AX i_i0_i5 (.D(i_31__N_1607[5]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i5.GSR = "ENABLED";
    FD1P3AX i_i0_i4 (.D(i_31__N_1607[4]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i4.GSR = "ENABLED";
    FD1P3AX i_i0_i3 (.D(i_31__N_1607[3]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i3.GSR = "ENABLED";
    FD1P3AX i_i0_i2 (.D(i_31__N_1607[2]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(i[2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i2.GSR = "ENABLED";
    LUT4 i14882_3_lut (.A(U_in_c_147), .B(\U[4] [19]), .C(done_N_1931), 
         .Z(U_0__31__N_967[371])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14882_3_lut.init = 16'hacac;
    FD1P3AX y_3___i1 (.D(y_in_c_96), .SP(clk_c_enable_708), .CK(clk_c), 
            .Q(\y[3] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam y_3___i1.GSR = "ENABLED";
    LUT4 div_4016_LessThan_2681_i32_3_lut_3_lut (.A(n4089), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n32_adj_531)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_3_i31_3_lut_rep_1086 (.A(n5326), .B(n3_adj_163), .C(n5325), 
         .Z(n42785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i31_3_lut_rep_1086.init = 16'hcaca;
    L6MUX21 div_4016_LessThan_2762_i62 (.D0(n34_adj_562), .D1(n60_adj_576), 
            .SD(n40108), .Z(n62_adj_577));
    LUT4 div_4016_LessThan_881_i54_4_lut (.A(n132), .B(n131_adj_234), .C(n1408), 
         .D(n683), .Z(n54)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i54_4_lut.init = 16'h0c8e;
    LUT4 i8737_2_lut_4_lut (.A(n5326), .B(n3_adj_163), .C(n5325), .D(n132), 
         .Z(n62_adj_800)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i8737_2_lut_4_lut.init = 16'hcaff;
    CCU2C div_4016_unary_minus_2_add_3_33 (.A0(n5325), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32870), .S0(n2));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_33.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_33.INIT1 = 16'h0000;
    defparam div_4016_unary_minus_2_add_3_33.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_33.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_31 (.A0(n5327), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5326), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32869), .COUT(n32870), .S0(n4_adj_164), .S1(n3_adj_163));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_31.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_31.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_31.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_31.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_29 (.A0(n5329), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5328), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32868), .COUT(n32869), .S0(n6_adj_166), .S1(n5_adj_165));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_29.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_29.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_29.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_29.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_27 (.A0(n5331), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5330), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32867), .COUT(n32868), .S0(n8_adj_168), .S1(n7_adj_167));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_27.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_27.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_27.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_27.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_25 (.A0(n5333), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5332), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32866), .COUT(n32867), .S0(n10_adj_170), .S1(n9_adj_169));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_25.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_25.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_25.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_25.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_23 (.A0(n5335), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5334), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32865), .COUT(n32866), .S0(n12_adj_172), .S1(n11_adj_171));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_23.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_23.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_23.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_23.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_21 (.A0(n5337), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5336), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32864), .COUT(n32865), .S0(n14_adj_174), .S1(n13_adj_173));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_21.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_21.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_21.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_21.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_19 (.A0(n5339), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5338), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32863), .COUT(n32864), .S0(n16_adj_176), .S1(n15_adj_175));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_19.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_19.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_19.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_19.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_17 (.A0(n5341), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5340), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32862), .COUT(n32863), .S0(n18_adj_178), .S1(n17_adj_177));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_17.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_17.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_17.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_17.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_15 (.A0(n5343), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5342), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32861), .COUT(n32862), .S0(n20_adj_180), .S1(n19_adj_179));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_15.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_15.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_15.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_15.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_13 (.A0(n5345), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5344), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32860), .COUT(n32861), .S0(n22_adj_182), .S1(n21_adj_181));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_13.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_13.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_13.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_13.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_11 (.A0(n5347), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5346), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32859), .COUT(n32860), .S0(n24_adj_184), .S1(n23_adj_183));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_11.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_11.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_11.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_11.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_9 (.A0(n5349), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5348), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32858), .COUT(n32859), .S0(n26_adj_186), .S1(n25_adj_185));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_9.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_9.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_9.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_9.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_7 (.A0(n5351), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5350), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32857), .COUT(n32858), .S0(n28_adj_188), .S1(n27_adj_187));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_7.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_7.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_7.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_7.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_5 (.A0(n5353), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5352), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32856), .COUT(n32857), .S0(n30_adj_190), .S1(n29_adj_189));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_5.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_5.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_5.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_5.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_3 (.A0(n5355), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5354), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32855), .COUT(n32856), .S0(n32_adj_192), .S1(n31_adj_191));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_3.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_3.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_2_add_3_3.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_3.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_2_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5356), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32855), .S1(n33_adj_193));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_2_add_3_1.INIT0 = 16'h0000;
    defparam div_4016_unary_minus_2_add_3_1.INIT1 = 16'haaaf;
    defparam div_4016_unary_minus_2_add_3_1.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_2_add_3_1.INJECT1_1 = "NO";
    LUT4 div_4016_i3274_2_lut_rep_1087 (.A(n5325), .B(n5460), .Z(n42786)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3274_2_lut_rep_1087.init = 16'h6666;
    LUT4 i25761_3_lut_4_lut (.A(n4089), .B(n121_adj_227), .C(n35_adj_533), 
         .D(n42579), .Z(n38655)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25761_3_lut_4_lut.init = 16'hfff6;
    PFUMX div_4016_LessThan_2762_i60 (.BLUT(n36_adj_563), .ALUT(n58_adj_575), 
          .C0(n40110), .Z(n60_adj_576));
    LUT4 div_4016_i3341_3_lut_4_lut (.A(n5325), .B(n5460), .C(n22305), 
         .D(n4783), .Z(n5524)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C)+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3341_3_lut_4_lut.init = 16'h60f9;
    LUT4 i14880_3_lut (.A(U_in_c_146), .B(\U[4] [18]), .C(done_N_1931), 
         .Z(U_0__31__N_967[370])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14880_3_lut.init = 16'hacac;
    LUT4 div_4016_i3315_3_lut_4_lut (.A(n5325), .B(n5460), .C(n22279), 
         .D(n1078), .Z(n5498)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C)+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3315_3_lut_4_lut.init = 16'h60f9;
    LUT4 i14878_3_lut (.A(U_in_c_145), .B(\U[4] [17]), .C(done_N_1931), 
         .Z(U_0__31__N_967[369])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14878_3_lut.init = 16'hacac;
    LUT4 div_4016_LessThan_2681_i39_2_lut_rep_880 (.A(n4088), .B(n120), 
         .Z(n42579)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i39_2_lut_rep_880.init = 16'h6666;
    LUT4 div_4016_i3314_3_lut_4_lut (.A(n5325), .B(n5460), .C(n22278), 
         .D(n36422), .Z(n5497)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C)+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3314_3_lut_4_lut.init = 16'h60f9;
    L6MUX21 div_4016_LessThan_2762_i52 (.D0(n40_adj_566), .D1(n50_adj_571), 
            .SD(n38840), .Z(n52_adj_572));
    LUT4 div_4016_LessThan_3066_i61_2_lut_rep_767 (.A(n4647), .B(n104_adj_216), 
         .Z(n42466)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i61_2_lut_rep_767.init = 16'h6666;
    LUT4 div_4016_i3342_3_lut_4_lut (.A(n5325), .B(n5460), .C(n22306), 
         .D(n4885), .Z(n5525)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C)+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3342_3_lut_4_lut.init = 16'h60f9;
    LUT4 i14876_3_lut (.A(U_in_c_144), .B(\U[4] [16]), .C(done_N_1931), 
         .Z(U_0__31__N_967[368])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14876_3_lut.init = 16'hacac;
    LUT4 div_4016_LessThan_2681_i34_3_lut_3_lut (.A(n4088), .B(n120), .C(n32_adj_531), 
         .Z(n34_adj_532)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i14874_3_lut (.A(U_in_c_143), .B(\U[4] [15]), .C(done_N_1931), 
         .Z(U_0__31__N_967[367])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14874_3_lut.init = 16'hacac;
    LUT4 i14872_3_lut (.A(U_in_c_142), .B(\U[4] [14]), .C(done_N_1931), 
         .Z(U_0__31__N_967[366])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14872_3_lut.init = 16'hacac;
    LUT4 i14870_3_lut (.A(U_in_c_141), .B(\U[4] [13]), .C(done_N_1931), 
         .Z(U_0__31__N_967[365])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14870_3_lut.init = 16'hacac;
    LUT4 i14868_3_lut (.A(U_in_c_140), .B(\U[4] [12]), .C(done_N_1931), 
         .Z(U_0__31__N_967[364])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14868_3_lut.init = 16'hacac;
    PFUMX div_4016_LessThan_2762_i50 (.BLUT(n42_adj_567), .ALUT(n48_adj_570), 
          .C0(n38842), .Z(n50_adj_571));
    LUT4 i14866_3_lut (.A(U_in_c_139), .B(\U[4] [11]), .C(done_N_1931), 
         .Z(U_0__31__N_967[363])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14866_3_lut.init = 16'hacac;
    LUT4 i14023_3_lut (.A(U_in_c_138), .B(\U[4] [10]), .C(done_N_1931), 
         .Z(U_0__31__N_967[362])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i14023_3_lut.init = 16'hacac;
    LUT4 i12644_3_lut (.A(U_in_c_137), .B(\U[4] [9]), .C(done_N_1931), 
         .Z(U_0__31__N_967[361])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12644_3_lut.init = 16'hacac;
    LUT4 i12404_3_lut (.A(U_in_c_136), .B(\U[4] [8]), .C(done_N_1931), 
         .Z(U_0__31__N_967[360])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12404_3_lut.init = 16'hacac;
    LUT4 i12402_3_lut (.A(U_in_c_135), .B(\U[4] [7]), .C(done_N_1931), 
         .Z(U_0__31__N_967[359])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12402_3_lut.init = 16'hacac;
    LUT4 i12400_3_lut (.A(U_in_c_134), .B(\U[4] [6]), .C(done_N_1931), 
         .Z(U_0__31__N_967[358])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12400_3_lut.init = 16'hacac;
    LUT4 i12398_3_lut (.A(U_in_c_133), .B(\U[4] [5]), .C(done_N_1931), 
         .Z(U_0__31__N_967[357])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12398_3_lut.init = 16'hacac;
    LUT4 i12396_3_lut (.A(U_in_c_132), .B(\U[4] [4]), .C(done_N_1931), 
         .Z(U_0__31__N_967[356])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12396_3_lut.init = 16'hacac;
    PFUMX div_4016_LessThan_2762_i40 (.BLUT(n16_adj_550), .ALUT(n38_adj_564), 
          .C0(n38808), .Z(n40_adj_566));
    LUT4 i12394_3_lut (.A(U_in_c_131), .B(\U[4] [3]), .C(done_N_1931), 
         .Z(U_0__31__N_967[355])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12394_3_lut.init = 16'hacac;
    LUT4 i12392_3_lut (.A(U_in_c_130), .B(\U[4] [2]), .C(done_N_1931), 
         .Z(U_0__31__N_967[354])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12392_3_lut.init = 16'hacac;
    LUT4 i12390_3_lut (.A(U_in_c_129), .B(\U[4] [1]), .C(done_N_1931), 
         .Z(U_0__31__N_967[353])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12390_3_lut.init = 16'hacac;
    LUT4 i12388_3_lut (.A(U_in_c_128), .B(\U[4] [0]), .C(done_N_1931), 
         .Z(U_0__31__N_967[352])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12388_3_lut.init = 16'hacac;
    LUT4 div_4016_LessThan_2681_i33_2_lut_rep_881 (.A(n4091), .B(n123), 
         .Z(n42580)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i33_2_lut_rep_881.init = 16'h6666;
    LUT4 div_4016_mux_3_i29_3_lut_rep_1088 (.A(n5328), .B(n5_adj_165), .C(n5325), 
         .Z(n42787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i29_3_lut_rep_1088.init = 16'hcaca;
    LUT4 div_4016_LessThan_3066_i54_3_lut_3_lut (.A(n4647), .B(n104_adj_216), 
         .C(n26_adj_683), .Z(n54_adj_698)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25785_4_lut (.A(n42452), .B(n42451), .C(n42454), .D(n39609), 
         .Z(n39634)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25785_4_lut.init = 16'hfeff;
    LUT4 i24349_4_lut (.A(n42453), .B(n42455), .C(n42456), .D(n39593), 
         .Z(n39609)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24349_4_lut.init = 16'h1011;
    LUT4 i24333_4_lut (.A(n42457), .B(n29_adj_719), .C(n17_adj_711), .D(n39546), 
         .Z(n39593)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24333_4_lut.init = 16'h1011;
    PFUMX div_4016_LessThan_2762_i34 (.BLUT(n18_adj_551), .ALUT(n32_adj_560), 
          .C0(n38786), .Z(n34_adj_562));
    LUT4 i25881_4_lut (.A(n42585), .B(n42587), .C(n42586), .D(n42597), 
         .Z(n40100)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25881_4_lut.init = 16'haaab;
    LUT4 i23468_2_lut_3_lut_4_lut (.A(n4091), .B(n123), .C(n111), .D(n4079), 
         .Z(n38728)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23468_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_i3332_4_lut (.A(n64_adj_469), .B(n22296), .C(n42786), 
         .D(n35922), .Z(n5515)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3332_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_2681_i31_2_lut_rep_882 (.A(n4092), .B(n124_adj_229), 
         .Z(n42581)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i31_2_lut_rep_882.init = 16'h6666;
    LUT4 div_4016_mux_3_i28_3_lut_rep_1089 (.A(n5329), .B(n6_adj_166), .C(n5325), 
         .Z(n42788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i28_3_lut_rep_1089.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i22_3_lut_3_lut (.A(n4092), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n22_adj_524)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3066_i55_2_lut_rep_768 (.A(n4650), .B(n107_adj_218), 
         .Z(n42467)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i55_2_lut_rep_768.init = 16'h6666;
    LUT4 div_4016_LessThan_2681_i25_2_lut_rep_883 (.A(n4095), .B(n127_adj_231), 
         .Z(n42582)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i25_2_lut_rep_883.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i48_3_lut_3_lut (.A(n4650), .B(n107_adj_218), 
         .C(n46_adj_694), .Z(n48_adj_695)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2681_i27_2_lut_rep_884 (.A(n4094), .B(n126), 
         .Z(n42583)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i27_2_lut_rep_884.init = 16'h6666;
    LUT4 i23361_2_lut_3_lut_4_lut (.A(n4094), .B(n126), .C(n127_adj_231), 
         .D(n4095), .Z(n38621)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23361_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_i3321_4_lut (.A(n64_adj_278), .B(n22285), .C(n42786), 
         .D(n30893), .Z(n5504)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3321_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_2426_i64_4_lut (.A(n60_adj_467), .B(n62_adj_468), 
         .C(n42619), .D(n38360), .Z(n64_adj_469)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i64_4_lut.init = 16'hccca;
    LUT4 i23100_4_lut (.A(n42621), .B(n42620), .C(n42622), .D(n38335), 
         .Z(n38360)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23100_4_lut.init = 16'h0100;
    LUT4 i23075_4_lut (.A(n42623), .B(n42625), .C(n42624), .D(n38314), 
         .Z(n38335)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23075_4_lut.init = 16'h0100;
    LUT4 i23054_4_lut (.A(n42626), .B(n47_adj_460), .C(n42627), .D(n38297), 
         .Z(n38314)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23054_4_lut.init = 16'h1011;
    LUT4 i23037_4_lut (.A(n42628), .B(n42630), .C(n42629), .D(n38282), 
         .Z(n38297)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23037_4_lut.init = 16'h0100;
    LUT4 i23022_4_lut (.A(n42631), .B(n35_adj_453), .C(n42632), .D(n38269), 
         .Z(n38282)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23022_4_lut.init = 16'h5455;
    LUT4 i23009_4_lut (.A(n42633), .B(n29_adj_449), .C(n42634), .D(n25_adj_446), 
         .Z(n38269)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23009_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_2426_i25_2_lut (.A(n3717), .B(n130_adj_233), 
         .Z(n25_adj_446)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i25_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_17 (.A(n42804), .B(n37298), .C(n42795), .D(n37286), 
         .Z(n35922)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_17.init = 16'hfffe;
    PFUMX div_4016_LessThan_3206_i38 (.BLUT(n30_adj_764), .ALUT(n36_adj_770), 
          .C0(n39991), .Z(n38_adj_772));
    LUT4 i1_2_lut_adj_18 (.A(n108), .B(n110_adj_220), .Z(n37286)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_18.init = 16'heeee;
    LUT4 div_4016_LessThan_2426_i29_2_lut (.A(n3715), .B(n128_adj_232), 
         .Z(n29_adj_449)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i29_2_lut.init = 16'h6666;
    L6MUX21 div_4016_LessThan_2681_i62 (.D0(n36_adj_534), .D1(n60_adj_547), 
            .SD(n40102), .Z(n62_adj_548));
    PFUMX div_4016_LessThan_2681_i60 (.BLUT(n38_adj_535), .ALUT(n58_adj_546), 
          .C0(n40104), .Z(n60_adj_547));
    LUT4 div_4016_LessThan_2426_i35_2_lut (.A(n3712), .B(n125_adj_230), 
         .Z(n35_adj_453)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i35_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_4_lut (.A(n36784), .B(n42792), .C(n36882), .D(n120), 
         .Z(n30896)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_19 (.A(n36992), .B(n42794), .C(n36994), .D(n42806), 
         .Z(n30893)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_19.init = 16'hfffe;
    L6MUX21 div_4016_LessThan_2681_i54 (.D0(n42_adj_538), .D1(n52_adj_543), 
            .SD(n38709), .Z(n54_adj_544));
    LUT4 div_4016_LessThan_2681_i24_3_lut_3_lut (.A(n4094), .B(n126), .C(n127_adj_231), 
         .Z(n24_adj_526)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_998_i52_4_lut (.A(n132), .B(n131_adj_234), .C(n1583), 
         .D(n684), .Z(n52)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i52_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2426_i47_2_lut (.A(n3706), .B(n119_adj_226), 
         .Z(n47_adj_460)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i47_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2681_i21_2_lut_rep_885 (.A(n4097), .B(n129), 
         .Z(n42584)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i21_2_lut_rep_885.init = 16'h6666;
    LUT4 i25783_4_lut (.A(n42452), .B(n42451), .C(n42454), .D(n39618), 
         .Z(n39636)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25783_4_lut.init = 16'hfffe;
    LUT4 div_4016_i3331_4_lut (.A(n64_adj_444), .B(n22295), .C(n42786), 
         .D(n30923), .Z(n5514)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3331_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_2681_i20_3_lut_3_lut (.A(n4097), .B(n129), .C(n130_adj_233), 
         .Z(n20_adj_523)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i20_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_2681_i52 (.BLUT(n44_adj_539), .ALUT(n50_adj_542), 
          .C0(n38711), .Z(n52_adj_543));
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 div_4016_LessThan_2598_i63_2_lut_rep_886 (.A(n3953), .B(n109_adj_219), 
         .Z(n42585)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i63_2_lut_rep_886.init = 16'h6666;
    LUT4 i1_2_lut_4_lut_adj_20 (.A(n42793), .B(n42803), .C(n42796), .D(n108), 
         .Z(n30932)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_20.init = 16'hfffe;
    LUT4 div_4016_LessThan_2598_i58_3_lut_3_lut (.A(n3953), .B(n109_adj_219), 
         .C(n24_adj_496), .Z(n58_adj_517)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25648_4_lut_4_lut (.A(n42589), .B(n38582), .C(n50_adj_513), 
         .D(n26_adj_498), .Z(n52_adj_514)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25648_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i23337_4_lut_4_lut (.A(n42589), .B(n38576), .C(n42586), .D(n42587), 
         .Z(n38597)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23337_4_lut_4_lut.init = 16'h000b;
    LUT4 div_4016_LessThan_2598_i59_2_lut_rep_887 (.A(n3955), .B(n111), 
         .Z(n42586)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i59_2_lut_rep_887.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i32_3_lut_3_lut (.A(n3955), .B(n111), .C(n123), 
         .Z(n32_adj_502)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2337_i64_4_lut (.A(n46_adj_434), .B(n62_adj_443), 
         .C(n42635), .D(n38244), .Z(n64_adj_444)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i64_4_lut.init = 16'hcacc;
    LUT4 i22984_4_lut (.A(n42636), .B(n42638), .C(n42637), .D(n38219), 
         .Z(n38244)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22984_4_lut.init = 16'h0100;
    LUT4 i22959_4_lut (.A(n42640), .B(n42639), .C(n42641), .D(n38204), 
         .Z(n38219)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22959_4_lut.init = 16'h0100;
    PFUMX div_4016_LessThan_2681_i42 (.BLUT(n18_adj_521), .ALUT(n40_adj_536), 
          .C0(n38677), .Z(n42_adj_538));
    LUT4 i22944_4_lut (.A(n49_adj_436), .B(n42643), .C(n42642), .D(n38183), 
         .Z(n38204)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22944_4_lut.init = 16'h5455;
    LUT4 i22923_4_lut (.A(n42645), .B(n42644), .C(n42646), .D(n38170), 
         .Z(n38183)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22923_4_lut.init = 16'h0001;
    LUT4 i22910_4_lut (.A(n37_adj_429), .B(n42648), .C(n42647), .D(n38159), 
         .Z(n38170)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22910_4_lut.init = 16'h0001;
    LUT4 i22899_4_lut (.A(n31_adj_425), .B(n42649), .C(n3584), .D(n130_adj_233), 
         .Z(n38159)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22899_4_lut.init = 16'h1001;
    LUT4 i1_4_lut_adj_21 (.A(n36992), .B(n42793), .C(n42810), .D(n42796), 
         .Z(n30923)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_21.init = 16'hfffe;
    PFUMX div_4016_LessThan_2681_i36 (.BLUT(n20_adj_523), .ALUT(n34_adj_532), 
          .C0(n38655), .Z(n36_adj_534));
    LUT4 i1_3_lut_rep_1090_4_lut (.A(n42798), .B(n42796), .C(n36882), 
         .D(n36784), .Z(n42789)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_rep_1090_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_1113_i50_4_lut (.A(n132), .B(n131_adj_234), .C(n1755), 
         .D(n685), .Z(n50)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i50_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2337_i31_2_lut (.A(n3582), .B(n128_adj_232), 
         .Z(n31_adj_425)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i31_2_lut.init = 16'h6666;
    L6MUX21 div_4016_LessThan_2598_i62 (.D0(n38_adj_506), .D1(n60_adj_518), 
            .SD(n40096), .Z(n62_adj_519));
    LUT4 div_4016_LessThan_2337_i37_2_lut (.A(n3579), .B(n125_adj_230), 
         .Z(n37_adj_429)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i37_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i49_2_lut (.A(n3573), .B(n119_adj_226), 
         .Z(n49_adj_436)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i49_2_lut.init = 16'h6666;
    L6MUX21 div_4016_LessThan_2598_i56 (.D0(n44_adj_510), .D1(n54_adj_515), 
            .SD(n38587), .Z(n56_adj_516));
    FD1P3IX x_3___i117 (.D(n5505), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i117.GSR = "ENABLED";
    PFUMX div_4016_LessThan_2598_i60 (.BLUT(n40_adj_507), .ALUT(n58_adj_517), 
          .C0(n40100), .Z(n60_adj_518));
    LUT4 div_4016_LessThan_3066_i57_2_lut_rep_769 (.A(n4649), .B(n106_adj_217), 
         .Z(n42468)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i57_2_lut_rep_769.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i61_2_lut_rep_888 (.A(n3954), .B(n110_adj_220), 
         .Z(n42587)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i61_2_lut_rep_888.init = 16'h6666;
    FD1P3IX x_3___i118 (.D(n5504), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i118.GSR = "ENABLED";
    PFUMX div_4016_LessThan_2598_i54 (.BLUT(n46_adj_511), .ALUT(n52_adj_514), 
          .C0(n38589), .Z(n54_adj_515));
    LUT4 i24260_2_lut_3_lut_4_lut (.A(n4649), .B(n106_adj_217), .C(n105), 
         .D(n4648), .Z(n39520)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24260_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_1226_i48_4_lut (.A(n132), .B(n131_adj_234), .C(n1924), 
         .D(n872), .Z(n48)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i48_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2598_i40_3_lut_3_lut (.A(n3954), .B(n110_adj_220), 
         .C(n32_adj_502), .Z(n40_adj_507)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2598_i55_2_lut_rep_889 (.A(n3957), .B(n113_adj_222), 
         .Z(n42588)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i55_2_lut_rep_889.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i53_2_lut_rep_770 (.A(n4651), .B(n108), 
         .Z(n42469)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i53_2_lut_rep_770.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i48_3_lut_3_lut (.A(n3957), .B(n113_adj_222), 
         .C(n114), .Z(n48_adj_512)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_3_lut_rep_1091_4_lut (.A(n42798), .B(n42800), .C(n42796), 
         .D(n42803), .Z(n42790)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_rep_1091_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2598_i57_2_lut_rep_890 (.A(n3956), .B(n112_adj_221), 
         .Z(n42589)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i57_2_lut_rep_890.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i50_3_lut_3_lut (.A(n3956), .B(n112_adj_221), 
         .C(n48_adj_512), .Z(n50_adj_513)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25796_4_lut (.A(n42464), .B(n42466), .C(n42465), .D(n39504), 
         .Z(n39525)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25796_4_lut.init = 16'hfeff;
    LUT4 i24244_4_lut (.A(n42468), .B(n42467), .C(n42469), .D(n39480), 
         .Z(n39504)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24244_4_lut.init = 16'h5455;
    LUT4 i24220_4_lut (.A(n42470), .B(n42472), .C(n42471), .D(n39400), 
         .Z(n39480)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24220_4_lut.init = 16'h0001;
    LUT4 i24140_4_lut (.A(n42481), .B(n42480), .C(n25_adj_682), .D(n39386), 
         .Z(n39400)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24140_4_lut.init = 16'h0001;
    PFUMX div_4016_LessThan_2598_i44 (.BLUT(n20_adj_494), .ALUT(n42_adj_508), 
          .C0(n38555), .Z(n44_adj_510));
    LUT4 div_4016_LessThan_3066_i25_2_lut (.A(n4665), .B(n122_adj_228), 
         .Z(n25_adj_682)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i25_2_lut.init = 16'h6666;
    PFUMX div_4016_LessThan_2598_i38 (.BLUT(n22_adj_495), .ALUT(n36_adj_504), 
          .C0(n38533), .Z(n38_adj_506));
    FD1P3IX x_3___i119 (.D(n5503), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i119.GSR = "ENABLED";
    LUT4 div_4016_LessThan_3066_i13_2_lut (.A(n4671), .B(n128_adj_232), 
         .Z(n13_adj_674)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i13_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_4_lut_adj_22 (.A(n42800), .B(n42798), .C(n42796), .D(n106_adj_217), 
         .Z(n30938)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_22.init = 16'hfffe;
    LUT4 div_4016_LessThan_2598_i53_2_lut_rep_891 (.A(n3958), .B(n114), 
         .Z(n42590)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i53_2_lut_rep_891.init = 16'h6666;
    LUT4 i23322_2_lut_3_lut_4_lut (.A(n3958), .B(n114), .C(n113_adj_222), 
         .D(n3957), .Z(n38582)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23322_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2598_i51_2_lut_rep_892 (.A(n3959), .B(n115_adj_223), 
         .Z(n42591)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i51_2_lut_rep_892.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i46_3_lut_3_lut (.A(n4651), .B(n108), .C(n109_adj_219), 
         .Z(n46_adj_694)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i46_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 div_4016_LessThan_2513_i58 (.D0(n46_adj_484), .D1(n56_adj_489), 
            .SD(n38472), .Z(n58_adj_490));
    LUT4 div_4016_LessThan_3066_i51_2_lut_rep_771 (.A(n4652), .B(n109_adj_219), 
         .Z(n42470)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i51_2_lut_rep_771.init = 16'h6666;
    FD1P3IX x_3___i120 (.D(n5502), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i120.GSR = "ENABLED";
    PFUMX div_4016_LessThan_2513_i62 (.BLUT(n40_adj_480), .ALUT(n60_adj_491), 
          .C0(n40092), .Z(n62_adj_492));
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(n42796), .B(n103_adj_215), .C(n36832), 
         .D(n42799), .Z(n37120)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'hfffe;
    LUT4 i24251_4_lut (.A(n42468), .B(n42481), .C(n42480), .D(n25_adj_682), 
         .Z(n39511)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24251_4_lut.init = 16'h5554;
    PFUMX div_4016_LessThan_2513_i56 (.BLUT(n48_adj_485), .ALUT(n54_adj_488), 
          .C0(n38474), .Z(n56_adj_489));
    LUT4 div_4016_i3330_4_lut (.A(n64_adj_421), .B(n22294), .C(n42786), 
         .D(n35925), .Z(n5513)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3330_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_2598_i46_3_lut_3_lut (.A(n3959), .B(n115_adj_223), 
         .C(n28_adj_499), .Z(n46_adj_511)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_3_lut_4_lut (.A(n42796), .B(n103_adj_215), .C(n104_adj_216), 
         .D(n102), .Z(n35961)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23311_3_lut_4_lut (.A(n3959), .B(n115_adj_223), .C(n31_adj_501), 
         .D(n42593), .Z(n38571)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23311_3_lut_4_lut.init = 16'h0009;
    LUT4 i10576_2_lut_rep_1097 (.A(n68_adj_194), .B(n5460), .Z(n42796)) /* synthesis lut_function=(A (B)) */ ;
    defparam i10576_2_lut_rep_1097.init = 16'h8888;
    LUT4 div_4016_LessThan_2598_i47_2_lut_rep_893 (.A(n3961), .B(n117), 
         .Z(n42592)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i47_2_lut_rep_893.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i56_rep_19_3_lut_3_lut_4_lut (.A(n68_adj_194), 
         .B(n5460), .C(n18_adj_752), .D(n42440), .Z(n37379)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam div_4016_LessThan_3206_i56_rep_19_3_lut_3_lut_4_lut.init = 16'h80f8;
    LUT4 div_4016_LessThan_2598_i42_3_lut_3_lut (.A(n3961), .B(n117), .C(n30_adj_500), 
         .Z(n42_adj_508)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24233_2_lut_3_lut_4_lut (.A(n4652), .B(n109_adj_219), .C(n108), 
         .D(n4651), .Z(n39493)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24233_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i25777_3_lut_4_lut (.A(n3961), .B(n117), .C(n43_adj_509), .D(n42594), 
         .Z(n38555)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25777_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_2598_i49_2_lut_rep_894 (.A(n3960), .B(n116_adj_224), 
         .Z(n42593)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i49_2_lut_rep_894.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i28_3_lut_3_lut (.A(n3960), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n28_adj_499)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut (.A(n68_adj_194), .B(n5460), .C(n102), .Z(n30950)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i25710_4_lut_4_lut (.A(n42474), .B(n39451), .C(n38_adj_690), 
         .D(n14_adj_675), .Z(n40_adj_691)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25710_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2246_i64_4_lut (.A(n48_adj_412), .B(n62_adj_420), 
         .C(n42650), .D(n38137), .Z(n64_adj_421)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i64_4_lut.init = 16'hcacc;
    LUT4 i22877_4_lut (.A(n38136), .B(n42651), .C(n42652), .D(n38114), 
         .Z(n38137)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22877_4_lut.init = 16'h0200;
    LUT4 i22854_4_lut (.A(n42653), .B(n42654), .C(n51_adj_414), .D(n38099), 
         .Z(n38114)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22854_4_lut.init = 16'h0001;
    LUT4 i22839_4_lut (.A(n42656), .B(n42655), .C(n42657), .D(n38080), 
         .Z(n38099)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22839_4_lut.init = 16'h0100;
    LUT4 i22820_4_lut (.A(n42658), .B(n42660), .C(n42659), .D(n38067), 
         .Z(n38080)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22820_4_lut.init = 16'h1011;
    PFUMX div_4016_LessThan_2513_i42 (.BLUT(n26_adj_472), .ALUT(n34_adj_477), 
          .C0(n40094), .Z(n42_adj_481));
    LUT4 i22807_4_lut (.A(n42661), .B(n35_adj_405), .C(n33_adj_403), .D(n38058), 
         .Z(n38067)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22807_4_lut.init = 16'h1011;
    LUT4 i1_4_lut_adj_24 (.A(n36832), .B(n42791), .C(n42807), .D(n36818), 
         .Z(n35925)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_24.init = 16'hfffe;
    FD1P3IX x_3___i121 (.D(n5501), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i121.GSR = "ENABLED";
    FD1P3AX U_15___i1 (.D(\U[15] [0]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[15] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i1.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_25 (.A(n110_adj_220), .B(n112_adj_221), .Z(n36818)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_25.init = 16'heeee;
    LUT4 div_4016_LessThan_2598_i45_2_lut_rep_895 (.A(n3962), .B(n118_adj_225), 
         .Z(n42594)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i45_2_lut_rep_895.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i30_3_lut_3_lut (.A(n3962), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n30_adj_500)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_rep_1096_3_lut (.A(n68_adj_194), .B(n5460), .C(n103_adj_215), 
         .Z(n42795)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_1096_3_lut.init = 16'hf8f8;
    LUT4 div_4016_LessThan_2598_i39_2_lut_rep_896 (.A(n3965), .B(n121_adj_227), 
         .Z(n42595)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i39_2_lut_rep_896.init = 16'h6666;
    LUT4 i24206_4_lut_4_lut (.A(n42474), .B(n39445), .C(n42471), .D(n42472), 
         .Z(n39466)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24206_4_lut_4_lut.init = 16'h000b;
    LUT4 i8027_2_lut_3_lut (.A(n68_adj_194), .B(n5460), .C(n64_adj_737), 
         .Z(n4783)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i8027_2_lut_3_lut.init = 16'hf8f8;
    LUT4 div_4016_LessThan_2246_i51_2_lut (.A(n3437), .B(n119_adj_226), 
         .Z(n51_adj_414)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i51_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2246_i61_2_lut (.A(n3432), .B(n114), .Z(n38136)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i61_2_lut.init = 16'h9999;
    LUT4 div_4016_LessThan_2246_i35_2_lut (.A(n3445), .B(n127_adj_231), 
         .Z(n35_adj_405)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i35_2_lut.init = 16'h6666;
    PFUMX div_4016_LessThan_2513_i46 (.BLUT(n22_adj_470), .ALUT(n44_adj_482), 
          .C0(n38440), .Z(n46_adj_484));
    LUT4 div_4016_LessThan_2246_i33_2_lut (.A(n3446), .B(n128_adj_232), 
         .Z(n33_adj_403)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i33_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_26 (.A(n68_adj_194), .B(n5460), .C(n104_adj_216), 
         .D(n42798), .Z(n30944)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_26.init = 16'hfff8;
    LUT4 i1_3_lut_rep_1095_4_lut (.A(n68_adj_194), .B(n5460), .C(n42798), 
         .D(n42800), .Z(n42794)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_rep_1095_4_lut.init = 16'hfff8;
    LUT4 div_4016_LessThan_1337_i46_4_lut (.A(n132), .B(n131_adj_234), .C(n2090), 
         .D(n873), .Z(n46)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i46_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_3066_i47_2_lut_rep_772 (.A(n4654), .B(n111), 
         .Z(n42471)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i47_2_lut_rep_772.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i34_3_lut_3_lut (.A(n3965), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n34_adj_503)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25781_3_lut_4_lut (.A(n3965), .B(n121_adj_227), .C(n37_adj_505), 
         .D(n42596), .Z(n38533)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25781_3_lut_4_lut.init = 16'hfff6;
    LUT4 i25763_4_lut (.A(n42589), .B(n42588), .C(n42590), .D(n38571), 
         .Z(n38589)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25763_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1092_3_lut_4_lut (.A(n68_adj_194), .B(n5460), .C(n42799), 
         .D(n103_adj_215), .Z(n42791)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_rep_1092_3_lut_4_lut.init = 16'hfff8;
    LUT4 div_4016_LessThan_2598_i41_2_lut_rep_897 (.A(n3964), .B(n120), 
         .Z(n42596)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i41_2_lut_rep_897.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i20_3_lut_3_lut (.A(n4654), .B(n111), .C(n123), 
         .Z(n20_adj_679)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25800_4_lut (.A(n42467), .B(n42469), .C(n42470), .D(n39482), 
         .Z(n39500)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25800_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1099 (.A(n103_adj_215), .B(n102), .Z(n42798)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1099.init = 16'heeee;
    LUT4 div_4016_mux_3_i9_3_lut (.A(n5348), .B(n25_adj_185), .C(n5325), 
         .Z(n886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2598_i36_3_lut_3_lut (.A(n3964), .B(n120), .C(n34_adj_503), 
         .Z(n36_adj_504)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i36_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 div_4016_LessThan_2426_i60 (.D0(n48_adj_461), .D1(n58_adj_466), 
            .SD(n38362), .Z(n60_adj_467));
    PFUMX div_4016_LessThan_2426_i58 (.BLUT(n50_adj_462), .ALUT(n56_adj_465), 
          .C0(n38364), .Z(n58_adj_466));
    LUT4 i24222_3_lut_4_lut (.A(n4654), .B(n111), .C(n42482), .D(n42472), 
         .Z(n39482)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24222_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_3066_i49_2_lut_rep_773 (.A(n4653), .B(n110_adj_220), 
         .Z(n42472)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i49_2_lut_rep_773.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i35_2_lut_rep_898 (.A(n3967), .B(n123), 
         .Z(n42597)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i35_2_lut_rep_898.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i28_3_lut_3_lut (.A(n4653), .B(n110_adj_220), 
         .C(n20_adj_679), .Z(n28_adj_684)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25808_4_lut (.A(n42474), .B(n42473), .C(n42475), .D(n39431), 
         .Z(n39456)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25808_4_lut.init = 16'hfeff;
    LUT4 i23257_3_lut_4_lut (.A(n3967), .B(n123), .C(n25_adj_497), .D(n42598), 
         .Z(n38517)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23257_3_lut_4_lut.init = 16'h0009;
    PFUMX div_4016_LessThan_2426_i62 (.BLUT(n42_adj_457), .ALUT(n44_adj_458), 
          .C0(n40090), .Z(n62_adj_468));
    LUT4 div_4016_LessThan_2598_i33_2_lut_rep_899 (.A(n3968), .B(n124_adj_229), 
         .Z(n42598)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i33_2_lut_rep_899.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i24_3_lut_3_lut (.A(n3968), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n24_adj_496)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24171_4_lut (.A(n42476), .B(n42478), .C(n42477), .D(n39415), 
         .Z(n39431)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24171_4_lut.init = 16'h1011;
    LUT4 i24155_4_lut (.A(n42479), .B(n31_adj_686), .C(n19_adj_678), .D(n39368), 
         .Z(n39415)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24155_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_3_lut_4_lut_adj_27 (.A(n103_adj_215), .B(n102), .C(n36992), 
         .D(n42800), .Z(n36606)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_27.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1093_3_lut_4_lut (.A(n103_adj_215), .B(n102), .C(n5460), 
         .D(n68_adj_194), .Z(n42792)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_2_lut_rep_1093_3_lut_4_lut.init = 16'hfeee;
    LUT4 div_4016_LessThan_3066_i31_2_lut (.A(n4662), .B(n119_adj_226), 
         .Z(n31_adj_686)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i31_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i19_2_lut (.A(n4668), .B(n125_adj_230), 
         .Z(n19_adj_678)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i19_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_1100 (.A(n102), .B(n105), .Z(n42799)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1100.init = 16'heeee;
    LUT4 div_4016_LessThan_2598_i27_2_lut_rep_900 (.A(n3971), .B(n127_adj_231), 
         .Z(n42599)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i27_2_lut_rep_900.init = 16'h6666;
    LUT4 div_4016_LessThan_1446_i44_4_lut (.A(n132), .B(n131_adj_234), .C(n2253), 
         .D(n874), .Z(n44)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i44_4_lut.init = 16'h0c8e;
    PFUMX div_4016_LessThan_2426_i48 (.BLUT(n24_adj_445), .ALUT(n46_adj_459), 
          .C0(n38330), .Z(n48_adj_461));
    ALU54B lat_alu_13 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n19191), .SIGNEDIB(n19264), .SIGNEDCIN(GND_net), 
           .A35(n19190), .A34(n19189), .A33(n19188), .A32(n19187), .A31(n19186), 
           .A30(n19185), .A29(n19184), .A28(n19183), .A27(n19182), .A26(n19181), 
           .A25(n19180), .A24(n19179), .A23(n19178), .A22(n19177), .A21(n19176), 
           .A20(n19175), .A19(n19174), .A18(n19173), .A17(n19172), .A16(n19171), 
           .A15(n19170), .A14(n19169), .A13(n19168), .A12(n19167), .A11(n19166), 
           .A10(n19165), .A9(n19164), .A8(n19163), .A7(n19162), .A6(n19161), 
           .A5(n19160), .A4(n19159), .A3(n19158), .A2(n19157), .A1(n19156), 
           .A0(n19155), .B35(n19263), .B34(n19262), .B33(n19261), .B32(n19260), 
           .B31(n19259), .B30(n19258), .B29(n19257), .B28(n19256), .B27(n19255), 
           .B26(n19254), .B25(n19253), .B24(n19252), .B23(n19251), .B22(n19250), 
           .B21(n19249), .B20(n19248), .B19(n19247), .B18(n19246), .B17(n19245), 
           .B16(n19244), .B15(n19243), .B14(n19242), .B13(n19241), .B12(n19240), 
           .B11(n19239), .B10(n19238), .B9(n19237), .B8(n19236), .B7(n19235), 
           .B6(n19234), .B5(n19233), .B4(n19232), .B3(n19231), .B2(n19230), 
           .B1(n19229), .B0(n19228), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n19227), .MA34(n19226), .MA33(n19225), .MA32(n19224), 
           .MA31(n19223), .MA30(n19222), .MA29(n19221), .MA28(n19220), 
           .MA27(n19219), .MA26(n19218), .MA25(n19217), .MA24(n19216), 
           .MA23(n19215), .MA22(n19214), .MA21(n19213), .MA20(n19212), 
           .MA19(n19211), .MA18(n19210), .MA17(n19209), .MA16(n19208), 
           .MA15(n19207), .MA14(n19206), .MA13(n19205), .MA12(n19204), 
           .MA11(n19203), .MA10(n19202), .MA9(n19201), .MA8(n19200), 
           .MA7(n19199), .MA6(n19198), .MA5(n19197), .MA4(n19196), .MA3(n19195), 
           .MA2(n19194), .MA1(n19193), .MA0(n19192), .MB35(n19300), 
           .MB34(n19299), .MB33(n19298), .MB32(n19297), .MB31(n19296), 
           .MB30(n19295), .MB29(n19294), .MB28(n19293), .MB27(n19292), 
           .MB26(n19291), .MB25(n19290), .MB24(n19289), .MB23(n19288), 
           .MB22(n19287), .MB21(n19286), .MB20(n19285), .MB19(n19284), 
           .MB18(n19283), .MB17(n19282), .MB16(n19281), .MB15(n19280), 
           .MB14(n19279), .MB13(n19278), .MB12(n19277), .MB11(n19276), 
           .MB10(n19275), .MB9(n19274), .MB8(n19273), .MB7(n19272), 
           .MB6(n19271), .MB5(n19270), .MB4(n19269), .MB3(n19268), .MB2(n19267), 
           .MB1(n19266), .MB0(n19265), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n19482), 
           .R52(n19481), .R51(n19480), .R50(n19479), .R49(n19478), .R48(n19477), 
           .R47(n19476), .R46(n19475), .R45(n19474), .R44(n19473), .R43(n19472), 
           .R42(n19471), .R41(n19470), .R40(n19469), .R39(n19468), .R38(n19467), 
           .R37(n19466), .R36(n19465), .R35(n19464), .R34(n19463), .R33(n19462), 
           .R32(n19461), .R31(n19460), .R30(n19459), .R29(n19458), .R28(n19457), 
           .R27(n19456), .R26(n19455), .R25(n19454), .R24(n19453), .R23(n19452), 
           .R22(n19451), .R21(n19450), .R20(n19449), .R19(n19448), .R18(n19447), 
           .R17(n177_adj_132), .R16(n178_adj_4), .R15(n179_adj_19), .R14(n180_adj_20), 
           .R13(n181_adj_21), .R12(n182_adj_127), .R11(n183_adj_126), 
           .R10(n184_adj_6), .R9(n185_adj_16), .R8(n186_adj_17), .R7(n187_adj_18), 
           .R6(n188_adj_121), .R5(n189_adj_120), .R4(n190_adj_7), .R3(n191_adj_13), 
           .R2(n192_adj_14), .R1(n193_adj_15), .R0(n194_adj_115), .SIGNEDR(n19483));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[19:38])
    defparam lat_alu_13.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_13.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_13.REG_FLAG_CLK = "NONE";
    defparam lat_alu_13.REG_FLAG_CE = "CE0";
    defparam lat_alu_13.REG_FLAG_RST = "RST0";
    defparam lat_alu_13.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASK01 = "0x00000000000000";
    defparam lat_alu_13.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_13.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_13.CLK0_DIV = "ENABLED";
    defparam lat_alu_13.CLK1_DIV = "ENABLED";
    defparam lat_alu_13.CLK2_DIV = "ENABLED";
    defparam lat_alu_13.CLK3_DIV = "ENABLED";
    defparam lat_alu_13.MCPAT = "0x00000000000000";
    defparam lat_alu_13.MASKPAT = "0x00000000000000";
    defparam lat_alu_13.RNDPAT = "0x00000000000000";
    defparam lat_alu_13.GSR = "ENABLED";
    defparam lat_alu_13.RESETMODE = "SYNC";
    defparam lat_alu_13.MULT9_MODE = "DISABLED";
    defparam lat_alu_13.LEGACY = "DISABLED";
    ALU54B lat_alu_14 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n19337), .SIGNEDIB(n19410), .SIGNEDCIN(n19483), .A35(n19336), 
           .A34(n19335), .A33(n19334), .A32(n19333), .A31(n19332), .A30(n19331), 
           .A29(n19330), .A28(n19329), .A27(n19328), .A26(n19327), .A25(n19326), 
           .A24(n19325), .A23(n19324), .A22(n19323), .A21(n19322), .A20(n19321), 
           .A19(n19320), .A18(n19319), .A17(n19318), .A16(n19317), .A15(n19316), 
           .A14(n19315), .A13(n19314), .A12(n19313), .A11(n19312), .A10(n19311), 
           .A9(n19310), .A8(n19309), .A7(n19308), .A6(n19307), .A5(n19306), 
           .A4(n19305), .A3(n19304), .A2(n19303), .A1(n19302), .A0(n19301), 
           .B35(n19409), .B34(n19408), .B33(n19407), .B32(n19406), .B31(n19405), 
           .B30(n19404), .B29(n19403), .B28(n19402), .B27(n19401), .B26(n19400), 
           .B25(n19399), .B24(n19398), .B23(n19397), .B22(n19396), .B21(n19395), 
           .B20(n19394), .B19(n19393), .B18(n19392), .B17(n19391), .B16(n19390), 
           .B15(n19389), .B14(n19388), .B13(n19387), .B12(n19386), .B11(n19385), 
           .B10(n19384), .B9(n19383), .B8(n19382), .B7(n19381), .B6(n19380), 
           .B5(n19379), .B4(n19378), .B3(n19377), .B2(n19376), .B1(n19375), 
           .B0(n19374), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n19373), .MA34(n19372), .MA33(n19371), .MA32(n19370), 
           .MA31(n19369), .MA30(n19368), .MA29(n19367), .MA28(n19366), 
           .MA27(n19365), .MA26(n19364), .MA25(n19363), .MA24(n19362), 
           .MA23(n19361), .MA22(n19360), .MA21(n19359), .MA20(n19358), 
           .MA19(n19357), .MA18(n19356), .MA17(n19355), .MA16(n19354), 
           .MA15(n19353), .MA14(n19352), .MA13(n19351), .MA12(n19350), 
           .MA11(n19349), .MA10(n19348), .MA9(n19347), .MA8(n19346), 
           .MA7(n19345), .MA6(n19344), .MA5(n19343), .MA4(n19342), .MA3(n19341), 
           .MA2(n19340), .MA1(n19339), .MA0(n19338), .MB35(n19446), 
           .MB34(n19445), .MB33(n19444), .MB32(n19443), .MB31(n19442), 
           .MB30(n19441), .MB29(n19440), .MB28(n19439), .MB27(n19438), 
           .MB26(n19437), .MB25(n19436), .MB24(n19435), .MB23(n19434), 
           .MB22(n19433), .MB21(n19432), .MB20(n19431), .MB19(n19430), 
           .MB18(n19429), .MB17(n19428), .MB16(n19427), .MB15(n19426), 
           .MB14(n19425), .MB13(n19424), .MB12(n19423), .MB11(n19422), 
           .MB10(n19421), .MB9(n19420), .MB8(n19419), .MB7(n19418), 
           .MB6(n19417), .MB5(n19416), .MB4(n19415), .MB3(n19414), .MB2(n19413), 
           .MB1(n19412), .MB0(n19411), .CIN53(n19482), .CIN52(n19481), 
           .CIN51(n19480), .CIN50(n19479), .CIN49(n19478), .CIN48(n19477), 
           .CIN47(n19476), .CIN46(n19475), .CIN45(n19474), .CIN44(n19473), 
           .CIN43(n19472), .CIN42(n19471), .CIN41(n19470), .CIN40(n19469), 
           .CIN39(n19468), .CIN38(n19467), .CIN37(n19466), .CIN36(n19465), 
           .CIN35(n19464), .CIN34(n19463), .CIN33(n19462), .CIN32(n19461), 
           .CIN31(n19460), .CIN30(n19459), .CIN29(n19458), .CIN28(n19457), 
           .CIN27(n19456), .CIN26(n19455), .CIN25(n19454), .CIN24(n19453), 
           .CIN23(n19452), .CIN22(n19451), .CIN21(n19450), .CIN20(n19449), 
           .CIN19(n19448), .CIN18(n19447), .CIN17(n177_adj_132), .CIN16(n178_adj_4), 
           .CIN15(n179_adj_19), .CIN14(n180_adj_20), .CIN13(n181_adj_21), 
           .CIN12(n182_adj_127), .CIN11(n183_adj_126), .CIN10(n184_adj_6), 
           .CIN9(n185_adj_16), .CIN8(n186_adj_17), .CIN7(n187_adj_18), 
           .CIN6(n188_adj_121), .CIN5(n189_adj_120), .CIN4(n190_adj_7), 
           .CIN3(n191_adj_13), .CIN2(n192_adj_14), .CIN1(n193_adj_15), 
           .CIN0(n194_adj_115), .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), 
           .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), 
           .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), 
           .R13(n163_adj_27), .R12(n164_adj_28), .R11(n165_adj_145), .R10(n166_adj_144), 
           .R9(n167_adj_34), .R8(n168_adj_25), .R7(n169_adj_26), .R6(n170_adj_139), 
           .R5(n171_adj_138), .R4(n172), .R3(n173_adj_22), .R2(n174_adj_23), 
           .R1(n175_adj_24), .R0(n176_adj_133));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[19:38])
    defparam lat_alu_14.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_14.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_14.REG_FLAG_CLK = "NONE";
    defparam lat_alu_14.REG_FLAG_CE = "CE0";
    defparam lat_alu_14.REG_FLAG_RST = "RST0";
    defparam lat_alu_14.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASK01 = "0x00000000000000";
    defparam lat_alu_14.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_14.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_14.CLK0_DIV = "ENABLED";
    defparam lat_alu_14.CLK1_DIV = "ENABLED";
    defparam lat_alu_14.CLK2_DIV = "ENABLED";
    defparam lat_alu_14.CLK3_DIV = "ENABLED";
    defparam lat_alu_14.MCPAT = "0x00000000000000";
    defparam lat_alu_14.MASKPAT = "0x00000000000000";
    defparam lat_alu_14.RNDPAT = "0x00000000000000";
    defparam lat_alu_14.GSR = "ENABLED";
    defparam lat_alu_14.RESETMODE = "SYNC";
    defparam lat_alu_14.MULT9_MODE = "DISABLED";
    defparam lat_alu_14.LEGACY = "DISABLED";
    MULT18X18D mult_4006 (.A17(\x[3] [17]), .A16(\x[3] [16]), .A15(\x[3] [15]), 
            .A14(\x[3] [14]), .A13(\x[3] [13]), .A12(\x[3] [12]), .A11(\x[3] [11]), 
            .A10(\x[3] [10]), .A9(\x[3] [9]), .A8(\x[3] [8]), .A7(\x[3] [7]), 
            .A6(\x[3] [6]), .A5(\x[3] [5]), .A4(\x[3] [4]), .A3(\x[3] [3]), 
            .A2(\x[3] [2]), .A1(\x[3] [1]), .A0(\x[3] [0]), .B17(\U[11] [17]), 
            .B16(\U[11] [16]), .B15(\U[11] [15]), .B14(\U[11] [14]), .B13(\U[11] [13]), 
            .B12(\U[11] [12]), .B11(\U[11] [11]), .B10(\U[11] [10]), .B9(\U[11] [9]), 
            .B8(\U[11] [8]), .B7(\U[11] [7]), .B6(\U[11] [6]), .B5(\U[11] [5]), 
            .B4(\U[11] [4]), .B3(\U[11] [3]), .B2(\U[11] [2]), .B1(\U[11] [1]), 
            .B0(\U[11] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19533), 
            .ROA16(n19532), .ROA15(n19531), .ROA14(n19530), .ROA13(n19529), 
            .ROA12(n19528), .ROA11(n19527), .ROA10(n19526), .ROA9(n19525), 
            .ROA8(n19524), .ROA7(n19523), .ROA6(n19522), .ROA5(n19521), 
            .ROA4(n19520), .ROA3(n19519), .ROA2(n19518), .ROA1(n19517), 
            .ROA0(n19516), .ROB17(n19551), .ROB16(n19550), .ROB15(n19549), 
            .ROB14(n19548), .ROB13(n19547), .ROB12(n19546), .ROB11(n19545), 
            .ROB10(n19544), .ROB9(n19543), .ROB8(n19542), .ROB7(n19541), 
            .ROB6(n19540), .ROB5(n19539), .ROB4(n19538), .ROB3(n19537), 
            .ROB2(n19536), .ROB1(n19535), .ROB0(n19534), .P35(n19588), 
            .P34(n19587), .P33(n19586), .P32(n19585), .P31(n19584), 
            .P30(n19583), .P29(n19582), .P28(n19581), .P27(n19580), 
            .P26(n19579), .P25(n19578), .P24(n19577), .P23(n19576), 
            .P22(n19575), .P21(n19574), .P20(n19573), .P19(n19572), 
            .P18(n19571), .P17(n19570), .P16(n19569), .P15(n19568), 
            .P14(n19567), .P13(n19566), .P12(n19565), .P11(n19564), 
            .P10(n19563), .P9(n19562), .P8(n19561), .P7(n19560), .P6(n19559), 
            .P5(n19558), .P4(n19557), .P3(n19556), .P2(n19555), .P1(n19554), 
            .P0(n19553), .SIGNEDP(n19552));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(109[16:35])
    defparam mult_4006.REG_INPUTA_CLK = "NONE";
    defparam mult_4006.REG_INPUTA_CE = "CE0";
    defparam mult_4006.REG_INPUTA_RST = "RST0";
    defparam mult_4006.REG_INPUTB_CLK = "NONE";
    defparam mult_4006.REG_INPUTB_CE = "CE0";
    defparam mult_4006.REG_INPUTB_RST = "RST0";
    defparam mult_4006.REG_INPUTC_CLK = "NONE";
    defparam mult_4006.REG_INPUTC_CE = "CE0";
    defparam mult_4006.REG_INPUTC_RST = "RST0";
    defparam mult_4006.REG_PIPELINE_CLK = "NONE";
    defparam mult_4006.REG_PIPELINE_CE = "CE0";
    defparam mult_4006.REG_PIPELINE_RST = "RST0";
    defparam mult_4006.REG_OUTPUT_CLK = "NONE";
    defparam mult_4006.REG_OUTPUT_CE = "CE0";
    defparam mult_4006.REG_OUTPUT_RST = "RST0";
    defparam mult_4006.CLK0_DIV = "ENABLED";
    defparam mult_4006.CLK1_DIV = "ENABLED";
    defparam mult_4006.CLK2_DIV = "ENABLED";
    defparam mult_4006.CLK3_DIV = "ENABLED";
    defparam mult_4006.HIGHSPEED_CLK = "NONE";
    defparam mult_4006.GSR = "ENABLED";
    defparam mult_4006.CAS_MATCH_REG = "FALSE";
    defparam mult_4006.SOURCEB_MODE = "B_SHIFT";
    defparam mult_4006.MULT_BYPASS = "DISABLED";
    defparam mult_4006.RESETMODE = "SYNC";
    MULT18X18D lat_mult_15 (.A17(\x[3] [31]), .A16(\x[3] [31]), .A15(\x[3] [31]), 
            .A14(\x[3] [31]), .A13(\x[3] [31]), .A12(\x[3] [30]), .A11(\x[3] [29]), 
            .A10(\x[3] [28]), .A9(\x[3] [27]), .A8(\x[3] [26]), .A7(\x[3] [25]), 
            .A6(\x[3] [24]), .A5(\x[3] [23]), .A4(\x[3] [22]), .A3(\x[3] [21]), 
            .A2(\x[3] [20]), .A1(\x[3] [19]), .A0(\x[3] [18]), .B17(\U[11] [17]), 
            .B16(\U[11] [16]), .B15(\U[11] [15]), .B14(\U[11] [14]), .B13(\U[11] [13]), 
            .B12(\U[11] [12]), .B11(\U[11] [11]), .B10(\U[11] [10]), .B9(\U[11] [9]), 
            .B8(\U[11] [8]), .B7(\U[11] [7]), .B6(\U[11] [6]), .B5(\U[11] [5]), 
            .B4(\U[11] [4]), .B3(\U[11] [3]), .B2(\U[11] [2]), .B1(\U[11] [1]), 
            .B0(\U[11] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19606), 
            .ROA16(n19605), .ROA15(n19604), .ROA14(n19603), .ROA13(n19602), 
            .ROA12(n19601), .ROA11(n19600), .ROA10(n19599), .ROA9(n19598), 
            .ROA8(n19597), .ROA7(n19596), .ROA6(n19595), .ROA5(n19594), 
            .ROA4(n19593), .ROA3(n19592), .ROA2(n19591), .ROA1(n19590), 
            .ROA0(n19589), .ROB17(n19624), .ROB16(n19623), .ROB15(n19622), 
            .ROB14(n19621), .ROB13(n19620), .ROB12(n19619), .ROB11(n19618), 
            .ROB10(n19617), .ROB9(n19616), .ROB8(n19615), .ROB7(n19614), 
            .ROB6(n19613), .ROB5(n19612), .ROB4(n19611), .ROB3(n19610), 
            .ROB2(n19609), .ROB1(n19608), .ROB0(n19607), .P35(n19661), 
            .P34(n19660), .P33(n19659), .P32(n19658), .P31(n19657), 
            .P30(n19656), .P29(n19655), .P28(n19654), .P27(n19653), 
            .P26(n19652), .P25(n19651), .P24(n19650), .P23(n19649), 
            .P22(n19648), .P21(n19647), .P20(n19646), .P19(n19645), 
            .P18(n19644), .P17(n19643), .P16(n19642), .P15(n19641), 
            .P14(n19640), .P13(n19639), .P12(n19638), .P11(n19637), 
            .P10(n19636), .P9(n19635), .P8(n19634), .P7(n19633), .P6(n19632), 
            .P5(n19631), .P4(n19630), .P3(n19629), .P2(n19628), .P1(n19627), 
            .P0(n19626), .SIGNEDP(n19625));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(109[16:35])
    defparam lat_mult_15.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTA_CE = "CE0";
    defparam lat_mult_15.REG_INPUTA_RST = "RST0";
    defparam lat_mult_15.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTB_CE = "CE0";
    defparam lat_mult_15.REG_INPUTB_RST = "RST0";
    defparam lat_mult_15.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTC_CE = "CE0";
    defparam lat_mult_15.REG_INPUTC_RST = "RST0";
    defparam lat_mult_15.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_15.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_15.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_15.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_15.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_15.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_15.CLK0_DIV = "ENABLED";
    defparam lat_mult_15.CLK1_DIV = "ENABLED";
    defparam lat_mult_15.CLK2_DIV = "ENABLED";
    defparam lat_mult_15.CLK3_DIV = "ENABLED";
    defparam lat_mult_15.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_15.GSR = "ENABLED";
    defparam lat_mult_15.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_15.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_15.MULT_BYPASS = "DISABLED";
    defparam lat_mult_15.RESETMODE = "SYNC";
    MULT18X18D lat_mult_16 (.A17(\x[3] [17]), .A16(\x[3] [16]), .A15(\x[3] [15]), 
            .A14(\x[3] [14]), .A13(\x[3] [13]), .A12(\x[3] [12]), .A11(\x[3] [11]), 
            .A10(\x[3] [10]), .A9(\x[3] [9]), .A8(\x[3] [8]), .A7(\x[3] [7]), 
            .A6(\x[3] [6]), .A5(\x[3] [5]), .A4(\x[3] [4]), .A3(\x[3] [3]), 
            .A2(\x[3] [2]), .A1(\x[3] [1]), .A0(\x[3] [0]), .B17(\U[11] [31]), 
            .B16(\U[11] [31]), .B15(\U[11] [31]), .B14(\U[11] [31]), .B13(\U[11] [31]), 
            .B12(\U[11] [30]), .B11(\U[11] [29]), .B10(\U[11] [28]), .B9(\U[11] [27]), 
            .B8(\U[11] [26]), .B7(\U[11] [25]), .B6(\U[11] [24]), .B5(\U[11] [23]), 
            .B4(\U[11] [22]), .B3(\U[11] [21]), .B2(\U[11] [20]), .B1(\U[11] [19]), 
            .B0(\U[11] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19679), 
            .ROA16(n19678), .ROA15(n19677), .ROA14(n19676), .ROA13(n19675), 
            .ROA12(n19674), .ROA11(n19673), .ROA10(n19672), .ROA9(n19671), 
            .ROA8(n19670), .ROA7(n19669), .ROA6(n19668), .ROA5(n19667), 
            .ROA4(n19666), .ROA3(n19665), .ROA2(n19664), .ROA1(n19663), 
            .ROA0(n19662), .ROB17(n19697), .ROB16(n19696), .ROB15(n19695), 
            .ROB14(n19694), .ROB13(n19693), .ROB12(n19692), .ROB11(n19691), 
            .ROB10(n19690), .ROB9(n19689), .ROB8(n19688), .ROB7(n19687), 
            .ROB6(n19686), .ROB5(n19685), .ROB4(n19684), .ROB3(n19683), 
            .ROB2(n19682), .ROB1(n19681), .ROB0(n19680), .P35(n19734), 
            .P34(n19733), .P33(n19732), .P32(n19731), .P31(n19730), 
            .P30(n19729), .P29(n19728), .P28(n19727), .P27(n19726), 
            .P26(n19725), .P25(n19724), .P24(n19723), .P23(n19722), 
            .P22(n19721), .P21(n19720), .P20(n19719), .P19(n19718), 
            .P18(n19717), .P17(n19716), .P16(n19715), .P15(n19714), 
            .P14(n19713), .P13(n19712), .P12(n19711), .P11(n19710), 
            .P10(n19709), .P9(n19708), .P8(n19707), .P7(n19706), .P6(n19705), 
            .P5(n19704), .P4(n19703), .P3(n19702), .P2(n19701), .P1(n19700), 
            .P0(n19699), .SIGNEDP(n19698));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(109[16:35])
    defparam lat_mult_16.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTA_CE = "CE0";
    defparam lat_mult_16.REG_INPUTA_RST = "RST0";
    defparam lat_mult_16.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTB_CE = "CE0";
    defparam lat_mult_16.REG_INPUTB_RST = "RST0";
    defparam lat_mult_16.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTC_CE = "CE0";
    defparam lat_mult_16.REG_INPUTC_RST = "RST0";
    defparam lat_mult_16.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_16.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_16.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_16.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_16.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_16.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_16.CLK0_DIV = "ENABLED";
    defparam lat_mult_16.CLK1_DIV = "ENABLED";
    defparam lat_mult_16.CLK2_DIV = "ENABLED";
    defparam lat_mult_16.CLK3_DIV = "ENABLED";
    defparam lat_mult_16.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_16.GSR = "ENABLED";
    defparam lat_mult_16.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_16.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_16.MULT_BYPASS = "DISABLED";
    defparam lat_mult_16.RESETMODE = "SYNC";
    MULT18X18D lat_mult_17 (.A17(\x[3] [31]), .A16(\x[3] [31]), .A15(\x[3] [31]), 
            .A14(\x[3] [31]), .A13(\x[3] [31]), .A12(\x[3] [30]), .A11(\x[3] [29]), 
            .A10(\x[3] [28]), .A9(\x[3] [27]), .A8(\x[3] [26]), .A7(\x[3] [25]), 
            .A6(\x[3] [24]), .A5(\x[3] [23]), .A4(\x[3] [22]), .A3(\x[3] [21]), 
            .A2(\x[3] [20]), .A1(\x[3] [19]), .A0(\x[3] [18]), .B17(\U[11] [31]), 
            .B16(\U[11] [31]), .B15(\U[11] [31]), .B14(\U[11] [31]), .B13(\U[11] [31]), 
            .B12(\U[11] [30]), .B11(\U[11] [29]), .B10(\U[11] [28]), .B9(\U[11] [27]), 
            .B8(\U[11] [26]), .B7(\U[11] [25]), .B6(\U[11] [24]), .B5(\U[11] [23]), 
            .B4(\U[11] [22]), .B3(\U[11] [21]), .B2(\U[11] [20]), .B1(\U[11] [19]), 
            .B0(\U[11] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19752), 
            .ROA16(n19751), .ROA15(n19750), .ROA14(n19749), .ROA13(n19748), 
            .ROA12(n19747), .ROA11(n19746), .ROA10(n19745), .ROA9(n19744), 
            .ROA8(n19743), .ROA7(n19742), .ROA6(n19741), .ROA5(n19740), 
            .ROA4(n19739), .ROA3(n19738), .ROA2(n19737), .ROA1(n19736), 
            .ROA0(n19735), .ROB17(n19770), .ROB16(n19769), .ROB15(n19768), 
            .ROB14(n19767), .ROB13(n19766), .ROB12(n19765), .ROB11(n19764), 
            .ROB10(n19763), .ROB9(n19762), .ROB8(n19761), .ROB7(n19760), 
            .ROB6(n19759), .ROB5(n19758), .ROB4(n19757), .ROB3(n19756), 
            .ROB2(n19755), .ROB1(n19754), .ROB0(n19753), .P35(n19807), 
            .P34(n19806), .P33(n19805), .P32(n19804), .P31(n19803), 
            .P30(n19802), .P29(n19801), .P28(n19800), .P27(n19799), 
            .P26(n19798), .P25(n19797), .P24(n19796), .P23(n19795), 
            .P22(n19794), .P21(n19793), .P20(n19792), .P19(n19791), 
            .P18(n19790), .P17(n19789), .P16(n19788), .P15(n19787), 
            .P14(n19786), .P13(n19785), .P12(n19784), .P11(n19783), 
            .P10(n19782), .P9(n19781), .P8(n19780), .P7(n19779), .P6(n19778), 
            .P5(n19777), .P4(n19776), .P3(n19775), .P2(n19774), .P1(n19773), 
            .P0(n19772), .SIGNEDP(n19771));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(109[16:35])
    defparam lat_mult_17.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTA_CE = "CE0";
    defparam lat_mult_17.REG_INPUTA_RST = "RST0";
    defparam lat_mult_17.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTB_CE = "CE0";
    defparam lat_mult_17.REG_INPUTB_RST = "RST0";
    defparam lat_mult_17.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTC_CE = "CE0";
    defparam lat_mult_17.REG_INPUTC_RST = "RST0";
    defparam lat_mult_17.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_17.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_17.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_17.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_17.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_17.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_17.CLK0_DIV = "ENABLED";
    defparam lat_mult_17.CLK1_DIV = "ENABLED";
    defparam lat_mult_17.CLK2_DIV = "ENABLED";
    defparam lat_mult_17.CLK3_DIV = "ENABLED";
    defparam lat_mult_17.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_17.GSR = "ENABLED";
    defparam lat_mult_17.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_17.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_17.MULT_BYPASS = "DISABLED";
    defparam lat_mult_17.RESETMODE = "SYNC";
    ALU54B lat_alu_18 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n19552), .SIGNEDIB(n19625), .SIGNEDCIN(GND_net), 
           .A35(n19551), .A34(n19550), .A33(n19549), .A32(n19548), .A31(n19547), 
           .A30(n19546), .A29(n19545), .A28(n19544), .A27(n19543), .A26(n19542), 
           .A25(n19541), .A24(n19540), .A23(n19539), .A22(n19538), .A21(n19537), 
           .A20(n19536), .A19(n19535), .A18(n19534), .A17(n19533), .A16(n19532), 
           .A15(n19531), .A14(n19530), .A13(n19529), .A12(n19528), .A11(n19527), 
           .A10(n19526), .A9(n19525), .A8(n19524), .A7(n19523), .A6(n19522), 
           .A5(n19521), .A4(n19520), .A3(n19519), .A2(n19518), .A1(n19517), 
           .A0(n19516), .B35(n19624), .B34(n19623), .B33(n19622), .B32(n19621), 
           .B31(n19620), .B30(n19619), .B29(n19618), .B28(n19617), .B27(n19616), 
           .B26(n19615), .B25(n19614), .B24(n19613), .B23(n19612), .B22(n19611), 
           .B21(n19610), .B20(n19609), .B19(n19608), .B18(n19607), .B17(n19606), 
           .B16(n19605), .B15(n19604), .B14(n19603), .B13(n19602), .B12(n19601), 
           .B11(n19600), .B10(n19599), .B9(n19598), .B8(n19597), .B7(n19596), 
           .B6(n19595), .B5(n19594), .B4(n19593), .B3(n19592), .B2(n19591), 
           .B1(n19590), .B0(n19589), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n19588), .MA34(n19587), .MA33(n19586), .MA32(n19585), 
           .MA31(n19584), .MA30(n19583), .MA29(n19582), .MA28(n19581), 
           .MA27(n19580), .MA26(n19579), .MA25(n19578), .MA24(n19577), 
           .MA23(n19576), .MA22(n19575), .MA21(n19574), .MA20(n19573), 
           .MA19(n19572), .MA18(n19571), .MA17(n19570), .MA16(n19569), 
           .MA15(n19568), .MA14(n19567), .MA13(n19566), .MA12(n19565), 
           .MA11(n19564), .MA10(n19563), .MA9(n19562), .MA8(n19561), 
           .MA7(n19560), .MA6(n19559), .MA5(n19558), .MA4(n19557), .MA3(n19556), 
           .MA2(n19555), .MA1(n19554), .MA0(n19553), .MB35(n19661), 
           .MB34(n19660), .MB33(n19659), .MB32(n19658), .MB31(n19657), 
           .MB30(n19656), .MB29(n19655), .MB28(n19654), .MB27(n19653), 
           .MB26(n19652), .MB25(n19651), .MB24(n19650), .MB23(n19649), 
           .MB22(n19648), .MB21(n19647), .MB20(n19646), .MB19(n19645), 
           .MB18(n19644), .MB17(n19643), .MB16(n19642), .MB15(n19641), 
           .MB14(n19640), .MB13(n19639), .MB12(n19638), .MB11(n19637), 
           .MB10(n19636), .MB9(n19635), .MB8(n19634), .MB7(n19633), 
           .MB6(n19632), .MB5(n19631), .MB4(n19630), .MB3(n19629), .MB2(n19628), 
           .MB1(n19627), .MB0(n19626), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n19843), 
           .R52(n19842), .R51(n19841), .R50(n19840), .R49(n19839), .R48(n19838), 
           .R47(n19837), .R46(n19836), .R45(n19835), .R44(n19834), .R43(n19833), 
           .R42(n19832), .R41(n19831), .R40(n19830), .R39(n19829), .R38(n19828), 
           .R37(n19827), .R36(n19826), .R35(n19825), .R34(n19824), .R33(n19823), 
           .R32(n19822), .R31(n19821), .R30(n19820), .R29(n19819), .R28(n19818), 
           .R27(n19817), .R26(n19816), .R25(n19815), .R24(n19814), .R23(n19813), 
           .R22(n19812), .R21(n19811), .R20(n19810), .R19(n19809), .R18(n19808), 
           .R17(n5207), .R16(n5208), .R15(n5209), .R14(n5210), .R13(n5211), 
           .R12(n5212), .R11(n5213), .R10(n5214), .R9(n5215), .R8(n5216), 
           .R7(n5217), .R6(n5218), .R5(n5219), .R4(n5220), .R3(n5221), 
           .R2(n5222), .R1(n5223), .R0(n5224), .SIGNEDR(n19844));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(109[16:35])
    defparam lat_alu_18.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_18.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_18.REG_FLAG_CLK = "NONE";
    defparam lat_alu_18.REG_FLAG_CE = "CE0";
    defparam lat_alu_18.REG_FLAG_RST = "RST0";
    defparam lat_alu_18.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASK01 = "0x00000000000000";
    defparam lat_alu_18.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_18.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_18.CLK0_DIV = "ENABLED";
    defparam lat_alu_18.CLK1_DIV = "ENABLED";
    defparam lat_alu_18.CLK2_DIV = "ENABLED";
    defparam lat_alu_18.CLK3_DIV = "ENABLED";
    defparam lat_alu_18.MCPAT = "0x00000000000000";
    defparam lat_alu_18.MASKPAT = "0x00000000000000";
    defparam lat_alu_18.RNDPAT = "0x00000000000000";
    defparam lat_alu_18.GSR = "ENABLED";
    defparam lat_alu_18.RESETMODE = "SYNC";
    defparam lat_alu_18.MULT9_MODE = "DISABLED";
    defparam lat_alu_18.LEGACY = "DISABLED";
    ALU54B lat_alu_19 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n19698), .SIGNEDIB(n19771), .SIGNEDCIN(n19844), .A35(n19697), 
           .A34(n19696), .A33(n19695), .A32(n19694), .A31(n19693), .A30(n19692), 
           .A29(n19691), .A28(n19690), .A27(n19689), .A26(n19688), .A25(n19687), 
           .A24(n19686), .A23(n19685), .A22(n19684), .A21(n19683), .A20(n19682), 
           .A19(n19681), .A18(n19680), .A17(n19679), .A16(n19678), .A15(n19677), 
           .A14(n19676), .A13(n19675), .A12(n19674), .A11(n19673), .A10(n19672), 
           .A9(n19671), .A8(n19670), .A7(n19669), .A6(n19668), .A5(n19667), 
           .A4(n19666), .A3(n19665), .A2(n19664), .A1(n19663), .A0(n19662), 
           .B35(n19770), .B34(n19769), .B33(n19768), .B32(n19767), .B31(n19766), 
           .B30(n19765), .B29(n19764), .B28(n19763), .B27(n19762), .B26(n19761), 
           .B25(n19760), .B24(n19759), .B23(n19758), .B22(n19757), .B21(n19756), 
           .B20(n19755), .B19(n19754), .B18(n19753), .B17(n19752), .B16(n19751), 
           .B15(n19750), .B14(n19749), .B13(n19748), .B12(n19747), .B11(n19746), 
           .B10(n19745), .B9(n19744), .B8(n19743), .B7(n19742), .B6(n19741), 
           .B5(n19740), .B4(n19739), .B3(n19738), .B2(n19737), .B1(n19736), 
           .B0(n19735), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n19734), .MA34(n19733), .MA33(n19732), .MA32(n19731), 
           .MA31(n19730), .MA30(n19729), .MA29(n19728), .MA28(n19727), 
           .MA27(n19726), .MA26(n19725), .MA25(n19724), .MA24(n19723), 
           .MA23(n19722), .MA22(n19721), .MA21(n19720), .MA20(n19719), 
           .MA19(n19718), .MA18(n19717), .MA17(n19716), .MA16(n19715), 
           .MA15(n19714), .MA14(n19713), .MA13(n19712), .MA12(n19711), 
           .MA11(n19710), .MA10(n19709), .MA9(n19708), .MA8(n19707), 
           .MA7(n19706), .MA6(n19705), .MA5(n19704), .MA4(n19703), .MA3(n19702), 
           .MA2(n19701), .MA1(n19700), .MA0(n19699), .MB35(n19807), 
           .MB34(n19806), .MB33(n19805), .MB32(n19804), .MB31(n19803), 
           .MB30(n19802), .MB29(n19801), .MB28(n19800), .MB27(n19799), 
           .MB26(n19798), .MB25(n19797), .MB24(n19796), .MB23(n19795), 
           .MB22(n19794), .MB21(n19793), .MB20(n19792), .MB19(n19791), 
           .MB18(n19790), .MB17(n19789), .MB16(n19788), .MB15(n19787), 
           .MB14(n19786), .MB13(n19785), .MB12(n19784), .MB11(n19783), 
           .MB10(n19782), .MB9(n19781), .MB8(n19780), .MB7(n19779), 
           .MB6(n19778), .MB5(n19777), .MB4(n19776), .MB3(n19775), .MB2(n19774), 
           .MB1(n19773), .MB0(n19772), .CIN53(n19843), .CIN52(n19842), 
           .CIN51(n19841), .CIN50(n19840), .CIN49(n19839), .CIN48(n19838), 
           .CIN47(n19837), .CIN46(n19836), .CIN45(n19835), .CIN44(n19834), 
           .CIN43(n19833), .CIN42(n19832), .CIN41(n19831), .CIN40(n19830), 
           .CIN39(n19829), .CIN38(n19828), .CIN37(n19827), .CIN36(n19826), 
           .CIN35(n19825), .CIN34(n19824), .CIN33(n19823), .CIN32(n19822), 
           .CIN31(n19821), .CIN30(n19820), .CIN29(n19819), .CIN28(n19818), 
           .CIN27(n19817), .CIN26(n19816), .CIN25(n19815), .CIN24(n19814), 
           .CIN23(n19813), .CIN22(n19812), .CIN21(n19811), .CIN20(n19810), 
           .CIN19(n19809), .CIN18(n19808), .CIN17(n5207), .CIN16(n5208), 
           .CIN15(n5209), .CIN14(n5210), .CIN13(n5211), .CIN12(n5212), 
           .CIN11(n5213), .CIN10(n5214), .CIN9(n5215), .CIN8(n5216), 
           .CIN7(n5217), .CIN6(n5218), .CIN5(n5219), .CIN4(n5220), .CIN3(n5221), 
           .CIN2(n5222), .CIN1(n5223), .CIN0(n5224), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(n5193), .R12(n5194), .R11(n5195), 
           .R10(n5196), .R9(n5197), .R8(n5198), .R7(n5199), .R6(n5200), 
           .R5(n5201), .R4(n5202), .R3(n5203), .R2(n5204), .R1(n5205), 
           .R0(n5206));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(109[16:35])
    defparam lat_alu_19.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_19.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_19.REG_FLAG_CLK = "NONE";
    defparam lat_alu_19.REG_FLAG_CE = "CE0";
    defparam lat_alu_19.REG_FLAG_RST = "RST0";
    defparam lat_alu_19.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASK01 = "0x00000000000000";
    defparam lat_alu_19.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_19.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_19.CLK0_DIV = "ENABLED";
    defparam lat_alu_19.CLK1_DIV = "ENABLED";
    defparam lat_alu_19.CLK2_DIV = "ENABLED";
    defparam lat_alu_19.CLK3_DIV = "ENABLED";
    defparam lat_alu_19.MCPAT = "0x00000000000000";
    defparam lat_alu_19.MASKPAT = "0x00000000000000";
    defparam lat_alu_19.RNDPAT = "0x00000000000000";
    defparam lat_alu_19.GSR = "ENABLED";
    defparam lat_alu_19.RESETMODE = "SYNC";
    defparam lat_alu_19.MULT9_MODE = "DISABLED";
    defparam lat_alu_19.LEGACY = "DISABLED";
    MULT18X18D mult_4001_mult_2 (.A17(\U[7] [17]), .A16(\U[7] [16]), .A15(\U[7] [15]), 
            .A14(\U[7] [14]), .A13(\U[7] [13]), .A12(\U[7] [12]), .A11(\U[7] [11]), 
            .A10(\U[7] [10]), .A9(\U[7] [9]), .A8(\U[7] [8]), .A7(\U[7] [7]), 
            .A6(\U[7] [6]), .A5(\U[7] [5]), .A4(\U[7] [4]), .A3(\U[7] [3]), 
            .A2(\U[7] [2]), .A1(\U[7] [1]), .A0(\U[7] [0]), .B17(\x[3] [17]), 
            .B16(\x[3] [16]), .B15(\x[3] [15]), .B14(\x[3] [14]), .B13(\x[3] [13]), 
            .B12(\x[3] [12]), .B11(\x[3] [11]), .B10(\x[3] [10]), .B9(\x[3] [9]), 
            .B8(\x[3] [8]), .B7(\x[3] [7]), .B6(\x[3] [6]), .B5(\x[3] [5]), 
            .B4(\x[3] [4]), .B3(\x[3] [3]), .B2(\x[3] [2]), .B1(\x[3] [1]), 
            .B0(\x[3] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n19894), 
            .ROA16(n19893), .ROA15(n19892), .ROA14(n19891), .ROA13(n19890), 
            .ROA12(n19889), .ROA11(n19888), .ROA10(n19887), .ROA9(n19886), 
            .ROA8(n19885), .ROA7(n19884), .ROA6(n19883), .ROA5(n19882), 
            .ROA4(n19881), .ROA3(n19880), .ROA2(n19879), .ROA1(n19878), 
            .ROA0(n19877), .ROB17(n19912), .ROB16(n19911), .ROB15(n19910), 
            .ROB14(n19909), .ROB13(n19908), .ROB12(n19907), .ROB11(n19906), 
            .ROB10(n19905), .ROB9(n19904), .ROB8(n19903), .ROB7(n19902), 
            .ROB6(n19901), .ROB5(n19900), .ROB4(n19899), .ROB3(n19898), 
            .ROB2(n19897), .ROB1(n19896), .ROB0(n19895), .P35(n19949), 
            .P34(n19948), .P33(n19947), .P32(n19946), .P31(n19945), 
            .P30(n19944), .P29(n19943), .P28(n19942), .P27(n19941), 
            .P26(n19940), .P25(n19939), .P24(n19938), .P23(n19937), 
            .P22(n19936), .P21(n19935), .P20(n19934), .P19(n19933), 
            .P18(n19932), .P17(n19931), .P16(n19930), .P15(n19929), 
            .P14(n19928), .P13(n19927), .P12(n19926), .P11(n19925), 
            .P10(n19924), .P9(n19923), .P8(n19922), .P7(n19921), .P6(n19920), 
            .P5(n19919), .P4(n19918), .P3(n19917), .P2(n19916), .P1(n19915), 
            .P0(n19914), .SIGNEDP(n19913));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(106[16:35])
    defparam mult_4001_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_4001_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_4001_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_4001_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_4001_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_4001_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_4001_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_4001_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_4001_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_4001_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_4001_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_4001_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_4001_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_4001_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_4001_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_4001_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_4001_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_4001_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_4001_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_4001_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_4001_mult_2.GSR = "ENABLED";
    defparam mult_4001_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_4001_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_4001_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_4001_mult_2.RESETMODE = "SYNC";
    MULT18X18D lat_mult_5 (.A17(\U[3] [31]), .A16(\U[3] [31]), .A15(\U[3] [31]), 
            .A14(\U[3] [31]), .A13(\U[3] [31]), .A12(\U[3] [30]), .A11(\U[3] [29]), 
            .A10(\U[3] [28]), .A9(\U[3] [27]), .A8(\U[3] [26]), .A7(\U[3] [25]), 
            .A6(\U[3] [24]), .A5(\U[3] [23]), .A4(\U[3] [22]), .A3(\U[3] [21]), 
            .A2(\U[3] [20]), .A1(\U[3] [19]), .A0(\U[3] [18]), .B17(\x[3] [17]), 
            .B16(\x[3] [16]), .B15(\x[3] [15]), .B14(\x[3] [14]), .B13(\x[3] [13]), 
            .B12(\x[3] [12]), .B11(\x[3] [11]), .B10(\x[3] [10]), .B9(\x[3] [9]), 
            .B8(\x[3] [8]), .B7(\x[3] [7]), .B6(\x[3] [6]), .B5(\x[3] [5]), 
            .B4(\x[3] [4]), .B3(\x[3] [3]), .B2(\x[3] [2]), .B1(\x[3] [1]), 
            .B0(\x[3] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18884), 
            .ROA16(n18883), .ROA15(n18882), .ROA14(n18881), .ROA13(n18880), 
            .ROA12(n18879), .ROA11(n18878), .ROA10(n18877), .ROA9(n18876), 
            .ROA8(n18875), .ROA7(n18874), .ROA6(n18873), .ROA5(n18872), 
            .ROA4(n18871), .ROA3(n18870), .ROA2(n18869), .ROA1(n18868), 
            .ROA0(n18867), .ROB17(n18902), .ROB16(n18901), .ROB15(n18900), 
            .ROB14(n18899), .ROB13(n18898), .ROB12(n18897), .ROB11(n18896), 
            .ROB10(n18895), .ROB9(n18894), .ROB8(n18893), .ROB7(n18892), 
            .ROB6(n18891), .ROB5(n18890), .ROB4(n18889), .ROB3(n18888), 
            .ROB2(n18887), .ROB1(n18886), .ROB0(n18885), .P35(n18939), 
            .P34(n18938), .P33(n18937), .P32(n18936), .P31(n18935), 
            .P30(n18934), .P29(n18933), .P28(n18932), .P27(n18931), 
            .P26(n18930), .P25(n18929), .P24(n18928), .P23(n18927), 
            .P22(n18926), .P21(n18925), .P20(n18924), .P19(n18923), 
            .P18(n18922), .P17(n18921), .P16(n18920), .P15(n18919), 
            .P14(n18918), .P13(n18917), .P12(n18916), .P11(n18915), 
            .P10(n18914), .P9(n18913), .P8(n18912), .P7(n18911), .P6(n18910), 
            .P5(n18909), .P4(n18908), .P3(n18907), .P2(n18906), .P1(n18905), 
            .P0(n18904), .SIGNEDP(n18903));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(102[16:35])
    defparam lat_mult_5.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTA_CE = "CE0";
    defparam lat_mult_5.REG_INPUTA_RST = "RST0";
    defparam lat_mult_5.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTB_CE = "CE0";
    defparam lat_mult_5.REG_INPUTB_RST = "RST0";
    defparam lat_mult_5.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTC_CE = "CE0";
    defparam lat_mult_5.REG_INPUTC_RST = "RST0";
    defparam lat_mult_5.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_5.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_5.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_5.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_5.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_5.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_5.CLK0_DIV = "ENABLED";
    defparam lat_mult_5.CLK1_DIV = "ENABLED";
    defparam lat_mult_5.CLK2_DIV = "ENABLED";
    defparam lat_mult_5.CLK3_DIV = "ENABLED";
    defparam lat_mult_5.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_5.GSR = "ENABLED";
    defparam lat_mult_5.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_5.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_5.MULT_BYPASS = "DISABLED";
    defparam lat_mult_5.RESETMODE = "SYNC";
    MULT18X18D lat_mult_22 (.A17(\U[7] [31]), .A16(\U[7] [31]), .A15(\U[7] [31]), 
            .A14(\U[7] [31]), .A13(\U[7] [31]), .A12(\U[7] [30]), .A11(\U[7] [29]), 
            .A10(\U[7] [28]), .A9(\U[7] [27]), .A8(\U[7] [26]), .A7(\U[7] [25]), 
            .A6(\U[7] [24]), .A5(\U[7] [23]), .A4(\U[7] [22]), .A3(\U[7] [21]), 
            .A2(\U[7] [20]), .A1(\U[7] [19]), .A0(\U[7] [18]), .B17(\x[3] [31]), 
            .B16(\x[3] [31]), .B15(\x[3] [31]), .B14(\x[3] [31]), .B13(\x[3] [31]), 
            .B12(\x[3] [30]), .B11(\x[3] [29]), .B10(\x[3] [28]), .B9(\x[3] [27]), 
            .B8(\x[3] [26]), .B7(\x[3] [25]), .B6(\x[3] [24]), .B5(\x[3] [23]), 
            .B4(\x[3] [22]), .B3(\x[3] [21]), .B2(\x[3] [20]), .B1(\x[3] [19]), 
            .B0(\x[3] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n20113), 
            .ROA16(n20112), .ROA15(n20111), .ROA14(n20110), .ROA13(n20109), 
            .ROA12(n20108), .ROA11(n20107), .ROA10(n20106), .ROA9(n20105), 
            .ROA8(n20104), .ROA7(n20103), .ROA6(n20102), .ROA5(n20101), 
            .ROA4(n20100), .ROA3(n20099), .ROA2(n20098), .ROA1(n20097), 
            .ROA0(n20096), .ROB17(n20131), .ROB16(n20130), .ROB15(n20129), 
            .ROB14(n20128), .ROB13(n20127), .ROB12(n20126), .ROB11(n20125), 
            .ROB10(n20124), .ROB9(n20123), .ROB8(n20122), .ROB7(n20121), 
            .ROB6(n20120), .ROB5(n20119), .ROB4(n20118), .ROB3(n20117), 
            .ROB2(n20116), .ROB1(n20115), .ROB0(n20114), .P35(n20168), 
            .P34(n20167), .P33(n20166), .P32(n20165), .P31(n20164), 
            .P30(n20163), .P29(n20162), .P28(n20161), .P27(n20160), 
            .P26(n20159), .P25(n20158), .P24(n20157), .P23(n20156), 
            .P22(n20155), .P21(n20154), .P20(n20153), .P19(n20152), 
            .P18(n20151), .P17(n20150), .P16(n20149), .P15(n20148), 
            .P14(n20147), .P13(n20146), .P12(n20145), .P11(n20144), 
            .P10(n20143), .P9(n20142), .P8(n20141), .P7(n20140), .P6(n20139), 
            .P5(n20138), .P4(n20137), .P3(n20136), .P2(n20135), .P1(n20134), 
            .P0(n20133), .SIGNEDP(n20132));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(106[16:35])
    defparam lat_mult_22.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_22.REG_INPUTA_CE = "CE0";
    defparam lat_mult_22.REG_INPUTA_RST = "RST0";
    defparam lat_mult_22.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_22.REG_INPUTB_CE = "CE0";
    defparam lat_mult_22.REG_INPUTB_RST = "RST0";
    defparam lat_mult_22.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_22.REG_INPUTC_CE = "CE0";
    defparam lat_mult_22.REG_INPUTC_RST = "RST0";
    defparam lat_mult_22.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_22.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_22.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_22.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_22.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_22.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_22.CLK0_DIV = "ENABLED";
    defparam lat_mult_22.CLK1_DIV = "ENABLED";
    defparam lat_mult_22.CLK2_DIV = "ENABLED";
    defparam lat_mult_22.CLK3_DIV = "ENABLED";
    defparam lat_mult_22.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_22.GSR = "ENABLED";
    defparam lat_mult_22.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_22.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_22.MULT_BYPASS = "DISABLED";
    defparam lat_mult_22.RESETMODE = "SYNC";
    MULT18X18D lat_mult_2 (.A17(\U[2] [31]), .A16(\U[2] [31]), .A15(\U[2] [31]), 
            .A14(\U[2] [31]), .A13(\U[2] [31]), .A12(\U[2] [30]), .A11(\U[2] [29]), 
            .A10(\U[2] [28]), .A9(\U[2] [27]), .A8(\U[2] [26]), .A7(\U[2] [25]), 
            .A6(\U[2] [24]), .A5(\U[2] [23]), .A4(\U[2] [22]), .A3(\U[2] [21]), 
            .A2(\U[2] [20]), .A1(\U[2] [19]), .A0(\U[2] [18]), .B17(\x[2] [31]), 
            .B16(\x[2] [31]), .B15(\x[2] [31]), .B14(\x[2] [31]), .B13(\x[2] [31]), 
            .B12(\x[2] [30]), .B11(\x[2] [29]), .B10(\x[2] [28]), .B9(\x[2] [27]), 
            .B8(\x[2] [26]), .B7(\x[2] [25]), .B6(\x[2] [24]), .B5(\x[2] [23]), 
            .B4(\x[2] [22]), .B3(\x[2] [21]), .B2(\x[2] [20]), .B1(\x[2] [19]), 
            .B0(\x[2] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18669), 
            .ROA16(n18668), .ROA15(n18667), .ROA14(n18666), .ROA13(n18665), 
            .ROA12(n18664), .ROA11(n18663), .ROA10(n18662), .ROA9(n18661), 
            .ROA8(n18660), .ROA7(n18659), .ROA6(n18658), .ROA5(n18657), 
            .ROA4(n18656), .ROA3(n18655), .ROA2(n18654), .ROA1(n18653), 
            .ROA0(n18652), .ROB17(n18687), .ROB16(n18686), .ROB15(n18685), 
            .ROB14(n18684), .ROB13(n18683), .ROB12(n18682), .ROB11(n18681), 
            .ROB10(n18680), .ROB9(n18679), .ROB8(n18678), .ROB7(n18677), 
            .ROB6(n18676), .ROB5(n18675), .ROB4(n18674), .ROB3(n18673), 
            .ROB2(n18672), .ROB1(n18671), .ROB0(n18670), .P35(n18724), 
            .P34(n18723), .P33(n18722), .P32(n18721), .P31(n18720), 
            .P30(n18719), .P29(n18718), .P28(n18717), .P27(n18716), 
            .P26(n18715), .P25(n18714), .P24(n18713), .P23(n18712), 
            .P22(n18711), .P21(n18710), .P20(n18709), .P19(n18708), 
            .P18(n18707), .P17(n18706), .P16(n18705), .P15(n18704), 
            .P14(n18703), .P13(n18702), .P12(n18701), .P11(n18700), 
            .P10(n18699), .P9(n18698), .P8(n18697), .P7(n18696), .P6(n18695), 
            .P5(n18694), .P4(n18693), .P3(n18692), .P2(n18691), .P1(n18690), 
            .P0(n18689), .SIGNEDP(n18688));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[16:35])
    defparam lat_mult_2.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTA_CE = "CE0";
    defparam lat_mult_2.REG_INPUTA_RST = "RST0";
    defparam lat_mult_2.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTB_CE = "CE0";
    defparam lat_mult_2.REG_INPUTB_RST = "RST0";
    defparam lat_mult_2.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTC_CE = "CE0";
    defparam lat_mult_2.REG_INPUTC_RST = "RST0";
    defparam lat_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_2.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_2.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_2.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_2.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_2.CLK0_DIV = "ENABLED";
    defparam lat_mult_2.CLK1_DIV = "ENABLED";
    defparam lat_mult_2.CLK2_DIV = "ENABLED";
    defparam lat_mult_2.CLK3_DIV = "ENABLED";
    defparam lat_mult_2.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_2.GSR = "ENABLED";
    defparam lat_mult_2.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_2.MULT_BYPASS = "DISABLED";
    defparam lat_mult_2.RESETMODE = "SYNC";
    LUT4 div_4016_mux_3_i14_3_lut (.A(n5343), .B(n20_adj_180), .C(n5325), 
         .Z(n881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i14_3_lut.init = 16'hcaca;
    LUT4 div_4016_i3329_4_lut (.A(n64_adj_399), .B(n22293), .C(n42786), 
         .D(n30917), .Z(n5512)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3329_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_3066_i43_2_lut_rep_774 (.A(n4656), .B(n113_adj_222), 
         .Z(n42473)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i43_2_lut_rep_774.init = 16'h6666;
    ALU54B lat_alu_23 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n19913), .SIGNEDIB(n19986), .SIGNEDCIN(GND_net), 
           .A35(n19912), .A34(n19911), .A33(n19910), .A32(n19909), .A31(n19908), 
           .A30(n19907), .A29(n19906), .A28(n19905), .A27(n19904), .A26(n19903), 
           .A25(n19902), .A24(n19901), .A23(n19900), .A22(n19899), .A21(n19898), 
           .A20(n19897), .A19(n19896), .A18(n19895), .A17(n19894), .A16(n19893), 
           .A15(n19892), .A14(n19891), .A13(n19890), .A12(n19889), .A11(n19888), 
           .A10(n19887), .A9(n19886), .A8(n19885), .A7(n19884), .A6(n19883), 
           .A5(n19882), .A4(n19881), .A3(n19880), .A2(n19879), .A1(n19878), 
           .A0(n19877), .B35(n19985), .B34(n19984), .B33(n19983), .B32(n19982), 
           .B31(n19981), .B30(n19980), .B29(n19979), .B28(n19978), .B27(n19977), 
           .B26(n19976), .B25(n19975), .B24(n19974), .B23(n19973), .B22(n19972), 
           .B21(n19971), .B20(n19970), .B19(n19969), .B18(n19968), .B17(n19967), 
           .B16(n19966), .B15(n19965), .B14(n19964), .B13(n19963), .B12(n19962), 
           .B11(n19961), .B10(n19960), .B9(n19959), .B8(n19958), .B7(n19957), 
           .B6(n19956), .B5(n19955), .B4(n19954), .B3(n19953), .B2(n19952), 
           .B1(n19951), .B0(n19950), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n19949), .MA34(n19948), .MA33(n19947), .MA32(n19946), 
           .MA31(n19945), .MA30(n19944), .MA29(n19943), .MA28(n19942), 
           .MA27(n19941), .MA26(n19940), .MA25(n19939), .MA24(n19938), 
           .MA23(n19937), .MA22(n19936), .MA21(n19935), .MA20(n19934), 
           .MA19(n19933), .MA18(n19932), .MA17(n19931), .MA16(n19930), 
           .MA15(n19929), .MA14(n19928), .MA13(n19927), .MA12(n19926), 
           .MA11(n19925), .MA10(n19924), .MA9(n19923), .MA8(n19922), 
           .MA7(n19921), .MA6(n19920), .MA5(n19919), .MA4(n19918), .MA3(n19917), 
           .MA2(n19916), .MA1(n19915), .MA0(n19914), .MB35(n20022), 
           .MB34(n20021), .MB33(n20020), .MB32(n20019), .MB31(n20018), 
           .MB30(n20017), .MB29(n20016), .MB28(n20015), .MB27(n20014), 
           .MB26(n20013), .MB25(n20012), .MB24(n20011), .MB23(n20010), 
           .MB22(n20009), .MB21(n20008), .MB20(n20007), .MB19(n20006), 
           .MB18(n20005), .MB17(n20004), .MB16(n20003), .MB15(n20002), 
           .MB14(n20001), .MB13(n20000), .MB12(n19999), .MB11(n19998), 
           .MB10(n19997), .MB9(n19996), .MB8(n19995), .MB7(n19994), 
           .MB6(n19993), .MB5(n19992), .MB4(n19991), .MB3(n19990), .MB2(n19989), 
           .MB1(n19988), .MB0(n19987), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n20204), 
           .R52(n20203), .R51(n20202), .R50(n20201), .R49(n20200), .R48(n20199), 
           .R47(n20198), .R46(n20197), .R45(n20196), .R44(n20195), .R43(n20194), 
           .R42(n20193), .R41(n20192), .R40(n20191), .R39(n20190), .R38(n20189), 
           .R37(n20188), .R36(n20187), .R35(n20186), .R34(n20185), .R33(n20184), 
           .R32(n20183), .R31(n20182), .R30(n20181), .R29(n20180), .R28(n20179), 
           .R27(n20178), .R26(n20177), .R25(n20176), .R24(n20175), .R23(n20174), 
           .R22(n20173), .R21(n20172), .R20(n20171), .R19(n20170), .R18(n20169), 
           .R17(n177_adj_40), .R16(n178_adj_39), .R15(n179_adj_89), .R14(n180_adj_88), 
           .R13(n181_adj_31), .R12(n182_adj_112), .R11(n183_adj_111), 
           .R10(n184_adj_110), .R9(n185_adj_109), .R8(n186_adj_108), .R7(n187_adj_51), 
           .R6(n188_adj_93), .R5(n189_adj_86), .R4(n190_adj_35), .R3(n191_adj_47), 
           .R2(n192_adj_42), .R1(n193_adj_44), .R0(n194_adj_48), .SIGNEDR(n20205));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(106[16:35])
    defparam lat_alu_23.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_23.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_23.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_23.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_23.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_23.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_23.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_23.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_23.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_23.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_23.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_23.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_23.REG_FLAG_CLK = "NONE";
    defparam lat_alu_23.REG_FLAG_CE = "CE0";
    defparam lat_alu_23.REG_FLAG_RST = "RST0";
    defparam lat_alu_23.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_23.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_23.MASK01 = "0x00000000000000";
    defparam lat_alu_23.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_23.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_23.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_23.CLK0_DIV = "ENABLED";
    defparam lat_alu_23.CLK1_DIV = "ENABLED";
    defparam lat_alu_23.CLK2_DIV = "ENABLED";
    defparam lat_alu_23.CLK3_DIV = "ENABLED";
    defparam lat_alu_23.MCPAT = "0x00000000000000";
    defparam lat_alu_23.MASKPAT = "0x00000000000000";
    defparam lat_alu_23.RNDPAT = "0x00000000000000";
    defparam lat_alu_23.GSR = "ENABLED";
    defparam lat_alu_23.RESETMODE = "SYNC";
    defparam lat_alu_23.MULT9_MODE = "DISABLED";
    defparam lat_alu_23.LEGACY = "DISABLED";
    MULT18X18D lat_mult_1 (.A17(\U[2] [17]), .A16(\U[2] [16]), .A15(\U[2] [15]), 
            .A14(\U[2] [14]), .A13(\U[2] [13]), .A12(\U[2] [12]), .A11(\U[2] [11]), 
            .A10(\U[2] [10]), .A9(\U[2] [9]), .A8(\U[2] [8]), .A7(\U[2] [7]), 
            .A6(\U[2] [6]), .A5(\U[2] [5]), .A4(\U[2] [4]), .A3(\U[2] [3]), 
            .A2(\U[2] [2]), .A1(\U[2] [1]), .A0(\U[2] [0]), .B17(\x[2] [31]), 
            .B16(\x[2] [31]), .B15(\x[2] [31]), .B14(\x[2] [31]), .B13(\x[2] [31]), 
            .B12(\x[2] [30]), .B11(\x[2] [29]), .B10(\x[2] [28]), .B9(\x[2] [27]), 
            .B8(\x[2] [26]), .B7(\x[2] [25]), .B6(\x[2] [24]), .B5(\x[2] [23]), 
            .B4(\x[2] [22]), .B3(\x[2] [21]), .B2(\x[2] [20]), .B1(\x[2] [19]), 
            .B0(\x[2] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18596), 
            .ROA16(n18595), .ROA15(n18594), .ROA14(n18593), .ROA13(n18592), 
            .ROA12(n18591), .ROA11(n18590), .ROA10(n18589), .ROA9(n18588), 
            .ROA8(n18587), .ROA7(n18586), .ROA6(n18585), .ROA5(n18584), 
            .ROA4(n18583), .ROA3(n18582), .ROA2(n18581), .ROA1(n18580), 
            .ROA0(n18579), .ROB17(n18614), .ROB16(n18613), .ROB15(n18612), 
            .ROB14(n18611), .ROB13(n18610), .ROB12(n18609), .ROB11(n18608), 
            .ROB10(n18607), .ROB9(n18606), .ROB8(n18605), .ROB7(n18604), 
            .ROB6(n18603), .ROB5(n18602), .ROB4(n18601), .ROB3(n18600), 
            .ROB2(n18599), .ROB1(n18598), .ROB0(n18597), .P35(n18651), 
            .P34(n18650), .P33(n18649), .P32(n18648), .P31(n18647), 
            .P30(n18646), .P29(n18645), .P28(n18644), .P27(n18643), 
            .P26(n18642), .P25(n18641), .P24(n18640), .P23(n18639), 
            .P22(n18638), .P21(n18637), .P20(n18636), .P19(n18635), 
            .P18(n18634), .P17(n18633), .P16(n18632), .P15(n18631), 
            .P14(n18630), .P13(n18629), .P12(n18628), .P11(n18627), 
            .P10(n18626), .P9(n18625), .P8(n18624), .P7(n18623), .P6(n18622), 
            .P5(n18621), .P4(n18620), .P3(n18619), .P2(n18618), .P1(n18617), 
            .P0(n18616), .SIGNEDP(n18615));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[16:35])
    defparam lat_mult_1.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTA_CE = "CE0";
    defparam lat_mult_1.REG_INPUTA_RST = "RST0";
    defparam lat_mult_1.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTB_CE = "CE0";
    defparam lat_mult_1.REG_INPUTB_RST = "RST0";
    defparam lat_mult_1.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTC_CE = "CE0";
    defparam lat_mult_1.REG_INPUTC_RST = "RST0";
    defparam lat_mult_1.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_1.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_1.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_1.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_1.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_1.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_1.CLK0_DIV = "ENABLED";
    defparam lat_mult_1.CLK1_DIV = "ENABLED";
    defparam lat_mult_1.CLK2_DIV = "ENABLED";
    defparam lat_mult_1.CLK3_DIV = "ENABLED";
    defparam lat_mult_1.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_1.GSR = "ENABLED";
    defparam lat_mult_1.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_1.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_1.MULT_BYPASS = "DISABLED";
    defparam lat_mult_1.RESETMODE = "SYNC";
    ALU54B lat_alu_24 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n20059), .SIGNEDIB(n20132), .SIGNEDCIN(n20205), .A35(n20058), 
           .A34(n20057), .A33(n20056), .A32(n20055), .A31(n20054), .A30(n20053), 
           .A29(n20052), .A28(n20051), .A27(n20050), .A26(n20049), .A25(n20048), 
           .A24(n20047), .A23(n20046), .A22(n20045), .A21(n20044), .A20(n20043), 
           .A19(n20042), .A18(n20041), .A17(n20040), .A16(n20039), .A15(n20038), 
           .A14(n20037), .A13(n20036), .A12(n20035), .A11(n20034), .A10(n20033), 
           .A9(n20032), .A8(n20031), .A7(n20030), .A6(n20029), .A5(n20028), 
           .A4(n20027), .A3(n20026), .A2(n20025), .A1(n20024), .A0(n20023), 
           .B35(n20131), .B34(n20130), .B33(n20129), .B32(n20128), .B31(n20127), 
           .B30(n20126), .B29(n20125), .B28(n20124), .B27(n20123), .B26(n20122), 
           .B25(n20121), .B24(n20120), .B23(n20119), .B22(n20118), .B21(n20117), 
           .B20(n20116), .B19(n20115), .B18(n20114), .B17(n20113), .B16(n20112), 
           .B15(n20111), .B14(n20110), .B13(n20109), .B12(n20108), .B11(n20107), 
           .B10(n20106), .B9(n20105), .B8(n20104), .B7(n20103), .B6(n20102), 
           .B5(n20101), .B4(n20100), .B3(n20099), .B2(n20098), .B1(n20097), 
           .B0(n20096), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n20095), .MA34(n20094), .MA33(n20093), .MA32(n20092), 
           .MA31(n20091), .MA30(n20090), .MA29(n20089), .MA28(n20088), 
           .MA27(n20087), .MA26(n20086), .MA25(n20085), .MA24(n20084), 
           .MA23(n20083), .MA22(n20082), .MA21(n20081), .MA20(n20080), 
           .MA19(n20079), .MA18(n20078), .MA17(n20077), .MA16(n20076), 
           .MA15(n20075), .MA14(n20074), .MA13(n20073), .MA12(n20072), 
           .MA11(n20071), .MA10(n20070), .MA9(n20069), .MA8(n20068), 
           .MA7(n20067), .MA6(n20066), .MA5(n20065), .MA4(n20064), .MA3(n20063), 
           .MA2(n20062), .MA1(n20061), .MA0(n20060), .MB35(n20168), 
           .MB34(n20167), .MB33(n20166), .MB32(n20165), .MB31(n20164), 
           .MB30(n20163), .MB29(n20162), .MB28(n20161), .MB27(n20160), 
           .MB26(n20159), .MB25(n20158), .MB24(n20157), .MB23(n20156), 
           .MB22(n20155), .MB21(n20154), .MB20(n20153), .MB19(n20152), 
           .MB18(n20151), .MB17(n20150), .MB16(n20149), .MB15(n20148), 
           .MB14(n20147), .MB13(n20146), .MB12(n20145), .MB11(n20144), 
           .MB10(n20143), .MB9(n20142), .MB8(n20141), .MB7(n20140), 
           .MB6(n20139), .MB5(n20138), .MB4(n20137), .MB3(n20136), .MB2(n20135), 
           .MB1(n20134), .MB0(n20133), .CIN53(n20204), .CIN52(n20203), 
           .CIN51(n20202), .CIN50(n20201), .CIN49(n20200), .CIN48(n20199), 
           .CIN47(n20198), .CIN46(n20197), .CIN45(n20196), .CIN44(n20195), 
           .CIN43(n20194), .CIN42(n20193), .CIN41(n20192), .CIN40(n20191), 
           .CIN39(n20190), .CIN38(n20189), .CIN37(n20188), .CIN36(n20187), 
           .CIN35(n20186), .CIN34(n20185), .CIN33(n20184), .CIN32(n20183), 
           .CIN31(n20182), .CIN30(n20181), .CIN29(n20180), .CIN28(n20179), 
           .CIN27(n20178), .CIN26(n20177), .CIN25(n20176), .CIN24(n20175), 
           .CIN23(n20174), .CIN22(n20173), .CIN21(n20172), .CIN20(n20171), 
           .CIN19(n20170), .CIN18(n20169), .CIN17(n177_adj_40), .CIN16(n178_adj_39), 
           .CIN15(n179_adj_89), .CIN14(n180_adj_88), .CIN13(n181_adj_31), 
           .CIN12(n182_adj_112), .CIN11(n183_adj_111), .CIN10(n184_adj_110), 
           .CIN9(n185_adj_109), .CIN8(n186_adj_108), .CIN7(n187_adj_51), 
           .CIN6(n188_adj_93), .CIN5(n189_adj_86), .CIN4(n190_adj_35), 
           .CIN3(n191_adj_47), .CIN2(n192_adj_42), .CIN1(n193_adj_44), 
           .CIN0(n194_adj_48), .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), 
           .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), 
           .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), 
           .R13(n163_adj_107), .R12(n164_adj_97), .R11(n165_adj_105), 
           .R10(n166_adj_33), .R9(n167_adj_32), .R8(n168_adj_46), .R7(n169_adj_37), 
           .R6(n170_adj_43), .R5(n171_adj_36), .R4(n172_adj_45), .R3(n173_adj_30), 
           .R2(n174_adj_29), .R1(n175_adj_38), .R0(n176_adj_41));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(106[16:35])
    defparam lat_alu_24.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_24.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_24.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_24.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_24.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_24.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_24.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_24.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_24.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_24.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_24.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_24.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_24.REG_FLAG_CLK = "NONE";
    defparam lat_alu_24.REG_FLAG_CE = "CE0";
    defparam lat_alu_24.REG_FLAG_RST = "RST0";
    defparam lat_alu_24.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_24.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_24.MASK01 = "0x00000000000000";
    defparam lat_alu_24.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_24.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_24.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_24.CLK0_DIV = "ENABLED";
    defparam lat_alu_24.CLK1_DIV = "ENABLED";
    defparam lat_alu_24.CLK2_DIV = "ENABLED";
    defparam lat_alu_24.CLK3_DIV = "ENABLED";
    defparam lat_alu_24.MCPAT = "0x00000000000000";
    defparam lat_alu_24.MASKPAT = "0x00000000000000";
    defparam lat_alu_24.RNDPAT = "0x00000000000000";
    defparam lat_alu_24.GSR = "ENABLED";
    defparam lat_alu_24.RESETMODE = "SYNC";
    defparam lat_alu_24.MULT9_MODE = "DISABLED";
    defparam lat_alu_24.LEGACY = "DISABLED";
    MULT18X18D mult_3998_mult_2 (.A17(\U[1] [17]), .A16(\U[1] [16]), .A15(\U[1] [15]), 
            .A14(\U[1] [14]), .A13(\U[1] [13]), .A12(\U[1] [12]), .A11(\U[1] [11]), 
            .A10(\U[1] [10]), .A9(\U[1] [9]), .A8(\U[1] [8]), .A7(\U[1] [7]), 
            .A6(\U[1] [6]), .A5(\U[1] [5]), .A4(\U[1] [4]), .A3(\U[1] [3]), 
            .A2(\U[1] [2]), .A1(\U[1] [1]), .A0(\U[1] [0]), .B17(\x[1] [17]), 
            .B16(\x[1] [16]), .B15(\x[1] [15]), .B14(\x[1] [14]), .B13(\x[1] [13]), 
            .B12(\x[1] [12]), .B11(\x[1] [11]), .B10(\x[1] [10]), .B9(\x[1] [9]), 
            .B8(\x[1] [8]), .B7(\x[1] [7]), .B6(\x[1] [6]), .B5(\x[1] [5]), 
            .B4(\x[1] [4]), .B3(\x[1] [3]), .B2(\x[1] [2]), .B1(\x[1] [1]), 
            .B0(\x[1] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n20255), 
            .ROA16(n20254), .ROA15(n20253), .ROA14(n20252), .ROA13(n20251), 
            .ROA12(n20250), .ROA11(n20249), .ROA10(n20248), .ROA9(n20247), 
            .ROA8(n20246), .ROA7(n20245), .ROA6(n20244), .ROA5(n20243), 
            .ROA4(n20242), .ROA3(n20241), .ROA2(n20240), .ROA1(n20239), 
            .ROA0(n20238), .ROB17(n20273), .ROB16(n20272), .ROB15(n20271), 
            .ROB14(n20270), .ROB13(n20269), .ROB12(n20268), .ROB11(n20267), 
            .ROB10(n20266), .ROB9(n20265), .ROB8(n20264), .ROB7(n20263), 
            .ROB6(n20262), .ROB5(n20261), .ROB4(n20260), .ROB3(n20259), 
            .ROB2(n20258), .ROB1(n20257), .ROB0(n20256), .P35(n20310), 
            .P34(n20309), .P33(n20308), .P32(n20307), .P31(n20306), 
            .P30(n20305), .P29(n20304), .P28(n20303), .P27(n20302), 
            .P26(n20301), .P25(n20300), .P24(n20299), .P23(n20298), 
            .P22(n20297), .P21(n20296), .P20(n20295), .P19(n20294), 
            .P18(n20293), .P17(n20292), .P16(n20291), .P15(n20290), 
            .P14(n20289), .P13(n20288), .P12(n20287), .P11(n20286), 
            .P10(n20285), .P9(n20284), .P8(n20283), .P7(n20282), .P6(n20281), 
            .P5(n20280), .P4(n20279), .P3(n20278), .P2(n20277), .P1(n20276), 
            .P0(n20275), .SIGNEDP(n20274));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(104[16:35])
    defparam mult_3998_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_3998_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_3998_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_3998_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_3998_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_3998_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_3998_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_3998_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_3998_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_3998_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_3998_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_3998_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_3998_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_3998_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_3998_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_3998_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_3998_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_3998_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_3998_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_3998_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_3998_mult_2.GSR = "ENABLED";
    defparam mult_3998_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_3998_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_3998_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_3998_mult_2.RESETMODE = "SYNC";
    MULT18X18D mult_3994_mult_2 (.A17(\U[3] [17]), .A16(\U[3] [16]), .A15(\U[3] [15]), 
            .A14(\U[3] [14]), .A13(\U[3] [13]), .A12(\U[3] [12]), .A11(\U[3] [11]), 
            .A10(\U[3] [10]), .A9(\U[3] [9]), .A8(\U[3] [8]), .A7(\U[3] [7]), 
            .A6(\U[3] [6]), .A5(\U[3] [5]), .A4(\U[3] [4]), .A3(\U[3] [3]), 
            .A2(\U[3] [2]), .A1(\U[3] [1]), .A0(\U[3] [0]), .B17(\x[3] [17]), 
            .B16(\x[3] [16]), .B15(\x[3] [15]), .B14(\x[3] [14]), .B13(\x[3] [13]), 
            .B12(\x[3] [12]), .B11(\x[3] [11]), .B10(\x[3] [10]), .B9(\x[3] [9]), 
            .B8(\x[3] [8]), .B7(\x[3] [7]), .B6(\x[3] [6]), .B5(\x[3] [5]), 
            .B4(\x[3] [4]), .B3(\x[3] [3]), .B2(\x[3] [2]), .B1(\x[3] [1]), 
            .B0(\x[3] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18811), 
            .ROA16(n18810), .ROA15(n18809), .ROA14(n18808), .ROA13(n18807), 
            .ROA12(n18806), .ROA11(n18805), .ROA10(n18804), .ROA9(n18803), 
            .ROA8(n18802), .ROA7(n18801), .ROA6(n18800), .ROA5(n18799), 
            .ROA4(n18798), .ROA3(n18797), .ROA2(n18796), .ROA1(n18795), 
            .ROA0(n18794), .ROB17(n18829), .ROB16(n18828), .ROB15(n18827), 
            .ROB14(n18826), .ROB13(n18825), .ROB12(n18824), .ROB11(n18823), 
            .ROB10(n18822), .ROB9(n18821), .ROB8(n18820), .ROB7(n18819), 
            .ROB6(n18818), .ROB5(n18817), .ROB4(n18816), .ROB3(n18815), 
            .ROB2(n18814), .ROB1(n18813), .ROB0(n18812), .P35(n18866), 
            .P34(n18865), .P33(n18864), .P32(n18863), .P31(n18862), 
            .P30(n18861), .P29(n18860), .P28(n18859), .P27(n18858), 
            .P26(n18857), .P25(n18856), .P24(n18855), .P23(n18854), 
            .P22(n18853), .P21(n18852), .P20(n18851), .P19(n18850), 
            .P18(n18849), .P17(n18848), .P16(n18847), .P15(n18846), 
            .P14(n18845), .P13(n18844), .P12(n18843), .P11(n18842), 
            .P10(n18841), .P9(n18840), .P8(n18839), .P7(n18838), .P6(n18837), 
            .P5(n18836), .P4(n18835), .P3(n18834), .P2(n18833), .P1(n18832), 
            .P0(n18831), .SIGNEDP(n18830));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(102[16:35])
    defparam mult_3994_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_3994_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_3994_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_3994_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_3994_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_3994_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_3994_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_3994_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_3994_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_3994_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_3994_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_3994_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_3994_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_3994_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_3994_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_3994_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_3994_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_3994_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_3994_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_3994_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_3994_mult_2.GSR = "ENABLED";
    defparam mult_3994_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_3994_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_3994_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_3994_mult_2.RESETMODE = "SYNC";
    MULT18X18D lat_mult_25 (.A17(\U[1] [31]), .A16(\U[1] [31]), .A15(\U[1] [31]), 
            .A14(\U[1] [31]), .A13(\U[1] [31]), .A12(\U[1] [30]), .A11(\U[1] [29]), 
            .A10(\U[1] [28]), .A9(\U[1] [27]), .A8(\U[1] [26]), .A7(\U[1] [25]), 
            .A6(\U[1] [24]), .A5(\U[1] [23]), .A4(\U[1] [22]), .A3(\U[1] [21]), 
            .A2(\U[1] [20]), .A1(\U[1] [19]), .A0(\U[1] [18]), .B17(\x[1] [17]), 
            .B16(\x[1] [16]), .B15(\x[1] [15]), .B14(\x[1] [14]), .B13(\x[1] [13]), 
            .B12(\x[1] [12]), .B11(\x[1] [11]), .B10(\x[1] [10]), .B9(\x[1] [9]), 
            .B8(\x[1] [8]), .B7(\x[1] [7]), .B6(\x[1] [6]), .B5(\x[1] [5]), 
            .B4(\x[1] [4]), .B3(\x[1] [3]), .B2(\x[1] [2]), .B1(\x[1] [1]), 
            .B0(\x[1] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n20328), 
            .ROA16(n20327), .ROA15(n20326), .ROA14(n20325), .ROA13(n20324), 
            .ROA12(n20323), .ROA11(n20322), .ROA10(n20321), .ROA9(n20320), 
            .ROA8(n20319), .ROA7(n20318), .ROA6(n20317), .ROA5(n20316), 
            .ROA4(n20315), .ROA3(n20314), .ROA2(n20313), .ROA1(n20312), 
            .ROA0(n20311), .ROB17(n20346), .ROB16(n20345), .ROB15(n20344), 
            .ROB14(n20343), .ROB13(n20342), .ROB12(n20341), .ROB11(n20340), 
            .ROB10(n20339), .ROB9(n20338), .ROB8(n20337), .ROB7(n20336), 
            .ROB6(n20335), .ROB5(n20334), .ROB4(n20333), .ROB3(n20332), 
            .ROB2(n20331), .ROB1(n20330), .ROB0(n20329), .P35(n20383), 
            .P34(n20382), .P33(n20381), .P32(n20380), .P31(n20379), 
            .P30(n20378), .P29(n20377), .P28(n20376), .P27(n20375), 
            .P26(n20374), .P25(n20373), .P24(n20372), .P23(n20371), 
            .P22(n20370), .P21(n20369), .P20(n20368), .P19(n20367), 
            .P18(n20366), .P17(n20365), .P16(n20364), .P15(n20363), 
            .P14(n20362), .P13(n20361), .P12(n20360), .P11(n20359), 
            .P10(n20358), .P9(n20357), .P8(n20356), .P7(n20355), .P6(n20354), 
            .P5(n20353), .P4(n20352), .P3(n20351), .P2(n20350), .P1(n20349), 
            .P0(n20348), .SIGNEDP(n20347));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(104[16:35])
    defparam lat_mult_25.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_25.REG_INPUTA_CE = "CE0";
    defparam lat_mult_25.REG_INPUTA_RST = "RST0";
    defparam lat_mult_25.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_25.REG_INPUTB_CE = "CE0";
    defparam lat_mult_25.REG_INPUTB_RST = "RST0";
    defparam lat_mult_25.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_25.REG_INPUTC_CE = "CE0";
    defparam lat_mult_25.REG_INPUTC_RST = "RST0";
    defparam lat_mult_25.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_25.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_25.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_25.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_25.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_25.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_25.CLK0_DIV = "ENABLED";
    defparam lat_mult_25.CLK1_DIV = "ENABLED";
    defparam lat_mult_25.CLK2_DIV = "ENABLED";
    defparam lat_mult_25.CLK3_DIV = "ENABLED";
    defparam lat_mult_25.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_25.GSR = "ENABLED";
    defparam lat_mult_25.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_25.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_25.MULT_BYPASS = "DISABLED";
    defparam lat_mult_25.RESETMODE = "SYNC";
    MULT18X18D lat_mult_26 (.A17(\U[1] [17]), .A16(\U[1] [16]), .A15(\U[1] [15]), 
            .A14(\U[1] [14]), .A13(\U[1] [13]), .A12(\U[1] [12]), .A11(\U[1] [11]), 
            .A10(\U[1] [10]), .A9(\U[1] [9]), .A8(\U[1] [8]), .A7(\U[1] [7]), 
            .A6(\U[1] [6]), .A5(\U[1] [5]), .A4(\U[1] [4]), .A3(\U[1] [3]), 
            .A2(\U[1] [2]), .A1(\U[1] [1]), .A0(\U[1] [0]), .B17(\x[1] [31]), 
            .B16(\x[1] [31]), .B15(\x[1] [31]), .B14(\x[1] [31]), .B13(\x[1] [31]), 
            .B12(\x[1] [30]), .B11(\x[1] [29]), .B10(\x[1] [28]), .B9(\x[1] [27]), 
            .B8(\x[1] [26]), .B7(\x[1] [25]), .B6(\x[1] [24]), .B5(\x[1] [23]), 
            .B4(\x[1] [22]), .B3(\x[1] [21]), .B2(\x[1] [20]), .B1(\x[1] [19]), 
            .B0(\x[1] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n20401), 
            .ROA16(n20400), .ROA15(n20399), .ROA14(n20398), .ROA13(n20397), 
            .ROA12(n20396), .ROA11(n20395), .ROA10(n20394), .ROA9(n20393), 
            .ROA8(n20392), .ROA7(n20391), .ROA6(n20390), .ROA5(n20389), 
            .ROA4(n20388), .ROA3(n20387), .ROA2(n20386), .ROA1(n20385), 
            .ROA0(n20384), .ROB17(n20419), .ROB16(n20418), .ROB15(n20417), 
            .ROB14(n20416), .ROB13(n20415), .ROB12(n20414), .ROB11(n20413), 
            .ROB10(n20412), .ROB9(n20411), .ROB8(n20410), .ROB7(n20409), 
            .ROB6(n20408), .ROB5(n20407), .ROB4(n20406), .ROB3(n20405), 
            .ROB2(n20404), .ROB1(n20403), .ROB0(n20402), .P35(n20456), 
            .P34(n20455), .P33(n20454), .P32(n20453), .P31(n20452), 
            .P30(n20451), .P29(n20450), .P28(n20449), .P27(n20448), 
            .P26(n20447), .P25(n20446), .P24(n20445), .P23(n20444), 
            .P22(n20443), .P21(n20442), .P20(n20441), .P19(n20440), 
            .P18(n20439), .P17(n20438), .P16(n20437), .P15(n20436), 
            .P14(n20435), .P13(n20434), .P12(n20433), .P11(n20432), 
            .P10(n20431), .P9(n20430), .P8(n20429), .P7(n20428), .P6(n20427), 
            .P5(n20426), .P4(n20425), .P3(n20424), .P2(n20423), .P1(n20422), 
            .P0(n20421), .SIGNEDP(n20420));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(104[16:35])
    defparam lat_mult_26.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_26.REG_INPUTA_CE = "CE0";
    defparam lat_mult_26.REG_INPUTA_RST = "RST0";
    defparam lat_mult_26.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_26.REG_INPUTB_CE = "CE0";
    defparam lat_mult_26.REG_INPUTB_RST = "RST0";
    defparam lat_mult_26.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_26.REG_INPUTC_CE = "CE0";
    defparam lat_mult_26.REG_INPUTC_RST = "RST0";
    defparam lat_mult_26.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_26.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_26.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_26.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_26.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_26.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_26.CLK0_DIV = "ENABLED";
    defparam lat_mult_26.CLK1_DIV = "ENABLED";
    defparam lat_mult_26.CLK2_DIV = "ENABLED";
    defparam lat_mult_26.CLK3_DIV = "ENABLED";
    defparam lat_mult_26.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_26.GSR = "ENABLED";
    defparam lat_mult_26.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_26.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_26.MULT_BYPASS = "DISABLED";
    defparam lat_mult_26.RESETMODE = "SYNC";
    MULT18X18D lat_mult_27 (.A17(\U[1] [31]), .A16(\U[1] [31]), .A15(\U[1] [31]), 
            .A14(\U[1] [31]), .A13(\U[1] [31]), .A12(\U[1] [30]), .A11(\U[1] [29]), 
            .A10(\U[1] [28]), .A9(\U[1] [27]), .A8(\U[1] [26]), .A7(\U[1] [25]), 
            .A6(\U[1] [24]), .A5(\U[1] [23]), .A4(\U[1] [22]), .A3(\U[1] [21]), 
            .A2(\U[1] [20]), .A1(\U[1] [19]), .A0(\U[1] [18]), .B17(\x[1] [31]), 
            .B16(\x[1] [31]), .B15(\x[1] [31]), .B14(\x[1] [31]), .B13(\x[1] [31]), 
            .B12(\x[1] [30]), .B11(\x[1] [29]), .B10(\x[1] [28]), .B9(\x[1] [27]), 
            .B8(\x[1] [26]), .B7(\x[1] [25]), .B6(\x[1] [24]), .B5(\x[1] [23]), 
            .B4(\x[1] [22]), .B3(\x[1] [21]), .B2(\x[1] [20]), .B1(\x[1] [19]), 
            .B0(\x[1] [18]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n20474), 
            .ROA16(n20473), .ROA15(n20472), .ROA14(n20471), .ROA13(n20470), 
            .ROA12(n20469), .ROA11(n20468), .ROA10(n20467), .ROA9(n20466), 
            .ROA8(n20465), .ROA7(n20464), .ROA6(n20463), .ROA5(n20462), 
            .ROA4(n20461), .ROA3(n20460), .ROA2(n20459), .ROA1(n20458), 
            .ROA0(n20457), .ROB17(n20492), .ROB16(n20491), .ROB15(n20490), 
            .ROB14(n20489), .ROB13(n20488), .ROB12(n20487), .ROB11(n20486), 
            .ROB10(n20485), .ROB9(n20484), .ROB8(n20483), .ROB7(n20482), 
            .ROB6(n20481), .ROB5(n20480), .ROB4(n20479), .ROB3(n20478), 
            .ROB2(n20477), .ROB1(n20476), .ROB0(n20475), .P35(n20529), 
            .P34(n20528), .P33(n20527), .P32(n20526), .P31(n20525), 
            .P30(n20524), .P29(n20523), .P28(n20522), .P27(n20521), 
            .P26(n20520), .P25(n20519), .P24(n20518), .P23(n20517), 
            .P22(n20516), .P21(n20515), .P20(n20514), .P19(n20513), 
            .P18(n20512), .P17(n20511), .P16(n20510), .P15(n20509), 
            .P14(n20508), .P13(n20507), .P12(n20506), .P11(n20505), 
            .P10(n20504), .P9(n20503), .P8(n20502), .P7(n20501), .P6(n20500), 
            .P5(n20499), .P4(n20498), .P3(n20497), .P2(n20496), .P1(n20495), 
            .P0(n20494), .SIGNEDP(n20493));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(104[16:35])
    defparam lat_mult_27.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_27.REG_INPUTA_CE = "CE0";
    defparam lat_mult_27.REG_INPUTA_RST = "RST0";
    defparam lat_mult_27.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_27.REG_INPUTB_CE = "CE0";
    defparam lat_mult_27.REG_INPUTB_RST = "RST0";
    defparam lat_mult_27.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_27.REG_INPUTC_CE = "CE0";
    defparam lat_mult_27.REG_INPUTC_RST = "RST0";
    defparam lat_mult_27.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_27.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_27.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_27.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_27.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_27.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_27.CLK0_DIV = "ENABLED";
    defparam lat_mult_27.CLK1_DIV = "ENABLED";
    defparam lat_mult_27.CLK2_DIV = "ENABLED";
    defparam lat_mult_27.CLK3_DIV = "ENABLED";
    defparam lat_mult_27.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_27.GSR = "ENABLED";
    defparam lat_mult_27.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_27.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_27.MULT_BYPASS = "DISABLED";
    defparam lat_mult_27.RESETMODE = "SYNC";
    ALU54B lat_alu_28 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n20274), .SIGNEDIB(n20347), .SIGNEDCIN(GND_net), 
           .A35(n20273), .A34(n20272), .A33(n20271), .A32(n20270), .A31(n20269), 
           .A30(n20268), .A29(n20267), .A28(n20266), .A27(n20265), .A26(n20264), 
           .A25(n20263), .A24(n20262), .A23(n20261), .A22(n20260), .A21(n20259), 
           .A20(n20258), .A19(n20257), .A18(n20256), .A17(n20255), .A16(n20254), 
           .A15(n20253), .A14(n20252), .A13(n20251), .A12(n20250), .A11(n20249), 
           .A10(n20248), .A9(n20247), .A8(n20246), .A7(n20245), .A6(n20244), 
           .A5(n20243), .A4(n20242), .A3(n20241), .A2(n20240), .A1(n20239), 
           .A0(n20238), .B35(n20346), .B34(n20345), .B33(n20344), .B32(n20343), 
           .B31(n20342), .B30(n20341), .B29(n20340), .B28(n20339), .B27(n20338), 
           .B26(n20337), .B25(n20336), .B24(n20335), .B23(n20334), .B22(n20333), 
           .B21(n20332), .B20(n20331), .B19(n20330), .B18(n20329), .B17(n20328), 
           .B16(n20327), .B15(n20326), .B14(n20325), .B13(n20324), .B12(n20323), 
           .B11(n20322), .B10(n20321), .B9(n20320), .B8(n20319), .B7(n20318), 
           .B6(n20317), .B5(n20316), .B4(n20315), .B3(n20314), .B2(n20313), 
           .B1(n20312), .B0(n20311), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n20310), .MA34(n20309), .MA33(n20308), .MA32(n20307), 
           .MA31(n20306), .MA30(n20305), .MA29(n20304), .MA28(n20303), 
           .MA27(n20302), .MA26(n20301), .MA25(n20300), .MA24(n20299), 
           .MA23(n20298), .MA22(n20297), .MA21(n20296), .MA20(n20295), 
           .MA19(n20294), .MA18(n20293), .MA17(n20292), .MA16(n20291), 
           .MA15(n20290), .MA14(n20289), .MA13(n20288), .MA12(n20287), 
           .MA11(n20286), .MA10(n20285), .MA9(n20284), .MA8(n20283), 
           .MA7(n20282), .MA6(n20281), .MA5(n20280), .MA4(n20279), .MA3(n20278), 
           .MA2(n20277), .MA1(n20276), .MA0(n20275), .MB35(n20383), 
           .MB34(n20382), .MB33(n20381), .MB32(n20380), .MB31(n20379), 
           .MB30(n20378), .MB29(n20377), .MB28(n20376), .MB27(n20375), 
           .MB26(n20374), .MB25(n20373), .MB24(n20372), .MB23(n20371), 
           .MB22(n20370), .MB21(n20369), .MB20(n20368), .MB19(n20367), 
           .MB18(n20366), .MB17(n20365), .MB16(n20364), .MB15(n20363), 
           .MB14(n20362), .MB13(n20361), .MB12(n20360), .MB11(n20359), 
           .MB10(n20358), .MB9(n20357), .MB8(n20356), .MB7(n20355), 
           .MB6(n20354), .MB5(n20353), .MB4(n20352), .MB3(n20351), .MB2(n20350), 
           .MB1(n20349), .MB0(n20348), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n20565), 
           .R52(n20564), .R51(n20563), .R50(n20562), .R49(n20561), .R48(n20560), 
           .R47(n20559), .R46(n20558), .R45(n20557), .R44(n20556), .R43(n20555), 
           .R42(n20554), .R41(n20553), .R40(n20552), .R39(n20551), .R38(n20550), 
           .R37(n20549), .R36(n20548), .R35(n20547), .R34(n20546), .R33(n20545), 
           .R32(n20544), .R31(n20543), .R30(n20542), .R29(n20541), .R28(n20540), 
           .R27(n20539), .R26(n20538), .R25(n20537), .R24(n20536), .R23(n20535), 
           .R22(n20534), .R21(n20533), .R20(n20532), .R19(n20531), .R18(n20530), 
           .R17(n177_adj_71), .R16(n178_adj_70), .R15(n179_adj_69), .R14(n180_adj_68), 
           .R13(n181_adj_67), .R12(n182_adj_66), .R11(n183_adj_65), .R10(n184_adj_64), 
           .R9(n185_adj_63), .R8(n186_adj_62), .R7(n187_adj_61), .R6(n188_adj_60), 
           .R5(n189_adj_59), .R4(n190_adj_58), .R3(n191_adj_57), .R2(n192_adj_56), 
           .R1(n193_adj_55), .R0(n194_adj_54), .SIGNEDR(n20566));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(104[16:35])
    defparam lat_alu_28.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_28.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_28.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_28.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_28.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_28.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_28.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_28.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_28.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_28.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_28.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_28.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_28.REG_FLAG_CLK = "NONE";
    defparam lat_alu_28.REG_FLAG_CE = "CE0";
    defparam lat_alu_28.REG_FLAG_RST = "RST0";
    defparam lat_alu_28.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_28.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_28.MASK01 = "0x00000000000000";
    defparam lat_alu_28.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_28.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_28.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_28.CLK0_DIV = "ENABLED";
    defparam lat_alu_28.CLK1_DIV = "ENABLED";
    defparam lat_alu_28.CLK2_DIV = "ENABLED";
    defparam lat_alu_28.CLK3_DIV = "ENABLED";
    defparam lat_alu_28.MCPAT = "0x00000000000000";
    defparam lat_alu_28.MASKPAT = "0x00000000000000";
    defparam lat_alu_28.RNDPAT = "0x00000000000000";
    defparam lat_alu_28.GSR = "ENABLED";
    defparam lat_alu_28.RESETMODE = "SYNC";
    defparam lat_alu_28.MULT9_MODE = "DISABLED";
    defparam lat_alu_28.LEGACY = "DISABLED";
    ALU54B lat_alu_29 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n20420), .SIGNEDIB(n20493), .SIGNEDCIN(n20566), .A35(n20419), 
           .A34(n20418), .A33(n20417), .A32(n20416), .A31(n20415), .A30(n20414), 
           .A29(n20413), .A28(n20412), .A27(n20411), .A26(n20410), .A25(n20409), 
           .A24(n20408), .A23(n20407), .A22(n20406), .A21(n20405), .A20(n20404), 
           .A19(n20403), .A18(n20402), .A17(n20401), .A16(n20400), .A15(n20399), 
           .A14(n20398), .A13(n20397), .A12(n20396), .A11(n20395), .A10(n20394), 
           .A9(n20393), .A8(n20392), .A7(n20391), .A6(n20390), .A5(n20389), 
           .A4(n20388), .A3(n20387), .A2(n20386), .A1(n20385), .A0(n20384), 
           .B35(n20492), .B34(n20491), .B33(n20490), .B32(n20489), .B31(n20488), 
           .B30(n20487), .B29(n20486), .B28(n20485), .B27(n20484), .B26(n20483), 
           .B25(n20482), .B24(n20481), .B23(n20480), .B22(n20479), .B21(n20478), 
           .B20(n20477), .B19(n20476), .B18(n20475), .B17(n20474), .B16(n20473), 
           .B15(n20472), .B14(n20471), .B13(n20470), .B12(n20469), .B11(n20468), 
           .B10(n20467), .B9(n20466), .B8(n20465), .B7(n20464), .B6(n20463), 
           .B5(n20462), .B4(n20461), .B3(n20460), .B2(n20459), .B1(n20458), 
           .B0(n20457), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n20456), .MA34(n20455), .MA33(n20454), .MA32(n20453), 
           .MA31(n20452), .MA30(n20451), .MA29(n20450), .MA28(n20449), 
           .MA27(n20448), .MA26(n20447), .MA25(n20446), .MA24(n20445), 
           .MA23(n20444), .MA22(n20443), .MA21(n20442), .MA20(n20441), 
           .MA19(n20440), .MA18(n20439), .MA17(n20438), .MA16(n20437), 
           .MA15(n20436), .MA14(n20435), .MA13(n20434), .MA12(n20433), 
           .MA11(n20432), .MA10(n20431), .MA9(n20430), .MA8(n20429), 
           .MA7(n20428), .MA6(n20427), .MA5(n20426), .MA4(n20425), .MA3(n20424), 
           .MA2(n20423), .MA1(n20422), .MA0(n20421), .MB35(n20529), 
           .MB34(n20528), .MB33(n20527), .MB32(n20526), .MB31(n20525), 
           .MB30(n20524), .MB29(n20523), .MB28(n20522), .MB27(n20521), 
           .MB26(n20520), .MB25(n20519), .MB24(n20518), .MB23(n20517), 
           .MB22(n20516), .MB21(n20515), .MB20(n20514), .MB19(n20513), 
           .MB18(n20512), .MB17(n20511), .MB16(n20510), .MB15(n20509), 
           .MB14(n20508), .MB13(n20507), .MB12(n20506), .MB11(n20505), 
           .MB10(n20504), .MB9(n20503), .MB8(n20502), .MB7(n20501), 
           .MB6(n20500), .MB5(n20499), .MB4(n20498), .MB3(n20497), .MB2(n20496), 
           .MB1(n20495), .MB0(n20494), .CIN53(n20565), .CIN52(n20564), 
           .CIN51(n20563), .CIN50(n20562), .CIN49(n20561), .CIN48(n20560), 
           .CIN47(n20559), .CIN46(n20558), .CIN45(n20557), .CIN44(n20556), 
           .CIN43(n20555), .CIN42(n20554), .CIN41(n20553), .CIN40(n20552), 
           .CIN39(n20551), .CIN38(n20550), .CIN37(n20549), .CIN36(n20548), 
           .CIN35(n20547), .CIN34(n20546), .CIN33(n20545), .CIN32(n20544), 
           .CIN31(n20543), .CIN30(n20542), .CIN29(n20541), .CIN28(n20540), 
           .CIN27(n20539), .CIN26(n20538), .CIN25(n20537), .CIN24(n20536), 
           .CIN23(n20535), .CIN22(n20534), .CIN21(n20533), .CIN20(n20532), 
           .CIN19(n20531), .CIN18(n20530), .CIN17(n177_adj_71), .CIN16(n178_adj_70), 
           .CIN15(n179_adj_69), .CIN14(n180_adj_68), .CIN13(n181_adj_67), 
           .CIN12(n182_adj_66), .CIN11(n183_adj_65), .CIN10(n184_adj_64), 
           .CIN9(n185_adj_63), .CIN8(n186_adj_62), .CIN7(n187_adj_61), 
           .CIN6(n188_adj_60), .CIN5(n189_adj_59), .CIN4(n190_adj_58), 
           .CIN3(n191_adj_57), .CIN2(n192_adj_56), .CIN1(n193_adj_55), 
           .CIN0(n194_adj_54), .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), 
           .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), 
           .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), 
           .R13(n163_adj_85), .R12(n164_adj_84), .R11(n165_adj_83), .R10(n166_adj_82), 
           .R9(n167_adj_81), .R8(n168_adj_80), .R7(n169_adj_79), .R6(n170_adj_78), 
           .R5(n171_adj_77), .R4(n172_adj_76), .R3(n173_adj_75), .R2(n174_adj_74), 
           .R1(n175_adj_73), .R0(n176_adj_72));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(104[16:35])
    defparam lat_alu_29.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_29.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_29.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_29.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_29.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_29.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_29.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_29.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_29.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_29.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_29.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_29.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_29.REG_FLAG_CLK = "NONE";
    defparam lat_alu_29.REG_FLAG_CE = "CE0";
    defparam lat_alu_29.REG_FLAG_RST = "RST0";
    defparam lat_alu_29.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_29.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_29.MASK01 = "0x00000000000000";
    defparam lat_alu_29.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_29.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_29.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_29.CLK0_DIV = "ENABLED";
    defparam lat_alu_29.CLK1_DIV = "ENABLED";
    defparam lat_alu_29.CLK2_DIV = "ENABLED";
    defparam lat_alu_29.CLK3_DIV = "ENABLED";
    defparam lat_alu_29.MCPAT = "0x00000000000000";
    defparam lat_alu_29.MASKPAT = "0x00000000000000";
    defparam lat_alu_29.RNDPAT = "0x00000000000000";
    defparam lat_alu_29.GSR = "ENABLED";
    defparam lat_alu_29.RESETMODE = "SYNC";
    defparam lat_alu_29.MULT9_MODE = "DISABLED";
    defparam lat_alu_29.LEGACY = "DISABLED";
    LUT4 i1_2_lut_rep_1101 (.A(n105), .B(n104_adj_216), .Z(n42800)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1101.init = 16'heeee;
    FD1S3IX done_4064 (.D(done_N_1928), .CK(clk_c), .CD(rst_c), .Q(done_c));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam done_4064.GSR = "ENABLED";
    MULT18X18D lat_mult_0 (.A17(\U[2] [31]), .A16(\U[2] [31]), .A15(\U[2] [31]), 
            .A14(\U[2] [31]), .A13(\U[2] [31]), .A12(\U[2] [30]), .A11(\U[2] [29]), 
            .A10(\U[2] [28]), .A9(\U[2] [27]), .A8(\U[2] [26]), .A7(\U[2] [25]), 
            .A6(\U[2] [24]), .A5(\U[2] [23]), .A4(\U[2] [22]), .A3(\U[2] [21]), 
            .A2(\U[2] [20]), .A1(\U[2] [19]), .A0(\U[2] [18]), .B17(\x[2] [17]), 
            .B16(\x[2] [16]), .B15(\x[2] [15]), .B14(\x[2] [14]), .B13(\x[2] [13]), 
            .B12(\x[2] [12]), .B11(\x[2] [11]), .B10(\x[2] [10]), .B9(\x[2] [9]), 
            .B8(\x[2] [8]), .B7(\x[2] [7]), .B6(\x[2] [6]), .B5(\x[2] [5]), 
            .B4(\x[2] [4]), .B3(\x[2] [3]), .B2(\x[2] [2]), .B1(\x[2] [1]), 
            .B0(\x[2] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18523), 
            .ROA16(n18522), .ROA15(n18521), .ROA14(n18520), .ROA13(n18519), 
            .ROA12(n18518), .ROA11(n18517), .ROA10(n18516), .ROA9(n18515), 
            .ROA8(n18514), .ROA7(n18513), .ROA6(n18512), .ROA5(n18511), 
            .ROA4(n18510), .ROA3(n18509), .ROA2(n18508), .ROA1(n18507), 
            .ROA0(n18506), .ROB17(n18541), .ROB16(n18540), .ROB15(n18539), 
            .ROB14(n18538), .ROB13(n18537), .ROB12(n18536), .ROB11(n18535), 
            .ROB10(n18534), .ROB9(n18533), .ROB8(n18532), .ROB7(n18531), 
            .ROB6(n18530), .ROB5(n18529), .ROB4(n18528), .ROB3(n18527), 
            .ROB2(n18526), .ROB1(n18525), .ROB0(n18524), .P35(n18578), 
            .P34(n18577), .P33(n18576), .P32(n18575), .P31(n18574), 
            .P30(n18573), .P29(n18572), .P28(n18571), .P27(n18570), 
            .P26(n18569), .P25(n18568), .P24(n18567), .P23(n18566), 
            .P22(n18565), .P21(n18564), .P20(n18563), .P19(n18562), 
            .P18(n18561), .P17(n18560), .P16(n18559), .P15(n18558), 
            .P14(n18557), .P13(n18556), .P12(n18555), .P11(n18554), 
            .P10(n18553), .P9(n18552), .P8(n18551), .P7(n18550), .P6(n18549), 
            .P5(n18548), .P4(n18547), .P3(n18546), .P2(n18545), .P1(n18544), 
            .P0(n18543), .SIGNEDP(n18542));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[16:35])
    defparam lat_mult_0.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTA_CE = "CE0";
    defparam lat_mult_0.REG_INPUTA_RST = "RST0";
    defparam lat_mult_0.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTB_CE = "CE0";
    defparam lat_mult_0.REG_INPUTB_RST = "RST0";
    defparam lat_mult_0.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTC_CE = "CE0";
    defparam lat_mult_0.REG_INPUTC_RST = "RST0";
    defparam lat_mult_0.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_0.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_0.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_0.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_0.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_0.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_0.CLK0_DIV = "ENABLED";
    defparam lat_mult_0.CLK1_DIV = "ENABLED";
    defparam lat_mult_0.CLK2_DIV = "ENABLED";
    defparam lat_mult_0.CLK3_DIV = "ENABLED";
    defparam lat_mult_0.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_0.GSR = "ENABLED";
    defparam lat_mult_0.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_0.MULT_BYPASS = "DISABLED";
    defparam lat_mult_0.RESETMODE = "SYNC";
    MULT18X18D mult_3996_mult_2 (.A17(\U[2] [17]), .A16(\U[2] [16]), .A15(\U[2] [15]), 
            .A14(\U[2] [14]), .A13(\U[2] [13]), .A12(\U[2] [12]), .A11(\U[2] [11]), 
            .A10(\U[2] [10]), .A9(\U[2] [9]), .A8(\U[2] [8]), .A7(\U[2] [7]), 
            .A6(\U[2] [6]), .A5(\U[2] [5]), .A4(\U[2] [4]), .A3(\U[2] [3]), 
            .A2(\U[2] [2]), .A1(\U[2] [1]), .A0(\U[2] [0]), .B17(\x[2] [17]), 
            .B16(\x[2] [16]), .B15(\x[2] [15]), .B14(\x[2] [14]), .B13(\x[2] [13]), 
            .B12(\x[2] [12]), .B11(\x[2] [11]), .B10(\x[2] [10]), .B9(\x[2] [9]), 
            .B8(\x[2] [8]), .B7(\x[2] [7]), .B6(\x[2] [6]), .B5(\x[2] [5]), 
            .B4(\x[2] [4]), .B3(\x[2] [3]), .B2(\x[2] [2]), .B1(\x[2] [1]), 
            .B0(\x[2] [0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18450), 
            .ROA16(n18449), .ROA15(n18448), .ROA14(n18447), .ROA13(n18446), 
            .ROA12(n18445), .ROA11(n18444), .ROA10(n18443), .ROA9(n18442), 
            .ROA8(n18441), .ROA7(n18440), .ROA6(n18439), .ROA5(n18438), 
            .ROA4(n18437), .ROA3(n18436), .ROA2(n18435), .ROA1(n18434), 
            .ROA0(n18433), .ROB17(n18468), .ROB16(n18467), .ROB15(n18466), 
            .ROB14(n18465), .ROB13(n18464), .ROB12(n18463), .ROB11(n18462), 
            .ROB10(n18461), .ROB9(n18460), .ROB8(n18459), .ROB7(n18458), 
            .ROB6(n18457), .ROB5(n18456), .ROB4(n18455), .ROB3(n18454), 
            .ROB2(n18453), .ROB1(n18452), .ROB0(n18451), .P35(n18505), 
            .P34(n18504), .P33(n18503), .P32(n18502), .P31(n18501), 
            .P30(n18500), .P29(n18499), .P28(n18498), .P27(n18497), 
            .P26(n18496), .P25(n18495), .P24(n18494), .P23(n18493), 
            .P22(n18492), .P21(n18491), .P20(n18490), .P19(n18489), 
            .P18(n18488), .P17(n18487), .P16(n18486), .P15(n18485), 
            .P14(n18484), .P13(n18483), .P12(n18482), .P11(n18481), 
            .P10(n18480), .P9(n18479), .P8(n18478), .P7(n18477), .P6(n18476), 
            .P5(n18475), .P4(n18474), .P3(n18473), .P2(n18472), .P1(n18471), 
            .P0(n18470), .SIGNEDP(n18469));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[16:35])
    defparam mult_3996_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_3996_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_3996_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_3996_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_3996_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_3996_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_3996_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_3996_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_3996_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_3996_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_3996_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_3996_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_3996_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_3996_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_3996_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_3996_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_3996_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_3996_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_3996_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_3996_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_3996_mult_2.GSR = "ENABLED";
    defparam mult_3996_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_3996_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_3996_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_3996_mult_2.RESETMODE = "SYNC";
    FD1P3AX U_15___i512 (.D(\U[0] [31]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i512.GSR = "ENABLED";
    IB U_in_pad_165 (.I(U_in[165]), .O(U_in_c_165));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_166 (.I(U_in[166]), .O(U_in_c_166));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_167 (.I(U_in[167]), .O(U_in_c_167));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_168 (.I(U_in[168]), .O(U_in_c_168));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_169 (.I(U_in[169]), .O(U_in_c_169));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_170 (.I(U_in[170]), .O(U_in_c_170));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_171 (.I(U_in[171]), .O(U_in_c_171));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_172 (.I(U_in[172]), .O(U_in_c_172));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_173 (.I(U_in[173]), .O(U_in_c_173));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_174 (.I(U_in[174]), .O(U_in_c_174));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_175 (.I(U_in[175]), .O(U_in_c_175));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_176 (.I(U_in[176]), .O(U_in_c_176));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_177 (.I(U_in[177]), .O(U_in_c_177));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_178 (.I(U_in[178]), .O(U_in_c_178));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_179 (.I(U_in[179]), .O(U_in_c_179));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_180 (.I(U_in[180]), .O(U_in_c_180));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_181 (.I(U_in[181]), .O(U_in_c_181));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_182 (.I(U_in[182]), .O(U_in_c_182));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_183 (.I(U_in[183]), .O(U_in_c_183));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_184 (.I(U_in[184]), .O(U_in_c_184));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_185 (.I(U_in[185]), .O(U_in_c_185));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_186 (.I(U_in[186]), .O(U_in_c_186));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_187 (.I(U_in[187]), .O(U_in_c_187));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_188 (.I(U_in[188]), .O(U_in_c_188));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_189 (.I(U_in[189]), .O(U_in_c_189));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_190 (.I(U_in[190]), .O(U_in_c_190));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_191 (.I(U_in[191]), .O(U_in_c_191));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_192 (.I(U_in[192]), .O(U_in_c_192));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    LUT4 div_4016_LessThan_2598_i29_2_lut_rep_901 (.A(n3970), .B(n126), 
         .Z(n42600)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i29_2_lut_rep_901.init = 16'h6666;
    LUT4 i1_2_lut_rep_1094_3_lut_4_lut (.A(n105), .B(n104_adj_216), .C(n102), 
         .D(n103_adj_215), .Z(n42793)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1094_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23239_2_lut_3_lut_4_lut (.A(n3970), .B(n126), .C(n127_adj_231), 
         .D(n3971), .Z(n38499)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23239_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2598_i26_3_lut_3_lut (.A(n3970), .B(n126), .C(n127_adj_231), 
         .Z(n26_adj_498)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2598_i23_2_lut_rep_902 (.A(n3973), .B(n129), 
         .Z(n42601)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i23_2_lut_rep_902.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i22_3_lut_3_lut (.A(n3973), .B(n129), .C(n130_adj_233), 
         .Z(n22_adj_495)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i3320_4_lut (.A(n37218), .B(n22284), .C(n42786), .D(n64_adj_269), 
         .Z(n5503)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3320_4_lut.init = 16'hc0c5;
    LUT4 i25640_4_lut_4_lut (.A(n42605), .B(n38467), .C(n52_adj_487), 
         .D(n28_adj_473), .Z(n54_adj_488)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25640_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i23219_4_lut_4_lut (.A(n42605), .B(n38452), .C(n42604), .D(n42602), 
         .Z(n38479)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23219_4_lut_4_lut.init = 16'h00fb;
    LUT4 i1_4_lut_adj_28 (.A(n37210), .B(n35955), .C(n37212), .D(n42805), 
         .Z(n37218)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_28.init = 16'hfffe;
    FD1P3IX x_3___i122 (.D(n5500), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i122.GSR = "ENABLED";
    LUT4 div_4016_LessThan_2153_i64_4_lut (.A(n50_adj_391), .B(n62_adj_398), 
         .C(n42662), .D(n38041), .Z(n64_adj_399)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i64_4_lut.init = 16'hcacc;
    LUT4 i22781_4_lut (.A(n42663), .B(n42665), .C(n42664), .D(n38020), 
         .Z(n38041)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22781_4_lut.init = 16'h0100;
    IB U_in_pad_193 (.I(U_in[193]), .O(U_in_c_193));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_194 (.I(U_in[194]), .O(U_in_c_194));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_195 (.I(U_in[195]), .O(U_in_c_195));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_196 (.I(U_in[196]), .O(U_in_c_196));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_197 (.I(U_in[197]), .O(U_in_c_197));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_198 (.I(U_in[198]), .O(U_in_c_198));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_199 (.I(U_in[199]), .O(U_in_c_199));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_200 (.I(U_in[200]), .O(U_in_c_200));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_201 (.I(U_in[201]), .O(U_in_c_201));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_202 (.I(U_in[202]), .O(U_in_c_202));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_203 (.I(U_in[203]), .O(U_in_c_203));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_204 (.I(U_in[204]), .O(U_in_c_204));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_205 (.I(U_in[205]), .O(U_in_c_205));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_206 (.I(U_in[206]), .O(U_in_c_206));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_207 (.I(U_in[207]), .O(U_in_c_207));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_208 (.I(U_in[208]), .O(U_in_c_208));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_209 (.I(U_in[209]), .O(U_in_c_209));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_210 (.I(U_in[210]), .O(U_in_c_210));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_211 (.I(U_in[211]), .O(U_in_c_211));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_212 (.I(U_in[212]), .O(U_in_c_212));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_213 (.I(U_in[213]), .O(U_in_c_213));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_214 (.I(U_in[214]), .O(U_in_c_214));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_215 (.I(U_in[215]), .O(U_in_c_215));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_216 (.I(U_in[216]), .O(U_in_c_216));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_217 (.I(U_in[217]), .O(U_in_c_217));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_218 (.I(U_in[218]), .O(U_in_c_218));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_219 (.I(U_in[219]), .O(U_in_c_219));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    LUT4 i22760_4_lut (.A(n42666), .B(n53_adj_393), .C(n42667), .D(n38003), 
         .Z(n38020)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22760_4_lut.init = 16'h1011;
    LUT4 i22743_4_lut (.A(n42668), .B(n42670), .C(n42669), .D(n37988), 
         .Z(n38003)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22743_4_lut.init = 16'h0100;
    L6MUX21 div_4016_LessThan_2337_i62 (.D0(n50_adj_437), .D1(n60_adj_442), 
            .SD(n38255), .Z(n62_adj_443));
    PFUMX div_4016_LessThan_2337_i60 (.BLUT(n52_adj_438), .ALUT(n58_adj_441), 
          .C0(n38257), .Z(n60_adj_442));
    LUT4 i22728_4_lut (.A(n42672), .B(n42671), .C(n42673), .D(n37975), 
         .Z(n37988)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22728_4_lut.init = 16'h5455;
    LUT4 i22715_4_lut (.A(n37_adj_384), .B(n35), .C(n42674), .D(n31_adj_380), 
         .Z(n37975)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22715_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_2153_i31_2_lut (.A(n3309), .B(n130_adj_233), 
         .Z(n31_adj_380)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i31_2_lut.init = 16'h6666;
    IB U_in_pad_220 (.I(U_in[220]), .O(U_in_c_220));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_221 (.I(U_in[221]), .O(U_in_c_221));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_222 (.I(U_in[222]), .O(U_in_c_222));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_223 (.I(U_in[223]), .O(U_in_c_223));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_224 (.I(U_in[224]), .O(U_in_c_224));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_225 (.I(U_in[225]), .O(U_in_c_225));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_226 (.I(U_in[226]), .O(U_in_c_226));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_227 (.I(U_in[227]), .O(U_in_c_227));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_228 (.I(U_in[228]), .O(U_in_c_228));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_229 (.I(U_in[229]), .O(U_in_c_229));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_230 (.I(U_in[230]), .O(U_in_c_230));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_231 (.I(U_in[231]), .O(U_in_c_231));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_232 (.I(U_in[232]), .O(U_in_c_232));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_233 (.I(U_in[233]), .O(U_in_c_233));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_234 (.I(U_in[234]), .O(U_in_c_234));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_235 (.I(U_in[235]), .O(U_in_c_235));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_236 (.I(U_in[236]), .O(U_in_c_236));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_237 (.I(U_in[237]), .O(U_in_c_237));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_238 (.I(U_in[238]), .O(U_in_c_238));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_239 (.I(U_in[239]), .O(U_in_c_239));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_240 (.I(U_in[240]), .O(U_in_c_240));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_241 (.I(U_in[241]), .O(U_in_c_241));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_242 (.I(U_in[242]), .O(U_in_c_242));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_243 (.I(U_in[243]), .O(U_in_c_243));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_244 (.I(U_in[244]), .O(U_in_c_244));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_245 (.I(U_in[245]), .O(U_in_c_245));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C div_4016_unary_minus_4_add_3_33 (.A0(n5460), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32854), .S0(n68_adj_194));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_33.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_33.INIT1 = 16'h0000;
    defparam div_4016_unary_minus_4_add_3_33.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_33.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_31 (.A0(n5462), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5461), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32853), .COUT(n32854), .S0(n70_adj_195), .S1(n69));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_31.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_31.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_31.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_31.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_29 (.A0(n5464), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5463), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32852), .COUT(n32853), .S0(n72), .S1(n71_adj_196));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_29.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_29.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_29.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_29.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_27 (.A0(n5466), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5465), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32851), .COUT(n32852), .S0(n74_adj_198), .S1(n73_adj_197));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_27.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_27.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_27.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_27.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_25 (.A0(n5468), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5467), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32850), .COUT(n32851), .S0(n76_adj_199), .S1(n75));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_25.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_25.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_25.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_25.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_23 (.A0(n5470), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5469), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32849), .COUT(n32850), .S0(n78), .S1(n77_adj_200));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_23.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_23.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_23.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_23.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_29 (.A(n36784), .B(n42813), .C(n42798), .D(n42796), 
         .Z(n30917)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_29.init = 16'hfffe;
    LUT4 div_4016_LessThan_2513_i61_2_lut_rep_903 (.A(n3828), .B(n111), 
         .Z(n42602)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i61_2_lut_rep_903.init = 16'h6666;
    LUT4 i1_4_lut_adj_30 (.A(n37206), .B(n42819), .C(n120), .D(n122_adj_228), 
         .Z(n37212)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_30.init = 16'hfffe;
    LUT4 div_4016_LessThan_2153_i37_2_lut (.A(n3306), .B(n127_adj_231), 
         .Z(n37_adj_384)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i37_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2513_i34_3_lut_3_lut (.A(n3828), .B(n111), .C(n123), 
         .Z(n34_adj_477)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_adj_31 (.A(n105), .B(n104_adj_216), .C(n42802), 
         .D(n42803), .Z(n36784)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_31.init = 16'hfffe;
    LUT4 div_4016_LessThan_2153_i35_2_lut (.A(n3307), .B(n128_adj_232), 
         .Z(n35)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i35_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i36_3_lut_3_lut (.A(n4656), .B(n113_adj_222), 
         .C(n114), .Z(n36_adj_689)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i36_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_2337_i50 (.BLUT(n26_adj_422), .ALUT(n48_adj_435), 
          .C0(n38223), .Z(n50_adj_437));
    LUT4 div_4016_LessThan_2153_i53_2_lut (.A(n3298), .B(n119_adj_226), 
         .Z(n53_adj_393)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i53_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_1102 (.A(n104_adj_216), .B(n107_adj_218), .Z(n42801)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1102.init = 16'heeee;
    IB U_in_pad_246 (.I(U_in[246]), .O(U_in_c_246));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_247 (.I(U_in[247]), .O(U_in_c_247));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_248 (.I(U_in[248]), .O(U_in_c_248));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_249 (.I(U_in[249]), .O(U_in_c_249));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_250 (.I(U_in[250]), .O(U_in_c_250));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_251 (.I(U_in[251]), .O(U_in_c_251));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_252 (.I(U_in[252]), .O(U_in_c_252));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_253 (.I(U_in[253]), .O(U_in_c_253));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_254 (.I(U_in[254]), .O(U_in_c_254));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_255 (.I(U_in[255]), .O(U_in_c_255));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_256 (.I(U_in[256]), .O(U_in_c_256));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_257 (.I(U_in[257]), .O(U_in_c_257));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_258 (.I(U_in[258]), .O(U_in_c_258));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_259 (.I(U_in[259]), .O(U_in_c_259));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_260 (.I(U_in[260]), .O(U_in_c_260));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_261 (.I(U_in[261]), .O(U_in_c_261));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_262 (.I(U_in[262]), .O(U_in_c_262));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_263 (.I(U_in[263]), .O(U_in_c_263));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_264 (.I(U_in[264]), .O(U_in_c_264));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_265 (.I(U_in[265]), .O(U_in_c_265));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_266 (.I(U_in[266]), .O(U_in_c_266));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_267 (.I(U_in[267]), .O(U_in_c_267));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_268 (.I(U_in[268]), .O(U_in_c_268));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_269 (.I(U_in[269]), .O(U_in_c_269));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_270 (.I(U_in[270]), .O(U_in_c_270));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C div_4016_unary_minus_4_add_3_21 (.A0(n5472), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5471), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32848), .COUT(n32849), .S0(n80_adj_202), .S1(n79_adj_201));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_21.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_21.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_21.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_21.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_19 (.A0(n5474), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5473), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32847), .COUT(n32848), .S0(n82_adj_203), .S1(n81));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_19.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_19.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_19.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_19.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_17 (.A0(n5476), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5475), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32846), .COUT(n32847), .S0(n84), .S1(n83_adj_204));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_17.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_17.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_17.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_17.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_15 (.A0(n5478), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5477), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32845), .COUT(n32846), .S0(n86_adj_206), .S1(n85_adj_205));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_15.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_15.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_15.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_15.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_13 (.A0(n5480), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5479), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32844), .COUT(n32845), .S0(n88_adj_207), .S1(n87));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_13.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_13.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_13.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_13.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_11 (.A0(n5482), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5481), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32843), .COUT(n32844), .S0(n90), .S1(n89_adj_208));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_11.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_11.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_11.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_11.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_9 (.A0(n5484), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5483), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32842), .COUT(n32843), .S0(n92_adj_210), .S1(n91_adj_209));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_9.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_9.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_9.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_9.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_3066_i45_2_lut_rep_775 (.A(n4655), .B(n112_adj_221), 
         .Z(n42474)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i45_2_lut_rep_775.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i64_4_lut (.A(n58_adj_266), .B(n62_adj_268), 
         .C(n42750), .D(n37508), .Z(n64_adj_269)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i64_4_lut.init = 16'hcacc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_32 (.A(n104_adj_216), .B(n107_adj_218), 
         .C(n105), .D(n102), .Z(n37298)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_32.init = 16'hfffe;
    LUT4 i22248_4_lut (.A(n42752), .B(n42751), .C(n42753), .D(n37495), 
         .Z(n37508)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22248_4_lut.init = 16'h5455;
    PFUMX div_4016_LessThan_2337_i46 (.BLUT(n38_adj_430), .ALUT(n44_adj_433), 
          .C0(n38199), .Z(n46_adj_434));
    LUT4 i1_3_lut_4_lut_adj_33 (.A(n104_adj_216), .B(n107_adj_218), .C(n105), 
         .D(n103_adj_215), .Z(n37146)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_33.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i38_3_lut_3_lut (.A(n4655), .B(n112_adj_221), 
         .C(n36_adj_689), .Z(n38_adj_690)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22235_4_lut (.A(n55_adj_264), .B(n42755), .C(n42754), .D(n49), 
         .Z(n37495)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22235_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_1226_i49_2_lut (.A(n1923), .B(n130_adj_233), 
         .Z(n49)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i49_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_1553_i42_4_lut (.A(n132), .B(n131_adj_234), .C(n2413), 
         .D(n875), .Z(n42)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i42_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2513_i63_2_lut_rep_904 (.A(n3827), .B(n110_adj_220), 
         .Z(n42603)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i63_2_lut_rep_904.init = 16'h6666;
    LUT4 div_4016_LessThan_1226_i55_2_lut (.A(n1920), .B(n127_adj_231), 
         .Z(n55_adj_264)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1226_i55_2_lut.init = 16'h6666;
    IB U_in_pad_271 (.I(U_in[271]), .O(U_in_c_271));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_272 (.I(U_in[272]), .O(U_in_c_272));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_273 (.I(U_in[273]), .O(U_in_c_273));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_274 (.I(U_in[274]), .O(U_in_c_274));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_275 (.I(U_in[275]), .O(U_in_c_275));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_276 (.I(U_in[276]), .O(U_in_c_276));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_277 (.I(U_in[277]), .O(U_in_c_277));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_278 (.I(U_in[278]), .O(U_in_c_278));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_279 (.I(U_in[279]), .O(U_in_c_279));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_280 (.I(U_in[280]), .O(U_in_c_280));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_281 (.I(U_in[281]), .O(U_in_c_281));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_282 (.I(U_in[282]), .O(U_in_c_282));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_283 (.I(U_in[283]), .O(U_in_c_283));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_284 (.I(U_in[284]), .O(U_in_c_284));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_285 (.I(U_in[285]), .O(U_in_c_285));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_286 (.I(U_in[286]), .O(U_in_c_286));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_287 (.I(U_in[287]), .O(U_in_c_287));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_288 (.I(U_in[288]), .O(U_in_c_288));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_289 (.I(U_in[289]), .O(U_in_c_289));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_290 (.I(U_in[290]), .O(U_in_c_290));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_291 (.I(U_in[291]), .O(U_in_c_291));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_292 (.I(U_in[292]), .O(U_in_c_292));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_293 (.I(U_in[293]), .O(U_in_c_293));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_294 (.I(U_in[294]), .O(U_in_c_294));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C div_4016_unary_minus_4_add_3_7 (.A0(n5486), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5485), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32841), .COUT(n32842), .S0(n94_adj_211), .S1(n93));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_7.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_7.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_7.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_7.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_5 (.A0(n5488), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5487), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32840), .COUT(n32841), .S0(n96), .S1(n95_adj_212));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_5.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_5.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_5.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_5.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_3 (.A0(n5490), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5489), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32839), .COUT(n32840), .S0(n98_adj_214), .S1(n97_adj_213));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_3.INIT0 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_3.INIT1 = 16'h5550;
    defparam div_4016_unary_minus_4_add_3_3.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_3.INJECT1_1 = "NO";
    CCU2C div_4016_unary_minus_4_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5491), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32839), .S1(n99));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_unary_minus_4_add_3_1.INIT0 = 16'h0000;
    defparam div_4016_unary_minus_4_add_3_1.INIT1 = 16'haaaf;
    defparam div_4016_unary_minus_4_add_3_1.INJECT1_0 = "NO";
    defparam div_4016_unary_minus_4_add_3_1.INJECT1_1 = "NO";
    CCU2C add_16626_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32838), 
          .S0(n16519));
    defparam add_16626_cout.INIT0 = 16'h0000;
    defparam add_16626_cout.INIT1 = 16'h0000;
    defparam add_16626_cout.INJECT1_0 = "NO";
    defparam add_16626_cout.INJECT1_1 = "NO";
    CCU2C add_16626_31 (.A0(i[30]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[31]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32837), 
          .COUT(n32838));
    defparam add_16626_31.INIT0 = 16'h5555;
    defparam add_16626_31.INIT1 = 16'h555f;
    defparam add_16626_31.INJECT1_0 = "NO";
    defparam add_16626_31.INJECT1_1 = "NO";
    CCU2C add_16626_29 (.A0(i[28]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[29]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32836), 
          .COUT(n32837));
    defparam add_16626_29.INIT0 = 16'h5555;
    defparam add_16626_29.INIT1 = 16'h5555;
    defparam add_16626_29.INJECT1_0 = "NO";
    defparam add_16626_29.INJECT1_1 = "NO";
    CCU2C add_16626_27 (.A0(i[26]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[27]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32835), 
          .COUT(n32836));
    defparam add_16626_27.INIT0 = 16'h5555;
    defparam add_16626_27.INIT1 = 16'h5555;
    defparam add_16626_27.INJECT1_0 = "NO";
    defparam add_16626_27.INJECT1_1 = "NO";
    LUT4 i25806_4_lut (.A(n42474), .B(n42473), .C(n42475), .D(n39440), 
         .Z(n39458)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25806_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2513_i60_3_lut_3_lut (.A(n3827), .B(n110_adj_220), 
         .C(n42_adj_481), .Z(n60_adj_491)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i3328_4_lut (.A(n37092), .B(n22292), .C(n42786), .D(n64_adj_378), 
         .Z(n5511)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3328_4_lut.init = 16'hc0c5;
    LUT4 i1_4_lut_adj_34 (.A(n37298), .B(n37082), .C(n37144), .D(n42795), 
         .Z(n37092)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_34.init = 16'hfffe;
    LUT4 div_4016_LessThan_2513_i57_2_lut_rep_905 (.A(n3830), .B(n113_adj_222), 
         .Z(n42604)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i57_2_lut_rep_905.init = 16'h6666;
    L6MUX21 div_4016_LessThan_2246_i62 (.D0(n52_adj_415), .D1(n60_adj_419), 
            .SD(n38148), .Z(n62_adj_420));
    LUT4 div_4016_mux_3_i3_3_lut (.A(n5354), .B(n31_adj_191), .C(n5325), 
         .Z(n892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i3_3_lut.init = 16'hcaca;
    LUT4 mux_4010_i3_4_lut (.A(n157), .B(n36646), .C(n15805), .D(i[1]), 
         .Z(n5354)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i3_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_35 (.A(i[0]), .B(\y[3] [2]), .Z(n36646)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_35.init = 16'h8888;
    IB U_in_pad_295 (.I(U_in[295]), .O(U_in_c_295));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_296 (.I(U_in[296]), .O(U_in_c_296));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_297 (.I(U_in[297]), .O(U_in_c_297));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_298 (.I(U_in[298]), .O(U_in_c_298));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_299 (.I(U_in[299]), .O(U_in_c_299));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_300 (.I(U_in[300]), .O(U_in_c_300));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_301 (.I(U_in[301]), .O(U_in_c_301));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_302 (.I(U_in[302]), .O(U_in_c_302));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_303 (.I(U_in[303]), .O(U_in_c_303));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_304 (.I(U_in[304]), .O(U_in_c_304));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_305 (.I(U_in[305]), .O(U_in_c_305));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_306 (.I(U_in[306]), .O(U_in_c_306));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_307 (.I(U_in[307]), .O(U_in_c_307));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_308 (.I(U_in[308]), .O(U_in_c_308));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_309 (.I(U_in[309]), .O(U_in_c_309));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_310 (.I(U_in[310]), .O(U_in_c_310));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_311 (.I(U_in[311]), .O(U_in_c_311));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_312 (.I(U_in[312]), .O(U_in_c_312));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_313 (.I(U_in[313]), .O(U_in_c_313));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_314 (.I(U_in[314]), .O(U_in_c_314));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_315 (.I(U_in[315]), .O(U_in_c_315));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_316 (.I(U_in[316]), .O(U_in_c_316));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_317 (.I(U_in[317]), .O(U_in_c_317));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_16626_25 (.A0(i[24]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[25]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32834), 
          .COUT(n32835));
    defparam add_16626_25.INIT0 = 16'h5555;
    defparam add_16626_25.INIT1 = 16'h5555;
    defparam add_16626_25.INJECT1_0 = "NO";
    defparam add_16626_25.INJECT1_1 = "NO";
    CCU2C add_16626_23 (.A0(i[22]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[23]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32833), 
          .COUT(n32834));
    defparam add_16626_23.INIT0 = 16'h5555;
    defparam add_16626_23.INIT1 = 16'h5555;
    defparam add_16626_23.INJECT1_0 = "NO";
    defparam add_16626_23.INJECT1_1 = "NO";
    CCU2C add_16626_21 (.A0(i[20]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[21]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32832), 
          .COUT(n32833));
    defparam add_16626_21.INIT0 = 16'h5555;
    defparam add_16626_21.INIT1 = 16'h5555;
    defparam add_16626_21.INJECT1_0 = "NO";
    defparam add_16626_21.INJECT1_1 = "NO";
    CCU2C add_16626_19 (.A0(i[18]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[19]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32831), 
          .COUT(n32832));
    defparam add_16626_19.INIT0 = 16'h5555;
    defparam add_16626_19.INIT1 = 16'h5555;
    defparam add_16626_19.INJECT1_0 = "NO";
    defparam add_16626_19.INJECT1_1 = "NO";
    CCU2C add_16626_17 (.A0(i[16]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32830), 
          .COUT(n32831));
    defparam add_16626_17.INIT0 = 16'h5555;
    defparam add_16626_17.INIT1 = 16'h5555;
    defparam add_16626_17.INJECT1_0 = "NO";
    defparam add_16626_17.INJECT1_1 = "NO";
    CCU2C add_16626_15 (.A0(i[14]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[15]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32829), 
          .COUT(n32830));
    defparam add_16626_15.INIT0 = 16'h5555;
    defparam add_16626_15.INIT1 = 16'h5555;
    defparam add_16626_15.INJECT1_0 = "NO";
    defparam add_16626_15.INJECT1_1 = "NO";
    CCU2C add_16626_13 (.A0(i[12]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[13]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32828), 
          .COUT(n32829));
    defparam add_16626_13.INIT0 = 16'h5555;
    defparam add_16626_13.INIT1 = 16'h5555;
    defparam add_16626_13.INJECT1_0 = "NO";
    defparam add_16626_13.INJECT1_1 = "NO";
    CCU2C add_16626_11 (.A0(i[10]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[11]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32827), 
          .COUT(n32828));
    defparam add_16626_11.INIT0 = 16'h5555;
    defparam add_16626_11.INIT1 = 16'h5555;
    defparam add_16626_11.INJECT1_0 = "NO";
    defparam add_16626_11.INJECT1_1 = "NO";
    CCU2C add_16626_9 (.A0(i[8]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[9]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32826), 
          .COUT(n32827));
    defparam add_16626_9.INIT0 = 16'h5555;
    defparam add_16626_9.INIT1 = 16'h5555;
    defparam add_16626_9.INJECT1_0 = "NO";
    defparam add_16626_9.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_3066_i41_2_lut_rep_776 (.A(n4657), .B(n114), 
         .Z(n42475)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i41_2_lut_rep_776.init = 16'h6666;
    LUT4 i24191_2_lut_3_lut_4_lut (.A(n4657), .B(n114), .C(n113_adj_222), 
         .D(n4656), .Z(n39451)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24191_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2513_i50_3_lut_3_lut (.A(n3830), .B(n113_adj_222), 
         .C(n114), .Z(n50_adj_486)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i50_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_2246_i60 (.BLUT(n54_adj_416), .ALUT(n58_adj_418), 
          .C0(n38150), .Z(n60_adj_419));
    LUT4 div_4016_LessThan_2513_i59_2_lut_rep_906 (.A(n3829), .B(n112_adj_221), 
         .Z(n42605)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i59_2_lut_rep_906.init = 16'h6666;
    IB U_in_pad_318 (.I(U_in[318]), .O(U_in_c_318));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_319 (.I(U_in[319]), .O(U_in_c_319));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_320 (.I(U_in[320]), .O(U_in_c_320));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_321 (.I(U_in[321]), .O(U_in_c_321));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_322 (.I(U_in[322]), .O(U_in_c_322));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_323 (.I(U_in[323]), .O(U_in_c_323));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_324 (.I(U_in[324]), .O(U_in_c_324));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_325 (.I(U_in[325]), .O(U_in_c_325));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_326 (.I(U_in[326]), .O(U_in_c_326));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_327 (.I(U_in[327]), .O(U_in_c_327));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_328 (.I(U_in[328]), .O(U_in_c_328));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_329 (.I(U_in[329]), .O(U_in_c_329));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_330 (.I(U_in[330]), .O(U_in_c_330));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_331 (.I(U_in[331]), .O(U_in_c_331));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_332 (.I(U_in[332]), .O(U_in_c_332));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_333 (.I(U_in[333]), .O(U_in_c_333));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_334 (.I(U_in[334]), .O(U_in_c_334));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_335 (.I(U_in[335]), .O(U_in_c_335));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_336 (.I(U_in[336]), .O(U_in_c_336));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_337 (.I(U_in[337]), .O(U_in_c_337));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_338 (.I(U_in[338]), .O(U_in_c_338));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_339 (.I(U_in[339]), .O(U_in_c_339));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_16626_7 (.A0(i[6]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[7]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32825), 
          .COUT(n32826));
    defparam add_16626_7.INIT0 = 16'h5555;
    defparam add_16626_7.INIT1 = 16'h5555;
    defparam add_16626_7.INJECT1_0 = "NO";
    defparam add_16626_7.INJECT1_1 = "NO";
    CCU2C add_16626_5 (.A0(i[4]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[5]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32824), 
          .COUT(n32825));
    defparam add_16626_5.INIT0 = 16'h5555;
    defparam add_16626_5.INIT1 = 16'h5555;
    defparam add_16626_5.INJECT1_0 = "NO";
    defparam add_16626_5.INJECT1_1 = "NO";
    CCU2C add_16626_3 (.A0(i[2]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[3]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32823), 
          .COUT(n32824));
    defparam add_16626_3.INIT0 = 16'h5555;
    defparam add_16626_3.INIT1 = 16'h5555;
    defparam add_16626_3.INJECT1_0 = "NO";
    defparam add_16626_3.INJECT1_1 = "NO";
    CCU2C add_16626_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[1]), .B1(i[0]), .C1(GND_net), .D1(VCC_net), .COUT(n32823));
    defparam add_16626_1.INIT0 = 16'h0000;
    defparam add_16626_1.INIT1 = 16'h6665;
    defparam add_16626_1.INJECT1_0 = "NO";
    defparam add_16626_1.INJECT1_1 = "NO";
    CCU2C add_17618_33 (.A0(n3), .B0(n163_adj_12), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32822), 
          .S0(n32354));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_33.INIT0 = 16'h666a;
    defparam add_17618_33.INIT1 = 16'h0000;
    defparam add_17618_33.INJECT1_0 = "NO";
    defparam add_17618_33.INJECT1_1 = "NO";
    CCU2C add_17618_31 (.A0(n5), .B0(n165), .C0(GND_net), .D0(VCC_net), 
          .A1(n4), .B1(n164), .C1(GND_net), .D1(VCC_net), .CIN(n32821), 
          .COUT(n32822), .S0(n32356), .S1(n32355));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_31.INIT0 = 16'h666a;
    defparam add_17618_31.INIT1 = 16'h666a;
    defparam add_17618_31.INJECT1_0 = "NO";
    defparam add_17618_31.INJECT1_1 = "NO";
    CCU2C add_17618_29 (.A0(n7), .B0(n167), .C0(GND_net), .D0(VCC_net), 
          .A1(n6), .B1(n166), .C1(GND_net), .D1(VCC_net), .CIN(n32820), 
          .COUT(n32821), .S0(n32358), .S1(n32357));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_29.INIT0 = 16'h666a;
    defparam add_17618_29.INIT1 = 16'h666a;
    defparam add_17618_29.INJECT1_0 = "NO";
    defparam add_17618_29.INJECT1_1 = "NO";
    CCU2C add_17618_27 (.A0(n9), .B0(n169), .C0(GND_net), .D0(VCC_net), 
          .A1(n8), .B1(n168_adj_10), .C1(GND_net), .D1(VCC_net), .CIN(n32819), 
          .COUT(n32820), .S0(n32360), .S1(n32359));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_27.INIT0 = 16'h666a;
    defparam add_17618_27.INIT1 = 16'h666a;
    defparam add_17618_27.INJECT1_0 = "NO";
    defparam add_17618_27.INJECT1_1 = "NO";
    CCU2C add_17618_25 (.A0(n11), .B0(n171), .C0(GND_net), .D0(VCC_net), 
          .A1(n10), .B1(n170), .C1(GND_net), .D1(VCC_net), .CIN(n32818), 
          .COUT(n32819), .S0(n32362), .S1(n32361));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_25.INIT0 = 16'h666a;
    defparam add_17618_25.INIT1 = 16'h666a;
    defparam add_17618_25.INJECT1_0 = "NO";
    defparam add_17618_25.INJECT1_1 = "NO";
    CCU2C add_17618_23 (.A0(n13), .B0(n173_adj_9), .C0(GND_net), .D0(VCC_net), 
          .A1(n12), .B1(n172_adj_8), .C1(GND_net), .D1(VCC_net), .CIN(n32817), 
          .COUT(n32818), .S0(n32364), .S1(n32363));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_23.INIT0 = 16'h666a;
    defparam add_17618_23.INIT1 = 16'h666a;
    defparam add_17618_23.INJECT1_0 = "NO";
    defparam add_17618_23.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_2513_i52_3_lut_3_lut (.A(n3829), .B(n112_adj_221), 
         .C(n50_adj_486), .Z(n52_adj_487)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i3327_4_lut (.A(n64_adj_360), .B(n22291), .C(n42786), 
         .D(n30911), .Z(n5510)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3327_4_lut.init = 16'hc0c5;
    LUT4 i1_4_lut_adj_36 (.A(n36606), .B(n42806), .C(n42816), .D(n42796), 
         .Z(n30911)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_36.init = 16'hfffe;
    LUT4 div_4016_i3326_4_lut (.A(n37122), .B(n22290), .C(n42786), .D(n64_adj_343), 
         .Z(n5509)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3326_4_lut.init = 16'hc0c5;
    LUT4 i1_4_lut_adj_37 (.A(n37120), .B(n37176), .C(n42812), .D(n36720), 
         .Z(n37122)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_37.init = 16'hfffe;
    LUT4 i1_2_lut_adj_38 (.A(n115_adj_223), .B(n116_adj_224), .Z(n36720)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_38.init = 16'heeee;
    PFUMX div_4016_LessThan_2246_i52 (.BLUT(n28_adj_400), .ALUT(n50_adj_413), 
          .C0(n38125), .Z(n52_adj_415));
    IB U_in_pad_340 (.I(U_in[340]), .O(U_in_c_340));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_341 (.I(U_in[341]), .O(U_in_c_341));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_342 (.I(U_in[342]), .O(U_in_c_342));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_343 (.I(U_in[343]), .O(U_in_c_343));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_344 (.I(U_in[344]), .O(U_in_c_344));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_345 (.I(U_in[345]), .O(U_in_c_345));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_346 (.I(U_in[346]), .O(U_in_c_346));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_347 (.I(U_in[347]), .O(U_in_c_347));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_348 (.I(U_in[348]), .O(U_in_c_348));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_349 (.I(U_in[349]), .O(U_in_c_349));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_350 (.I(U_in[350]), .O(U_in_c_350));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_351 (.I(U_in[351]), .O(U_in_c_351));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_352 (.I(U_in[352]), .O(U_in_c_352));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_353 (.I(U_in[353]), .O(U_in_c_353));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_354 (.I(U_in[354]), .O(U_in_c_354));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_355 (.I(U_in[355]), .O(U_in_c_355));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_356 (.I(U_in[356]), .O(U_in_c_356));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_357 (.I(U_in[357]), .O(U_in_c_357));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_358 (.I(U_in[358]), .O(U_in_c_358));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_359 (.I(U_in[359]), .O(U_in_c_359));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_360 (.I(U_in[360]), .O(U_in_c_360));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_17618_21 (.A0(n15), .B0(n175), .C0(GND_net), .D0(VCC_net), 
          .A1(n14), .B1(n174), .C1(GND_net), .D1(VCC_net), .CIN(n32816), 
          .COUT(n32817), .S0(n32366), .S1(n32365));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_21.INIT0 = 16'h666a;
    defparam add_17618_21.INIT1 = 16'h666a;
    defparam add_17618_21.INJECT1_0 = "NO";
    defparam add_17618_21.INJECT1_1 = "NO";
    CCU2C add_17618_19 (.A0(n17), .B0(n177), .C0(GND_net), .D0(VCC_net), 
          .A1(n16), .B1(n176), .C1(GND_net), .D1(VCC_net), .CIN(n32815), 
          .COUT(n32816), .S0(n32368), .S1(n32367));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_19.INIT0 = 16'h666a;
    defparam add_17618_19.INIT1 = 16'h666a;
    defparam add_17618_19.INJECT1_0 = "NO";
    defparam add_17618_19.INJECT1_1 = "NO";
    CCU2C add_17618_17 (.A0(n19), .B0(n179), .C0(GND_net), .D0(VCC_net), 
          .A1(n18), .B1(n178_adj_5), .C1(GND_net), .D1(VCC_net), .CIN(n32814), 
          .COUT(n32815), .S0(n32370), .S1(n32369));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_17.INIT0 = 16'h666a;
    defparam add_17618_17.INIT1 = 16'h666a;
    defparam add_17618_17.INJECT1_0 = "NO";
    defparam add_17618_17.INJECT1_1 = "NO";
    CCU2C add_17618_15 (.A0(n21), .B0(n181), .C0(GND_net), .D0(VCC_net), 
          .A1(n20), .B1(n180), .C1(GND_net), .D1(VCC_net), .CIN(n32813), 
          .COUT(n32814), .S0(n32372), .S1(n32371));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_15.INIT0 = 16'h666a;
    defparam add_17618_15.INIT1 = 16'h666a;
    defparam add_17618_15.INJECT1_0 = "NO";
    defparam add_17618_15.INJECT1_1 = "NO";
    CCU2C add_17618_13 (.A0(n23), .B0(n183_adj_3), .C0(GND_net), .D0(VCC_net), 
          .A1(n22), .B1(n182), .C1(GND_net), .D1(VCC_net), .CIN(n32812), 
          .COUT(n32813), .S0(n32374), .S1(n32373));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_13.INIT0 = 16'h666a;
    defparam add_17618_13.INIT1 = 16'h666a;
    defparam add_17618_13.INJECT1_0 = "NO";
    defparam add_17618_13.INJECT1_1 = "NO";
    CCU2C add_17618_11 (.A0(n25), .B0(n185), .C0(GND_net), .D0(VCC_net), 
          .A1(n24), .B1(n184), .C1(GND_net), .D1(VCC_net), .CIN(n32811), 
          .COUT(n32812), .S0(n32376), .S1(n32375));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_11.INIT0 = 16'h666a;
    defparam add_17618_11.INIT1 = 16'h666a;
    defparam add_17618_11.INJECT1_0 = "NO";
    defparam add_17618_11.INJECT1_1 = "NO";
    CCU2C add_17618_9 (.A0(n27), .B0(n187), .C0(GND_net), .D0(VCC_net), 
          .A1(n26), .B1(n186), .C1(GND_net), .D1(VCC_net), .CIN(n32810), 
          .COUT(n32811), .S0(n32378), .S1(n32377));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_9.INIT0 = 16'h666a;
    defparam add_17618_9.INIT1 = 16'h666a;
    defparam add_17618_9.INJECT1_0 = "NO";
    defparam add_17618_9.INJECT1_1 = "NO";
    CCU2C add_17618_7 (.A0(n29), .B0(n189), .C0(GND_net), .D0(VCC_net), 
          .A1(n28), .B1(n188_adj_2), .C1(GND_net), .D1(VCC_net), .CIN(n32809), 
          .COUT(n32810), .S0(n32380), .S1(n32379));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_7.INIT0 = 16'h666a;
    defparam add_17618_7.INIT1 = 16'h666a;
    defparam add_17618_7.INJECT1_0 = "NO";
    defparam add_17618_7.INJECT1_1 = "NO";
    CCU2C add_17618_5 (.A0(n31), .B0(n191), .C0(GND_net), .D0(VCC_net), 
          .A1(n30), .B1(n190), .C1(GND_net), .D1(VCC_net), .CIN(n32808), 
          .COUT(n32809), .S0(n32382), .S1(n32381));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_5.INIT0 = 16'h666a;
    defparam add_17618_5.INIT1 = 16'h666a;
    defparam add_17618_5.INJECT1_0 = "NO";
    defparam add_17618_5.INJECT1_1 = "NO";
    CCU2C add_17618_3 (.A0(n33), .B0(n193_adj_1), .C0(GND_net), .D0(VCC_net), 
          .A1(n32), .B1(n192), .C1(GND_net), .D1(VCC_net), .CIN(n32807), 
          .COUT(n32808), .S0(n32384), .S1(n32383));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_3.INIT0 = 16'h666a;
    defparam add_17618_3.INIT1 = 16'h666a;
    defparam add_17618_3.INJECT1_0 = "NO";
    defparam add_17618_3.INJECT1_1 = "NO";
    CCU2C add_17618_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n194_adj_114), .B1(n194_adj_54), .C1(n194), .D1(VCC_net), 
          .COUT(n32807), .S1(n32385));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam add_17618_1.INIT0 = 16'h0000;
    defparam add_17618_1.INIT1 = 16'h9696;
    defparam add_17618_1.INJECT1_0 = "NO";
    defparam add_17618_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1104 (.A(n107_adj_218), .B(n106_adj_217), .Z(n42803)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1104.init = 16'heeee;
    LUT4 div_4016_LessThan_3066_i39_2_lut_rep_777 (.A(n4658), .B(n115_adj_223), 
         .Z(n42476)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i39_2_lut_rep_777.init = 16'h6666;
    PFUMX div_4016_LessThan_2246_i48 (.BLUT(n40_adj_408), .ALUT(n46_adj_411), 
          .C0(n38101), .Z(n48_adj_412));
    LUT4 div_4016_LessThan_3066_i34_3_lut_3_lut (.A(n4658), .B(n115_adj_223), 
         .C(n16_adj_676), .Z(n34_adj_688)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_4_lut_adj_39 (.A(n42799), .B(n42795), .C(n104_adj_216), .D(n106_adj_217), 
         .Z(n35955)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_39.init = 16'hfffe;
    LUT4 div_4016_LessThan_2513_i55_2_lut_rep_907 (.A(n3831), .B(n114), 
         .Z(n42606)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i55_2_lut_rep_907.init = 16'h6666;
    LUT4 i24180_3_lut_4_lut (.A(n4658), .B(n115_adj_223), .C(n19_adj_678), 
         .D(n42478), .Z(n39440)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24180_3_lut_4_lut.init = 16'h0009;
    LUT4 i1_2_lut_rep_1098_3_lut_4_lut (.A(n107_adj_218), .B(n106_adj_217), 
         .C(n104_adj_216), .D(n105), .Z(n42797)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1098_3_lut_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i35_2_lut_rep_778 (.A(n4660), .B(n117), 
         .Z(n42477)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i35_2_lut_rep_778.init = 16'h6666;
    IB U_in_pad_361 (.I(U_in[361]), .O(U_in_c_361));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_362 (.I(U_in[362]), .O(U_in_c_362));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_363 (.I(U_in[363]), .O(U_in_c_363));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_364 (.I(U_in[364]), .O(U_in_c_364));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_365 (.I(U_in[365]), .O(U_in_c_365));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_366 (.I(U_in[366]), .O(U_in_c_366));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_367 (.I(U_in[367]), .O(U_in_c_367));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_368 (.I(U_in[368]), .O(U_in_c_368));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_369 (.I(U_in[369]), .O(U_in_c_369));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_370 (.I(U_in[370]), .O(U_in_c_370));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_371 (.I(U_in[371]), .O(U_in_c_371));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_372 (.I(U_in[372]), .O(U_in_c_372));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_373 (.I(U_in[373]), .O(U_in_c_373));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_374 (.I(U_in[374]), .O(U_in_c_374));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_375 (.I(U_in[375]), .O(U_in_c_375));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_376 (.I(U_in[376]), .O(U_in_c_376));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_377 (.I(U_in[377]), .O(U_in_c_377));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_378 (.I(U_in[378]), .O(U_in_c_378));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_379 (.I(U_in[379]), .O(U_in_c_379));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_380 (.I(U_in[380]), .O(U_in_c_380));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7646_33 (.A0(n30962), .B0(n4_adj_235), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32806), 
          .S0(n22275));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_33.INIT0 = 16'heeee;
    defparam add_7646_33.INIT1 = 16'h0000;
    defparam add_7646_33.INJECT1_0 = "NO";
    defparam add_7646_33.INJECT1_1 = "NO";
    CCU2C add_7646_31 (.A0(n42776), .B0(n30965), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_799), .B1(n30962), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32805), .COUT(n32806), .S0(n22277), .S1(n22276));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_31.INIT0 = 16'heeee;
    defparam add_7646_31.INIT1 = 16'heeee;
    defparam add_7646_31.INJECT1_0 = "NO";
    defparam add_7646_31.INJECT1_1 = "NO";
    CCU2C add_7646_29 (.A0(n64), .B0(n30872), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_797), .B1(n30968), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32804), .COUT(n32805), .S0(n22279), .S1(n22278));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_29.INIT0 = 16'heeee;
    defparam add_7646_29.INIT1 = 16'heeee;
    defparam add_7646_29.INJECT1_0 = "NO";
    defparam add_7646_29.INJECT1_1 = "NO";
    CCU2C add_7646_27 (.A0(n64_adj_246), .B0(n30881), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_241), .B1(n30878), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32803), .COUT(n32804), .S0(n22281), .S1(n22280));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_27.INIT0 = 16'heeee;
    defparam add_7646_27.INIT1 = 16'heeee;
    defparam add_7646_27.INJECT1_0 = "NO";
    defparam add_7646_27.INJECT1_1 = "NO";
    CCU2C add_7646_25 (.A0(n64_adj_260), .B0(n30887), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_252), .B1(n30884), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32802), .COUT(n32803), .S0(n22283), .S1(n22282));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_25.INIT0 = 16'heeee;
    defparam add_7646_25.INIT1 = 16'heeee;
    defparam add_7646_25.INJECT1_0 = "NO";
    defparam add_7646_25.INJECT1_1 = "NO";
    CCU2C add_7646_23 (.A0(n64_adj_278), .B0(n30893), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_269), .B1(n30890), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32801), .COUT(n32802), .S0(n22285), .S1(n22284));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_23.INIT0 = 16'heeee;
    defparam add_7646_23.INIT1 = 16'heeee;
    defparam add_7646_23.INJECT1_0 = "NO";
    defparam add_7646_23.INJECT1_1 = "NO";
    CCU2C add_7646_21 (.A0(n64_adj_301), .B0(n42789), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_289), .B1(n30896), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32800), .COUT(n32801), .S0(n22287), .S1(n22286));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_21.INIT0 = 16'heeee;
    defparam add_7646_21.INIT1 = 16'heeee;
    defparam add_7646_21.INJECT1_0 = "NO";
    defparam add_7646_21.INJECT1_1 = "NO";
    CCU2C add_7646_19 (.A0(n64_adj_328), .B0(n30905), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_315), .B1(n30902), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32799), .COUT(n32800), .S0(n22289), .S1(n22288));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_19.INIT0 = 16'heeee;
    defparam add_7646_19.INIT1 = 16'heeee;
    defparam add_7646_19.INJECT1_0 = "NO";
    defparam add_7646_19.INJECT1_1 = "NO";
    CCU2C add_7646_17 (.A0(n64_adj_360), .B0(n30911), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_343), .B1(n30908), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32798), .COUT(n32799), .S0(n22291), .S1(n22290));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_17.INIT0 = 16'heeee;
    defparam add_7646_17.INIT1 = 16'heeee;
    defparam add_7646_17.INJECT1_0 = "NO";
    defparam add_7646_17.INJECT1_1 = "NO";
    CCU2C add_7646_15 (.A0(n64_adj_399), .B0(n30917), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_378), .B1(n30914), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32797), .COUT(n32798), .S0(n22293), .S1(n22292));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_15.INIT0 = 16'heeee;
    defparam add_7646_15.INIT1 = 16'heeee;
    defparam add_7646_15.INJECT1_0 = "NO";
    defparam add_7646_15.INJECT1_1 = "NO";
    CCU2C add_7646_13 (.A0(n64_adj_444), .B0(n30923), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_421), .B1(n30920), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32796), .COUT(n32797), .S0(n22295), .S1(n22294));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_13.INIT0 = 16'heeee;
    defparam add_7646_13.INIT1 = 16'heeee;
    defparam add_7646_13.INJECT1_0 = "NO";
    defparam add_7646_13.INJECT1_1 = "NO";
    CCU2C add_7646_11 (.A0(n64_adj_493), .B0(n30929), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_469), .B1(n30926), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32795), .COUT(n32796), .S0(n22297), .S1(n22296));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_11.INIT0 = 16'heeee;
    defparam add_7646_11.INIT1 = 16'heeee;
    defparam add_7646_11.INJECT1_0 = "NO";
    defparam add_7646_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1105 (.A(n106_adj_217), .B(n109_adj_219), .Z(n42804)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1105.init = 16'heeee;
    LUT4 i23207_2_lut_3_lut_4_lut (.A(n3831), .B(n114), .C(n113_adj_222), 
         .D(n3830), .Z(n38467)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23207_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i1_2_lut_3_lut_4_lut_adj_40 (.A(n106_adj_217), .B(n109_adj_219), 
         .C(n107_adj_218), .D(n104_adj_216), .Z(n36832)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_40.init = 16'hfffe;
    LUT4 i24064_4_lut (.A(n42491), .B(n42490), .C(n42492), .D(n39308), 
         .Z(n39324)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24064_4_lut.init = 16'h1011;
    IB U_in_pad_381 (.I(U_in[381]), .O(U_in_c_381));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_382 (.I(U_in[382]), .O(U_in_c_382));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_383 (.I(U_in[383]), .O(U_in_c_383));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_384 (.I(U_in[384]), .O(U_in_c_384));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_385 (.I(U_in[385]), .O(U_in_c_385));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_386 (.I(U_in[386]), .O(U_in_c_386));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_387 (.I(U_in[387]), .O(U_in_c_387));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_388 (.I(U_in[388]), .O(U_in_c_388));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_389 (.I(U_in[389]), .O(U_in_c_389));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_390 (.I(U_in[390]), .O(U_in_c_390));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_391 (.I(U_in[391]), .O(U_in_c_391));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_392 (.I(U_in[392]), .O(U_in_c_392));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_393 (.I(U_in[393]), .O(U_in_c_393));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_394 (.I(U_in[394]), .O(U_in_c_394));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_395 (.I(U_in[395]), .O(U_in_c_395));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_396 (.I(U_in[396]), .O(U_in_c_396));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_397 (.I(U_in[397]), .O(U_in_c_397));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_398 (.I(U_in[398]), .O(U_in_c_398));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_399 (.I(U_in[399]), .O(U_in_c_399));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7646_9 (.A0(n64_adj_549), .B0(n42790), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_520), .B1(n30932), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32794), .COUT(n32795), .S0(n22299), .S1(n22298));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_9.INIT0 = 16'heeee;
    defparam add_7646_9.INIT1 = 16'heeee;
    defparam add_7646_9.INJECT1_0 = "NO";
    defparam add_7646_9.INJECT1_1 = "NO";
    CCU2C add_7646_7 (.A0(n64_adj_608), .B0(n42794), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_578), .B1(n30938), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32793), .COUT(n32794), .S0(n22301), .S1(n22300));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_7.INIT0 = 16'heeee;
    defparam add_7646_7.INIT1 = 16'heeee;
    defparam add_7646_7.INJECT1_0 = "NO";
    defparam add_7646_7.INJECT1_1 = "NO";
    CCU2C add_7646_5 (.A0(n64_adj_670), .B0(n42792), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_640), .B1(n30944), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32792), .COUT(n32793), .S0(n22303), .S1(n22302));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_5.INIT0 = 16'heeee;
    defparam add_7646_5.INIT1 = 16'heeee;
    defparam add_7646_5.INJECT1_0 = "NO";
    defparam add_7646_5.INJECT1_1 = "NO";
    CCU2C add_7646_3 (.A0(n64_adj_737), .B0(n42796), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_703), .B1(n30950), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32791), .COUT(n32792), .S0(n22305), .S1(n22304));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_3.INIT0 = 16'heeee;
    defparam add_7646_3.INIT1 = 16'heeee;
    defparam add_7646_3.INJECT1_0 = "NO";
    defparam add_7646_3.INJECT1_1 = "NO";
    CCU2C add_7646_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n42440), .B1(n5460), .C1(n68_adj_194), .D1(n62_adj_794), 
          .COUT(n32791), .S1(n22306));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7646_1.INIT0 = 16'h0000;
    defparam add_7646_1.INIT1 = 16'h2abf;
    defparam add_7646_1.INJECT1_0 = "NO";
    defparam add_7646_1.INJECT1_1 = "NO";
    CCU2C add_7645_33 (.A0(n4751), .B0(n102), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32790), 
          .S0(n22241));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_33.INIT0 = 16'h999a;
    defparam add_7645_33.INIT1 = 16'h0000;
    defparam add_7645_33.INJECT1_0 = "NO";
    defparam add_7645_33.INJECT1_1 = "NO";
    CCU2C add_7645_31 (.A0(n4753), .B0(n104_adj_216), .C0(GND_net), .D0(VCC_net), 
          .A1(n4752), .B1(n103_adj_215), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32789), .COUT(n32790), .S0(n22243), .S1(n22242));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_31.INIT0 = 16'h999a;
    defparam add_7645_31.INIT1 = 16'h999a;
    defparam add_7645_31.INJECT1_0 = "NO";
    defparam add_7645_31.INJECT1_1 = "NO";
    CCU2C add_7645_29 (.A0(n4755), .B0(n106_adj_217), .C0(GND_net), .D0(VCC_net), 
          .A1(n4754), .B1(n105), .C1(GND_net), .D1(VCC_net), .CIN(n32788), 
          .COUT(n32789), .S0(n22245), .S1(n22244));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_29.INIT0 = 16'h999a;
    defparam add_7645_29.INIT1 = 16'h999a;
    defparam add_7645_29.INJECT1_0 = "NO";
    defparam add_7645_29.INJECT1_1 = "NO";
    CCU2C add_7645_27 (.A0(n4757), .B0(n108), .C0(GND_net), .D0(VCC_net), 
          .A1(n4756), .B1(n107_adj_218), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32787), .COUT(n32788), .S0(n22247), .S1(n22246));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_27.INIT0 = 16'h999a;
    defparam add_7645_27.INIT1 = 16'h999a;
    defparam add_7645_27.INJECT1_0 = "NO";
    defparam add_7645_27.INJECT1_1 = "NO";
    CCU2C add_7645_25 (.A0(n4759), .B0(n110_adj_220), .C0(GND_net), .D0(VCC_net), 
          .A1(n4758), .B1(n109_adj_219), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32786), .COUT(n32787), .S0(n22249), .S1(n22248));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_25.INIT0 = 16'h999a;
    defparam add_7645_25.INIT1 = 16'h999a;
    defparam add_7645_25.INJECT1_0 = "NO";
    defparam add_7645_25.INJECT1_1 = "NO";
    CCU2C add_7645_23 (.A0(n4761), .B0(n112_adj_221), .C0(GND_net), .D0(VCC_net), 
          .A1(n4760), .B1(n111), .C1(GND_net), .D1(VCC_net), .CIN(n32785), 
          .COUT(n32786), .S0(n22251), .S1(n22250));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_23.INIT0 = 16'h999a;
    defparam add_7645_23.INIT1 = 16'h999a;
    defparam add_7645_23.INJECT1_0 = "NO";
    defparam add_7645_23.INJECT1_1 = "NO";
    CCU2C add_7645_21 (.A0(n4763), .B0(n114), .C0(GND_net), .D0(VCC_net), 
          .A1(n4762), .B1(n113_adj_222), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32784), .COUT(n32785), .S0(n22253), .S1(n22252));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_21.INIT0 = 16'h999a;
    defparam add_7645_21.INIT1 = 16'h999a;
    defparam add_7645_21.INJECT1_0 = "NO";
    defparam add_7645_21.INJECT1_1 = "NO";
    CCU2C add_7645_19 (.A0(n4765), .B0(n116_adj_224), .C0(GND_net), .D0(VCC_net), 
          .A1(n4764), .B1(n115_adj_223), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32783), .COUT(n32784), .S0(n22255), .S1(n22254));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_19.INIT0 = 16'h999a;
    defparam add_7645_19.INIT1 = 16'h999a;
    defparam add_7645_19.INJECT1_0 = "NO";
    defparam add_7645_19.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_3066_i30_3_lut_3_lut (.A(n4660), .B(n117), .C(n18_adj_677), 
         .Z(n30_adj_685)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2513_i53_2_lut_rep_908 (.A(n3832), .B(n115_adj_223), 
         .Z(n42607)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i53_2_lut_rep_908.init = 16'h6666;
    LUT4 div_4016_LessThan_2513_i48_3_lut_3_lut (.A(n3832), .B(n115_adj_223), 
         .C(n30_adj_474), .Z(n48_adj_485)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23196_3_lut_4_lut (.A(n3832), .B(n115_adj_223), .C(n33_adj_476), 
         .D(n42609), .Z(n38456)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23196_3_lut_4_lut.init = 16'h0009;
    L6MUX21 div_4016_LessThan_2153_i62 (.D0(n54_adj_394), .D1(n60_adj_397), 
            .SD(n38050), .Z(n62_adj_398));
    LUT4 div_4016_LessThan_2513_i49_2_lut_rep_909 (.A(n3834), .B(n117), 
         .Z(n42608)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i49_2_lut_rep_909.init = 16'h6666;
    PFUMX div_4016_LessThan_2153_i60 (.BLUT(n56_adj_395), .ALUT(n58_adj_396), 
          .C0(n38054), .Z(n60_adj_397));
    LUT4 i1_3_lut_4_lut_adj_41 (.A(n106_adj_217), .B(n109_adj_219), .C(n107_adj_218), 
         .D(n105), .Z(n37178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_41.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1108 (.A(n108), .B(n111), .Z(n42807)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1108.init = 16'heeee;
    LUT4 div_4016_LessThan_2513_i44_3_lut_3_lut (.A(n3834), .B(n117), .C(n32_adj_475), 
         .Z(n44_adj_482)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(n108), .B(n111), .C(n109_adj_219), 
         .D(n106_adj_217), .Z(n37144)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'hfffe;
    IB U_in_pad_400 (.I(U_in[400]), .O(U_in_c_400));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_401 (.I(U_in[401]), .O(U_in_c_401));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_402 (.I(U_in[402]), .O(U_in_c_402));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_403 (.I(U_in[403]), .O(U_in_c_403));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_404 (.I(U_in[404]), .O(U_in_c_404));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_405 (.I(U_in[405]), .O(U_in_c_405));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_406 (.I(U_in[406]), .O(U_in_c_406));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_407 (.I(U_in[407]), .O(U_in_c_407));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_408 (.I(U_in[408]), .O(U_in_c_408));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_409 (.I(U_in[409]), .O(U_in_c_409));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_410 (.I(U_in[410]), .O(U_in_c_410));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_411 (.I(U_in[411]), .O(U_in_c_411));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_412 (.I(U_in[412]), .O(U_in_c_412));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_413 (.I(U_in[413]), .O(U_in_c_413));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_414 (.I(U_in[414]), .O(U_in_c_414));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_415 (.I(U_in[415]), .O(U_in_c_415));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_416 (.I(U_in[416]), .O(U_in_c_416));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_417 (.I(U_in[417]), .O(U_in_c_417));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7645_17 (.A0(n4767), .B0(n118_adj_225), .C0(GND_net), .D0(VCC_net), 
          .A1(n4766), .B1(n117), .C1(GND_net), .D1(VCC_net), .CIN(n32782), 
          .COUT(n32783), .S0(n22257), .S1(n22256));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_17.INIT0 = 16'h999a;
    defparam add_7645_17.INIT1 = 16'h999a;
    defparam add_7645_17.INJECT1_0 = "NO";
    defparam add_7645_17.INJECT1_1 = "NO";
    CCU2C add_7645_15 (.A0(n4769), .B0(n120), .C0(GND_net), .D0(VCC_net), 
          .A1(n4768), .B1(n119_adj_226), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32781), .COUT(n32782), .S0(n22259), .S1(n22258));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_15.INIT0 = 16'h999a;
    defparam add_7645_15.INIT1 = 16'h999a;
    defparam add_7645_15.INJECT1_0 = "NO";
    defparam add_7645_15.INJECT1_1 = "NO";
    CCU2C add_7645_13 (.A0(n4771), .B0(n122_adj_228), .C0(GND_net), .D0(VCC_net), 
          .A1(n4770), .B1(n121_adj_227), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32780), .COUT(n32781), .S0(n22261), .S1(n22260));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_13.INIT0 = 16'h999a;
    defparam add_7645_13.INIT1 = 16'h999a;
    defparam add_7645_13.INJECT1_0 = "NO";
    defparam add_7645_13.INJECT1_1 = "NO";
    CCU2C add_7645_11 (.A0(n4773), .B0(n124_adj_229), .C0(GND_net), .D0(VCC_net), 
          .A1(n4772), .B1(n123), .C1(GND_net), .D1(VCC_net), .CIN(n32779), 
          .COUT(n32780), .S0(n22263), .S1(n22262));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_11.INIT0 = 16'h999a;
    defparam add_7645_11.INIT1 = 16'h999a;
    defparam add_7645_11.INJECT1_0 = "NO";
    defparam add_7645_11.INJECT1_1 = "NO";
    CCU2C add_7645_9 (.A0(n4775), .B0(n126), .C0(GND_net), .D0(VCC_net), 
          .A1(n4774), .B1(n125_adj_230), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32778), .COUT(n32779), .S0(n22265), .S1(n22264));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_9.INIT0 = 16'h999a;
    defparam add_7645_9.INIT1 = 16'h999a;
    defparam add_7645_9.INJECT1_0 = "NO";
    defparam add_7645_9.INJECT1_1 = "NO";
    CCU2C add_7645_7 (.A0(n4777), .B0(n128_adj_232), .C0(GND_net), .D0(VCC_net), 
          .A1(n4776), .B1(n127_adj_231), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32777), .COUT(n32778), .S0(n22267), .S1(n22266));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_7.INIT0 = 16'h999a;
    defparam add_7645_7.INIT1 = 16'h999a;
    defparam add_7645_7.INJECT1_0 = "NO";
    defparam add_7645_7.INJECT1_1 = "NO";
    CCU2C add_7645_5 (.A0(n4779), .B0(n130_adj_233), .C0(GND_net), .D0(VCC_net), 
          .A1(n4778), .B1(n129), .C1(GND_net), .D1(VCC_net), .CIN(n32776), 
          .COUT(n32777), .S0(n22269), .S1(n22268));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_5.INIT0 = 16'h999a;
    defparam add_7645_5.INIT1 = 16'h999a;
    defparam add_7645_5.INJECT1_0 = "NO";
    defparam add_7645_5.INJECT1_1 = "NO";
    CCU2C add_7645_3 (.A0(n132), .B0(n32_adj_192), .C0(n5325), .D0(n5355), 
          .A1(n4780), .B1(n131_adj_234), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32775), .COUT(n32776), .S0(n22271), .S1(n22270));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_3.INIT0 = 16'h9a95;
    defparam add_7645_3.INIT1 = 16'h999a;
    defparam add_7645_3.INJECT1_0 = "NO";
    defparam add_7645_3.INJECT1_1 = "NO";
    CCU2C add_7645_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n708), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .COUT(n32775));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7645_1.INIT0 = 16'h000F;
    defparam add_7645_1.INIT1 = 16'h555a;
    defparam add_7645_1.INJECT1_0 = "NO";
    defparam add_7645_1.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_32 (.A0(n164_adj_149), .B0(n164_adj_84), 
          .C0(GND_net), .D0(VCC_net), .A1(n163), .B1(n163_adj_85), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32773), .S0(n4), .S1(n3));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_32.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_32.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_32.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_32.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_30 (.A0(n166_adj_147), .B0(n166_adj_82), 
          .C0(GND_net), .D0(VCC_net), .A1(n165_adj_148), .B1(n165_adj_83), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32772), .COUT(n32773), .S0(n6), 
          .S1(n5));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_30.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_30.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_30.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_30.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_28 (.A0(n168), .B0(n168_adj_80), 
          .C0(GND_net), .D0(VCC_net), .A1(n167_adj_146), .B1(n167_adj_81), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32771), .COUT(n32772), .S0(n8), 
          .S1(n7));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_28.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_28.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_28.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_28.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_26 (.A0(n170_adj_142), .B0(n170_adj_78), 
          .C0(GND_net), .D0(VCC_net), .A1(n169_adj_143), .B1(n169_adj_79), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32770), .COUT(n32771), .S0(n10), 
          .S1(n9));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_26.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_26.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_26.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_26.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_24 (.A0(n172_adj_140), .B0(n172_adj_76), 
          .C0(GND_net), .D0(VCC_net), .A1(n171_adj_141), .B1(n171_adj_77), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32769), .COUT(n32770), .S0(n12), 
          .S1(n11));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_24.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_24.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_24.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_24.INJECT1_1 = "NO";
    LUT4 i25793_3_lut_4_lut (.A(n3834), .B(n117), .C(n45_adj_483), .D(n42610), 
         .Z(n38440)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25793_3_lut_4_lut.init = 16'hfff6;
    LUT4 i25812_3_lut_4_lut (.A(n4660), .B(n117), .C(n31_adj_686), .D(n42479), 
         .Z(n39424)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25812_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_3066_i37_2_lut_rep_779 (.A(n4659), .B(n116_adj_224), 
         .Z(n42478)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i37_2_lut_rep_779.init = 16'h6666;
    PFUMX div_4016_LessThan_2153_i54 (.BLUT(n30_adj_379), .ALUT(n52_adj_392), 
          .C0(n38036), .Z(n54_adj_394));
    LUT4 i25791_4_lut (.A(n42605), .B(n42604), .C(n42606), .D(n38447), 
         .Z(n38472)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25791_4_lut.init = 16'hfeff;
    IB U_in_pad_418 (.I(U_in[418]), .O(U_in_c_418));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_419 (.I(U_in[419]), .O(U_in_c_419));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_420 (.I(U_in[420]), .O(U_in_c_420));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_421 (.I(U_in[421]), .O(U_in_c_421));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_422 (.I(U_in[422]), .O(U_in_c_422));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_423 (.I(U_in[423]), .O(U_in_c_423));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_424 (.I(U_in[424]), .O(U_in_c_424));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_425 (.I(U_in[425]), .O(U_in_c_425));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_426 (.I(U_in[426]), .O(U_in_c_426));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_427 (.I(U_in[427]), .O(U_in_c_427));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_428 (.I(U_in[428]), .O(U_in_c_428));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_429 (.I(U_in[429]), .O(U_in_c_429));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_430 (.I(U_in[430]), .O(U_in_c_430));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_431 (.I(U_in[431]), .O(U_in_c_431));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_432 (.I(U_in[432]), .O(U_in_c_432));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_433 (.I(U_in[433]), .O(U_in_c_433));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_434 (.I(U_in[434]), .O(U_in_c_434));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C _add_1_7035_add_4_add_1_add_1_22 (.A0(n174_adj_137), .B0(n174_adj_74), 
          .C0(GND_net), .D0(VCC_net), .A1(n173), .B1(n173_adj_75), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32768), .COUT(n32769), .S0(n14), .S1(n13));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_22.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_22.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_22.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_22.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_20 (.A0(n176_adj_135), .B0(n176_adj_72), 
          .C0(GND_net), .D0(VCC_net), .A1(n175_adj_136), .B1(n175_adj_73), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32767), .COUT(n32768), .S0(n16), 
          .S1(n15));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_20.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_20.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_20.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_20.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_18 (.A0(n178), .B0(n178_adj_70), 
          .C0(GND_net), .D0(VCC_net), .A1(n177_adj_134), .B1(n177_adj_71), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32766), .COUT(n32767), .S0(n18), 
          .S1(n17));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_18.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_18.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_18.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_18.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_16 (.A0(n180_adj_130), .B0(n180_adj_68), 
          .C0(GND_net), .D0(VCC_net), .A1(n179_adj_131), .B1(n179_adj_69), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32765), .COUT(n32766), .S0(n20), 
          .S1(n19));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_16.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_16.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_16.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_16.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_14 (.A0(n182_adj_128), .B0(n182_adj_66), 
          .C0(GND_net), .D0(VCC_net), .A1(n181_adj_129), .B1(n181_adj_67), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32764), .COUT(n32765), .S0(n22), 
          .S1(n21));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_14.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_14.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_14.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_14.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_12 (.A0(n184_adj_125), .B0(n184_adj_64), 
          .C0(GND_net), .D0(VCC_net), .A1(n183), .B1(n183_adj_65), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32763), .COUT(n32764), .S0(n24), .S1(n23));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_12.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_12.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_12.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_12.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_10 (.A0(n186_adj_123), .B0(n186_adj_62), 
          .C0(GND_net), .D0(VCC_net), .A1(n185_adj_124), .B1(n185_adj_63), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32762), .COUT(n32763), .S0(n26), 
          .S1(n25));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_10.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_10.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_10.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_10.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_8 (.A0(n188), .B0(n188_adj_60), 
          .C0(GND_net), .D0(VCC_net), .A1(n187_adj_122), .B1(n187_adj_61), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32761), .COUT(n32762), .S0(n28), 
          .S1(n27));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_8.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_8.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_8.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_8.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_6 (.A0(n190_adj_118), .B0(n190_adj_58), 
          .C0(GND_net), .D0(VCC_net), .A1(n189_adj_119), .B1(n189_adj_59), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32760), .COUT(n32761), .S0(n30), 
          .S1(n29));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_6.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_6.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_6.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_6.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_4 (.A0(n192_adj_116), .B0(n192_adj_56), 
          .C0(GND_net), .D0(VCC_net), .A1(n191_adj_117), .B1(n191_adj_57), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32759), .COUT(n32760), .S0(n32), 
          .S1(n31));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_4.INIT0 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_4.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_4.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_4.INJECT1_1 = "NO";
    CCU2C _add_1_7035_add_4_add_1_add_1_2 (.A0(n194_adj_114), .B0(n194_adj_54), 
          .C0(GND_net), .D0(VCC_net), .A1(n193), .B1(n193_adj_55), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32759), .S1(n33));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(103[10:35])
    defparam _add_1_7035_add_4_add_1_add_1_2.INIT0 = 16'h0008;
    defparam _add_1_7035_add_4_add_1_add_1_2.INIT1 = 16'h666a;
    defparam _add_1_7035_add_4_add_1_add_1_2.INJECT1_0 = "NO";
    defparam _add_1_7035_add_4_add_1_add_1_2.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_43 (.A(n108), .B(n111), .C(n109_adj_219), 
         .D(n107_adj_218), .Z(n37210)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_43.init = 16'hfffe;
    CCU2C add_7644_31 (.A0(n4647), .B0(n30950), .C0(n64_adj_703), .D0(n4683), 
          .A1(n4646), .B1(n30950), .C1(n64_adj_703), .D1(n4682), .CIN(n32756), 
          .S0(n4752), .S1(n4751));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_31.INIT0 = 16'ha9aa;
    defparam add_7644_31.INIT1 = 16'ha9aa;
    defparam add_7644_31.INJECT1_0 = "NO";
    defparam add_7644_31.INJECT1_1 = "NO";
    CCU2C add_7644_29 (.A0(n4649), .B0(n30950), .C0(n64_adj_703), .D0(n4352), 
          .A1(n4648), .B1(n30950), .C1(n64_adj_703), .D1(n4465), .CIN(n32755), 
          .COUT(n32756), .S0(n4754), .S1(n4753));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_29.INIT0 = 16'ha9aa;
    defparam add_7644_29.INIT1 = 16'ha9aa;
    defparam add_7644_29.INJECT1_0 = "NO";
    defparam add_7644_29.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1109 (.A(n109_adj_219), .B(n108), .Z(n42808)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1109.init = 16'heeee;
    LUT4 i25772_4_lut (.A(n42442), .B(n42441), .C(n42443), .D(n39685), 
         .Z(n39712)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25772_4_lut.init = 16'hfeff;
    LUT4 div_4016_LessThan_3066_i16_3_lut_3_lut (.A(n4659), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n16_adj_676)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i16_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_2153_i50 (.BLUT(n42_adj_387), .ALUT(n48_adj_390), 
          .C0(n38012), .Z(n50_adj_391));
    LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.A(n109_adj_219), .B(n108), .C(n42809), 
         .D(n42810), .Z(n36956)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_44.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i33_2_lut_rep_780 (.A(n4661), .B(n118_adj_225), 
         .Z(n42479)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i33_2_lut_rep_780.init = 16'h6666;
    LUT4 i23187_4_lut (.A(n42607), .B(n42609), .C(n42608), .D(n38431), 
         .Z(n38447)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23187_4_lut.init = 16'h1011;
    LUT4 i24425_4_lut (.A(n42444), .B(n42446), .C(n42445), .D(n39656), 
         .Z(n39685)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24425_4_lut.init = 16'h0100;
    IB U_in_pad_435 (.I(U_in[435]), .O(U_in_c_435));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_436 (.I(U_in[436]), .O(U_in_c_436));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_437 (.I(U_in[437]), .O(U_in_c_437));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_438 (.I(U_in[438]), .O(U_in_c_438));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_439 (.I(U_in[439]), .O(U_in_c_439));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_440 (.I(U_in[440]), .O(U_in_c_440));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_441 (.I(U_in[441]), .O(U_in_c_441));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_442 (.I(U_in[442]), .O(U_in_c_442));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_443 (.I(U_in[443]), .O(U_in_c_443));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_444 (.I(U_in[444]), .O(U_in_c_444));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_445 (.I(U_in[445]), .O(U_in_c_445));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_446 (.I(U_in[446]), .O(U_in_c_446));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_447 (.I(U_in[447]), .O(U_in_c_447));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_448 (.I(U_in[448]), .O(U_in_c_448));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_449 (.I(U_in[449]), .O(U_in_c_449));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_450 (.I(U_in[450]), .O(U_in_c_450));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7644_27 (.A0(n4651), .B0(n30950), .C0(n64_adj_703), .D0(n4117), 
          .A1(n4650), .B1(n30950), .C1(n64_adj_703), .D1(n4236), .CIN(n32754), 
          .COUT(n32755), .S0(n4756), .S1(n4755));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_27.INIT0 = 16'ha9aa;
    defparam add_7644_27.INIT1 = 16'ha9aa;
    defparam add_7644_27.INJECT1_0 = "NO";
    defparam add_7644_27.INJECT1_1 = "NO";
    CCU2C add_7644_25 (.A0(n4653), .B0(n30950), .C0(n64_adj_703), .D0(n3870), 
          .A1(n4652), .B1(n30950), .C1(n64_adj_703), .D1(n3995), .CIN(n32753), 
          .COUT(n32754), .S0(n4758), .S1(n4757));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_25.INIT0 = 16'ha9aa;
    defparam add_7644_25.INIT1 = 16'ha9aa;
    defparam add_7644_25.INJECT1_0 = "NO";
    defparam add_7644_25.INJECT1_1 = "NO";
    CCU2C add_7644_23 (.A0(n4655), .B0(n30950), .C0(n64_adj_703), .D0(n3611), 
          .A1(n4654), .B1(n30950), .C1(n64_adj_703), .D1(n3871), .CIN(n32752), 
          .COUT(n32753), .S0(n4760), .S1(n4759));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_23.INIT0 = 16'ha9aa;
    defparam add_7644_23.INIT1 = 16'ha9aa;
    defparam add_7644_23.INJECT1_0 = "NO";
    defparam add_7644_23.INJECT1_1 = "NO";
    CCU2C add_7644_21 (.A0(n4657), .B0(n30950), .C0(n64_adj_703), .D0(n3340), 
          .A1(n4656), .B1(n30950), .C1(n64_adj_703), .D1(n3477), .CIN(n32751), 
          .COUT(n32752), .S0(n4762), .S1(n4761));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_21.INIT0 = 16'ha9aa;
    defparam add_7644_21.INIT1 = 16'ha9aa;
    defparam add_7644_21.INJECT1_0 = "NO";
    defparam add_7644_21.INJECT1_1 = "NO";
    CCU2C add_7644_19 (.A0(n4659), .B0(n30950), .C0(n64_adj_703), .D0(n3057), 
          .A1(n4658), .B1(n30950), .C1(n64_adj_703), .D1(n3479), .CIN(n32750), 
          .COUT(n32751), .S0(n4764), .S1(n4763));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_19.INIT0 = 16'ha9aa;
    defparam add_7644_19.INIT1 = 16'ha9aa;
    defparam add_7644_19.INJECT1_0 = "NO";
    defparam add_7644_19.INJECT1_1 = "NO";
    CCU2C add_7644_17 (.A0(n4661), .B0(n30950), .C0(n64_adj_703), .D0(n2762), 
          .A1(n4660), .B1(n30950), .C1(n64_adj_703), .D1(n2911), .CIN(n32749), 
          .COUT(n32750), .S0(n4766), .S1(n4765));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_17.INIT0 = 16'ha9aa;
    defparam add_7644_17.INIT1 = 16'ha9aa;
    defparam add_7644_17.INJECT1_0 = "NO";
    defparam add_7644_17.INJECT1_1 = "NO";
    CCU2C add_7644_15 (.A0(n4663), .B0(n30950), .C0(n64_adj_703), .D0(n2455), 
          .A1(n4662), .B1(n30950), .C1(n64_adj_703), .D1(n3060), .CIN(n32748), 
          .COUT(n32749), .S0(n4768), .S1(n4767));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_15.INIT0 = 16'ha9aa;
    defparam add_7644_15.INIT1 = 16'ha9aa;
    defparam add_7644_15.INJECT1_0 = "NO";
    defparam add_7644_15.INJECT1_1 = "NO";
    CCU2C add_7644_13 (.A0(n4665), .B0(n30950), .C0(n64_adj_703), .D0(n2298), 
          .A1(n4664), .B1(n30950), .C1(n64_adj_703), .D1(n2456), .CIN(n32747), 
          .COUT(n32748), .S0(n4770), .S1(n4769));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_13.INIT0 = 16'ha9aa;
    defparam add_7644_13.INIT1 = 16'ha9aa;
    defparam add_7644_13.INJECT1_0 = "NO";
    defparam add_7644_13.INJECT1_1 = "NO";
    CCU2C add_7644_11 (.A0(n4667), .B0(n30950), .C0(n64_adj_703), .D0(n1805), 
          .A1(n4666), .B1(n30950), .C1(n64_adj_703), .D1(n2137), .CIN(n32746), 
          .COUT(n32747), .S0(n4772), .S1(n4771));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_11.INIT0 = 16'ha9aa;
    defparam add_7644_11.INIT1 = 16'ha9aa;
    defparam add_7644_11.INJECT1_0 = "NO";
    defparam add_7644_11.INJECT1_1 = "NO";
    CCU2C add_7644_9 (.A0(n4669), .B0(n30950), .C0(n64_adj_703), .D0(n1462), 
          .A1(n4668), .B1(n30950), .C1(n64_adj_703), .D1(n1635), .CIN(n32745), 
          .COUT(n32746), .S0(n4774), .S1(n4773));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_9.INIT0 = 16'ha9aa;
    defparam add_7644_9.INIT1 = 16'ha9aa;
    defparam add_7644_9.INJECT1_0 = "NO";
    defparam add_7644_9.INJECT1_1 = "NO";
    CCU2C add_7644_7 (.A0(n4671), .B0(n30950), .C0(n64_adj_703), .D0(n2142), 
          .A1(n4670), .B1(n30950), .C1(n64_adj_703), .D1(n2141), .CIN(n32744), 
          .COUT(n32745), .S0(n4776), .S1(n4775));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_7.INIT0 = 16'ha9aa;
    defparam add_7644_7.INIT1 = 16'ha9aa;
    defparam add_7644_7.INJECT1_0 = "NO";
    defparam add_7644_7.INJECT1_1 = "NO";
    CCU2C add_7644_5 (.A0(n4673), .B0(n30950), .C0(n64_adj_703), .D0(n42824), 
          .A1(n4672), .B1(n30950), .C1(n64_adj_703), .D1(n42822), .CIN(n32743), 
          .COUT(n32744), .S0(n4778), .S1(n4777));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_5.INIT0 = 16'ha9aa;
    defparam add_7644_5.INIT1 = 16'ha9aa;
    defparam add_7644_5.INJECT1_0 = "NO";
    defparam add_7644_5.INJECT1_1 = "NO";
    CCU2C add_7644_3 (.A0(n892), .B0(n30950), .C0(n64_adj_703), .D0(n42827), 
          .A1(n4674), .B1(n30950), .C1(n64_adj_703), .D1(n42823), .CIN(n32742), 
          .COUT(n32743), .S0(n4780), .S1(n4779));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_3.INIT0 = 16'ha9aa;
    defparam add_7644_3.INIT1 = 16'ha9aa;
    defparam add_7644_3.INJECT1_0 = "NO";
    defparam add_7644_3.INJECT1_1 = "NO";
    CCU2C add_7644_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_703), .B1(n30950), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32742));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7644_1.INIT0 = 16'h0000;
    defparam add_7644_1.INIT1 = 16'heee1;
    defparam add_7644_1.INJECT1_0 = "NO";
    defparam add_7644_1.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_1761_i38_4_lut (.A(n132), .B(n131_adj_234), .C(n2724), 
         .D(n877), .Z(n38)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i38_4_lut.init = 16'h0c8e;
    CCU2C add_7643_31 (.A0(n4538), .B0(n42792), .C0(n64_adj_670), .D0(n4683), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32738), 
          .S0(n4646));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_31.INIT0 = 16'ha9aa;
    defparam add_7643_31.INIT1 = 16'h0000;
    defparam add_7643_31.INJECT1_0 = "NO";
    defparam add_7643_31.INJECT1_1 = "NO";
    LUT4 i24396_4_lut (.A(n42448), .B(n42447), .C(n42449), .D(n39641), 
         .Z(n39656)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24396_4_lut.init = 16'h0100;
    LUT4 div_4016_LessThan_2513_i51_2_lut_rep_910 (.A(n3833), .B(n116_adj_224), 
         .Z(n42609)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i51_2_lut_rep_910.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_45 (.A(n109_adj_219), .B(n108), .C(n106_adj_217), 
         .D(n107_adj_218), .Z(n36992)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_45.init = 16'hfffe;
    LUT4 i25824_4_lut (.A(n42488), .B(n42487), .C(n39328), .D(n39331), 
         .Z(n39349)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25824_4_lut.init = 16'hffef;
    LUT4 i23171_4_lut (.A(n42610), .B(n45_adj_483), .C(n33_adj_476), .D(n38384), 
         .Z(n38431)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23171_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_2513_i30_3_lut_3_lut (.A(n3833), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n30_adj_474)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24046_4_lut (.A(n42492), .B(n42493), .C(n42502), .D(n39226), 
         .Z(n39306)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24046_4_lut.init = 16'h1011;
    LUT4 i23966_4_lut (.A(n42501), .B(n42503), .C(n42504), .D(n39214), 
         .Z(n39226)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23966_4_lut.init = 16'h1011;
    IB U_in_pad_451 (.I(U_in[451]), .O(U_in_c_451));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_452 (.I(U_in[452]), .O(U_in_c_452));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_453 (.I(U_in[453]), .O(U_in_c_453));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_454 (.I(U_in[454]), .O(U_in_c_454));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_455 (.I(U_in[455]), .O(U_in_c_455));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_456 (.I(U_in[456]), .O(U_in_c_456));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_457 (.I(U_in[457]), .O(U_in_c_457));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_458 (.I(U_in[458]), .O(U_in_c_458));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_459 (.I(U_in[459]), .O(U_in_c_459));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_460 (.I(U_in[460]), .O(U_in_c_460));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_461 (.I(U_in[461]), .O(U_in_c_461));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_462 (.I(U_in[462]), .O(U_in_c_462));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_463 (.I(U_in[463]), .O(U_in_c_463));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_464 (.I(U_in[464]), .O(U_in_c_464));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_465 (.I(U_in[465]), .O(U_in_c_465));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7643_29 (.A0(n4540), .B0(n42792), .C0(n64_adj_670), .D0(n4352), 
          .A1(n4539), .B1(n42792), .C1(n64_adj_670), .D1(n4465), .CIN(n32737), 
          .COUT(n32738), .S0(n4648), .S1(n4647));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_29.INIT0 = 16'ha9aa;
    defparam add_7643_29.INIT1 = 16'ha9aa;
    defparam add_7643_29.INJECT1_0 = "NO";
    defparam add_7643_29.INJECT1_1 = "NO";
    CCU2C add_7643_27 (.A0(n4542), .B0(n42792), .C0(n64_adj_670), .D0(n4117), 
          .A1(n4541), .B1(n42792), .C1(n64_adj_670), .D1(n4236), .CIN(n32736), 
          .COUT(n32737), .S0(n4650), .S1(n4649));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_27.INIT0 = 16'ha9aa;
    defparam add_7643_27.INIT1 = 16'ha9aa;
    defparam add_7643_27.INJECT1_0 = "NO";
    defparam add_7643_27.INJECT1_1 = "NO";
    CCU2C add_7643_25 (.A0(n4544), .B0(n42792), .C0(n64_adj_670), .D0(n3870), 
          .A1(n4543), .B1(n42792), .C1(n64_adj_670), .D1(n3995), .CIN(n32735), 
          .COUT(n32736), .S0(n4652), .S1(n4651));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_25.INIT0 = 16'ha9aa;
    defparam add_7643_25.INIT1 = 16'ha9aa;
    defparam add_7643_25.INJECT1_0 = "NO";
    defparam add_7643_25.INJECT1_1 = "NO";
    CCU2C add_7643_23 (.A0(n4546), .B0(n42792), .C0(n64_adj_670), .D0(n3611), 
          .A1(n4545), .B1(n42792), .C1(n64_adj_670), .D1(n3871), .CIN(n32734), 
          .COUT(n32735), .S0(n4654), .S1(n4653));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_23.INIT0 = 16'ha9aa;
    defparam add_7643_23.INIT1 = 16'ha9aa;
    defparam add_7643_23.INJECT1_0 = "NO";
    defparam add_7643_23.INJECT1_1 = "NO";
    CCU2C add_7643_21 (.A0(n4548), .B0(n42792), .C0(n64_adj_670), .D0(n3340), 
          .A1(n4547), .B1(n42792), .C1(n64_adj_670), .D1(n3477), .CIN(n32733), 
          .COUT(n32734), .S0(n4656), .S1(n4655));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_21.INIT0 = 16'ha9aa;
    defparam add_7643_21.INIT1 = 16'ha9aa;
    defparam add_7643_21.INJECT1_0 = "NO";
    defparam add_7643_21.INJECT1_1 = "NO";
    CCU2C add_7643_19 (.A0(n4550), .B0(n42792), .C0(n64_adj_670), .D0(n3057), 
          .A1(n4549), .B1(n42792), .C1(n64_adj_670), .D1(n3479), .CIN(n32732), 
          .COUT(n32733), .S0(n4658), .S1(n4657));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_19.INIT0 = 16'ha9aa;
    defparam add_7643_19.INIT1 = 16'ha9aa;
    defparam add_7643_19.INJECT1_0 = "NO";
    defparam add_7643_19.INJECT1_1 = "NO";
    CCU2C add_7643_17 (.A0(n4552), .B0(n42792), .C0(n64_adj_670), .D0(n2762), 
          .A1(n4551), .B1(n42792), .C1(n64_adj_670), .D1(n2911), .CIN(n32731), 
          .COUT(n32732), .S0(n4660), .S1(n4659));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_17.INIT0 = 16'ha9aa;
    defparam add_7643_17.INIT1 = 16'ha9aa;
    defparam add_7643_17.INJECT1_0 = "NO";
    defparam add_7643_17.INJECT1_1 = "NO";
    CCU2C add_7643_15 (.A0(n4554), .B0(n42792), .C0(n64_adj_670), .D0(n2455), 
          .A1(n4553), .B1(n42792), .C1(n64_adj_670), .D1(n3060), .CIN(n32730), 
          .COUT(n32731), .S0(n4662), .S1(n4661));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_15.INIT0 = 16'ha9aa;
    defparam add_7643_15.INIT1 = 16'ha9aa;
    defparam add_7643_15.INJECT1_0 = "NO";
    defparam add_7643_15.INJECT1_1 = "NO";
    CCU2C add_7643_13 (.A0(n4556), .B0(n42792), .C0(n64_adj_670), .D0(n2298), 
          .A1(n4555), .B1(n42792), .C1(n64_adj_670), .D1(n2456), .CIN(n32729), 
          .COUT(n32730), .S0(n4664), .S1(n4663));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_13.INIT0 = 16'ha9aa;
    defparam add_7643_13.INIT1 = 16'ha9aa;
    defparam add_7643_13.INJECT1_0 = "NO";
    defparam add_7643_13.INJECT1_1 = "NO";
    CCU2C add_7643_11 (.A0(n4558), .B0(n42792), .C0(n64_adj_670), .D0(n1805), 
          .A1(n4557), .B1(n42792), .C1(n64_adj_670), .D1(n2137), .CIN(n32728), 
          .COUT(n32729), .S0(n4666), .S1(n4665));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_11.INIT0 = 16'ha9aa;
    defparam add_7643_11.INIT1 = 16'ha9aa;
    defparam add_7643_11.INJECT1_0 = "NO";
    defparam add_7643_11.INJECT1_1 = "NO";
    CCU2C add_7643_9 (.A0(n4560), .B0(n42792), .C0(n64_adj_670), .D0(n1462), 
          .A1(n4559), .B1(n42792), .C1(n64_adj_670), .D1(n1635), .CIN(n32727), 
          .COUT(n32728), .S0(n4668), .S1(n4667));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_9.INIT0 = 16'ha9aa;
    defparam add_7643_9.INIT1 = 16'ha9aa;
    defparam add_7643_9.INJECT1_0 = "NO";
    defparam add_7643_9.INJECT1_1 = "NO";
    CCU2C add_7643_7 (.A0(n4562), .B0(n42792), .C0(n64_adj_670), .D0(n2142), 
          .A1(n4561), .B1(n42792), .C1(n64_adj_670), .D1(n2141), .CIN(n32726), 
          .COUT(n32727), .S0(n4670), .S1(n4669));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_7.INIT0 = 16'ha9aa;
    defparam add_7643_7.INIT1 = 16'ha9aa;
    defparam add_7643_7.INJECT1_0 = "NO";
    defparam add_7643_7.INJECT1_1 = "NO";
    CCU2C add_7643_5 (.A0(n4564), .B0(n42792), .C0(n64_adj_670), .D0(n42824), 
          .A1(n4563), .B1(n42792), .C1(n64_adj_670), .D1(n42822), .CIN(n32725), 
          .COUT(n32726), .S0(n4672), .S1(n4671));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_5.INIT0 = 16'ha9aa;
    defparam add_7643_5.INIT1 = 16'ha9aa;
    defparam add_7643_5.INJECT1_0 = "NO";
    defparam add_7643_5.INJECT1_1 = "NO";
    CCU2C add_7643_3 (.A0(n891), .B0(n42792), .C0(n64_adj_670), .D0(n42827), 
          .A1(n4565), .B1(n42792), .C1(n64_adj_670), .D1(n42823), .CIN(n32724), 
          .COUT(n32725), .S0(n4674), .S1(n4673));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_3.INIT0 = 16'ha9aa;
    defparam add_7643_3.INIT1 = 16'ha9aa;
    defparam add_7643_3.INJECT1_0 = "NO";
    defparam add_7643_3.INJECT1_1 = "NO";
    CCU2C add_7643_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_670), .B1(n42792), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32724));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7643_1.INIT0 = 16'h0000;
    defparam add_7643_1.INIT1 = 16'heee1;
    defparam add_7643_1.INJECT1_0 = "NO";
    defparam add_7643_1.INJECT1_1 = "NO";
    LUT4 i25642_4_lut_4_lut (.A(n42611), .B(n38411), .C(n38_adj_479), 
         .D(n24_adj_471), .Z(n40_adj_480)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25642_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_3066_i18_3_lut_3_lut (.A(n4661), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n18_adj_677)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24381_4_lut (.A(n42450), .B(n42452), .C(n42451), .D(n39614), 
         .Z(n39641)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24381_4_lut.init = 16'h5455;
    PFUMX div_4016_LessThan_2058_i62 (.BLUT(n56_adj_374), .ALUT(n60_adj_376), 
          .C0(n37963), .Z(n62_adj_377));
    LUT4 i24354_4_lut (.A(n42454), .B(n42453), .C(n42455), .D(n39591), 
         .Z(n39614)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24354_4_lut.init = 16'h0100;
    IB U_in_pad_466 (.I(U_in[466]), .O(U_in_c_466));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_467 (.I(U_in[467]), .O(U_in_c_467));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_468 (.I(U_in[468]), .O(U_in_c_468));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_469 (.I(U_in[469]), .O(U_in_c_469));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_470 (.I(U_in[470]), .O(U_in_c_470));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_471 (.I(U_in[471]), .O(U_in_c_471));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_472 (.I(U_in[472]), .O(U_in_c_472));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_473 (.I(U_in[473]), .O(U_in_c_473));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_474 (.I(U_in[474]), .O(U_in_c_474));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_475 (.I(U_in[475]), .O(U_in_c_475));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_476 (.I(U_in[476]), .O(U_in_c_476));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_477 (.I(U_in[477]), .O(U_in_c_477));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_478 (.I(U_in[478]), .O(U_in_c_478));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_479 (.I(U_in[479]), .O(U_in_c_479));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7642_29 (.A0(n4428), .B0(n30944), .C0(n64_adj_640), .D0(n4352), 
          .A1(n4427), .B1(n30944), .C1(n64_adj_640), .D1(n4465), .CIN(n32719), 
          .S0(n4539), .S1(n4538));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_29.INIT0 = 16'ha9aa;
    defparam add_7642_29.INIT1 = 16'ha9aa;
    defparam add_7642_29.INJECT1_0 = "NO";
    defparam add_7642_29.INJECT1_1 = "NO";
    CCU2C add_7642_27 (.A0(n4430), .B0(n30944), .C0(n64_adj_640), .D0(n4117), 
          .A1(n4429), .B1(n30944), .C1(n64_adj_640), .D1(n4236), .CIN(n32718), 
          .COUT(n32719), .S0(n4541), .S1(n4540));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_27.INIT0 = 16'ha9aa;
    defparam add_7642_27.INIT1 = 16'ha9aa;
    defparam add_7642_27.INJECT1_0 = "NO";
    defparam add_7642_27.INJECT1_1 = "NO";
    CCU2C add_7642_25 (.A0(n4432), .B0(n30944), .C0(n64_adj_640), .D0(n3870), 
          .A1(n4431), .B1(n30944), .C1(n64_adj_640), .D1(n3995), .CIN(n32717), 
          .COUT(n32718), .S0(n4543), .S1(n4542));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_25.INIT0 = 16'ha9aa;
    defparam add_7642_25.INIT1 = 16'ha9aa;
    defparam add_7642_25.INJECT1_0 = "NO";
    defparam add_7642_25.INJECT1_1 = "NO";
    CCU2C add_7642_23 (.A0(n4434), .B0(n30944), .C0(n64_adj_640), .D0(n3611), 
          .A1(n4433), .B1(n30944), .C1(n64_adj_640), .D1(n3871), .CIN(n32716), 
          .COUT(n32717), .S0(n4545), .S1(n4544));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_23.INIT0 = 16'ha9aa;
    defparam add_7642_23.INIT1 = 16'ha9aa;
    defparam add_7642_23.INJECT1_0 = "NO";
    defparam add_7642_23.INJECT1_1 = "NO";
    CCU2C add_7642_21 (.A0(n4436), .B0(n30944), .C0(n64_adj_640), .D0(n3340), 
          .A1(n4435), .B1(n30944), .C1(n64_adj_640), .D1(n3477), .CIN(n32715), 
          .COUT(n32716), .S0(n4547), .S1(n4546));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_21.INIT0 = 16'ha9aa;
    defparam add_7642_21.INIT1 = 16'ha9aa;
    defparam add_7642_21.INJECT1_0 = "NO";
    defparam add_7642_21.INJECT1_1 = "NO";
    CCU2C add_7642_19 (.A0(n4438), .B0(n30944), .C0(n64_adj_640), .D0(n3057), 
          .A1(n4437), .B1(n30944), .C1(n64_adj_640), .D1(n3479), .CIN(n32714), 
          .COUT(n32715), .S0(n4549), .S1(n4548));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_19.INIT0 = 16'ha9aa;
    defparam add_7642_19.INIT1 = 16'ha9aa;
    defparam add_7642_19.INJECT1_0 = "NO";
    defparam add_7642_19.INJECT1_1 = "NO";
    CCU2C add_7642_17 (.A0(n4440), .B0(n30944), .C0(n64_adj_640), .D0(n2762), 
          .A1(n4439), .B1(n30944), .C1(n64_adj_640), .D1(n2911), .CIN(n32713), 
          .COUT(n32714), .S0(n4551), .S1(n4550));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_17.INIT0 = 16'ha9aa;
    defparam add_7642_17.INIT1 = 16'ha9aa;
    defparam add_7642_17.INJECT1_0 = "NO";
    defparam add_7642_17.INJECT1_1 = "NO";
    CCU2C add_7642_15 (.A0(n4442), .B0(n30944), .C0(n64_adj_640), .D0(n2455), 
          .A1(n4441), .B1(n30944), .C1(n64_adj_640), .D1(n3060), .CIN(n32712), 
          .COUT(n32713), .S0(n4553), .S1(n4552));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_15.INIT0 = 16'ha9aa;
    defparam add_7642_15.INIT1 = 16'ha9aa;
    defparam add_7642_15.INJECT1_0 = "NO";
    defparam add_7642_15.INJECT1_1 = "NO";
    CCU2C add_7642_13 (.A0(n4444), .B0(n30944), .C0(n64_adj_640), .D0(n2298), 
          .A1(n4443), .B1(n30944), .C1(n64_adj_640), .D1(n2456), .CIN(n32711), 
          .COUT(n32712), .S0(n4555), .S1(n4554));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_13.INIT0 = 16'ha9aa;
    defparam add_7642_13.INIT1 = 16'ha9aa;
    defparam add_7642_13.INJECT1_0 = "NO";
    defparam add_7642_13.INJECT1_1 = "NO";
    CCU2C add_7642_11 (.A0(n4446), .B0(n30944), .C0(n64_adj_640), .D0(n1805), 
          .A1(n4445), .B1(n30944), .C1(n64_adj_640), .D1(n2137), .CIN(n32710), 
          .COUT(n32711), .S0(n4557), .S1(n4556));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_11.INIT0 = 16'ha9aa;
    defparam add_7642_11.INIT1 = 16'ha9aa;
    defparam add_7642_11.INJECT1_0 = "NO";
    defparam add_7642_11.INJECT1_1 = "NO";
    CCU2C add_7642_9 (.A0(n4448), .B0(n30944), .C0(n64_adj_640), .D0(n1462), 
          .A1(n4447), .B1(n30944), .C1(n64_adj_640), .D1(n1635), .CIN(n32709), 
          .COUT(n32710), .S0(n4559), .S1(n4558));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_9.INIT0 = 16'ha9aa;
    defparam add_7642_9.INIT1 = 16'ha9aa;
    defparam add_7642_9.INJECT1_0 = "NO";
    defparam add_7642_9.INJECT1_1 = "NO";
    CCU2C add_7642_7 (.A0(n4450), .B0(n30944), .C0(n64_adj_640), .D0(n2142), 
          .A1(n4449), .B1(n30944), .C1(n64_adj_640), .D1(n2141), .CIN(n32708), 
          .COUT(n32709), .S0(n4561), .S1(n4560));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_7.INIT0 = 16'ha9aa;
    defparam add_7642_7.INIT1 = 16'ha9aa;
    defparam add_7642_7.INJECT1_0 = "NO";
    defparam add_7642_7.INJECT1_1 = "NO";
    CCU2C add_7642_5 (.A0(n4452), .B0(n30944), .C0(n64_adj_640), .D0(n42824), 
          .A1(n4451), .B1(n30944), .C1(n64_adj_640), .D1(n42822), .CIN(n32707), 
          .COUT(n32708), .S0(n4563), .S1(n4562));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_5.INIT0 = 16'ha9aa;
    defparam add_7642_5.INIT1 = 16'ha9aa;
    defparam add_7642_5.INJECT1_0 = "NO";
    defparam add_7642_5.INJECT1_1 = "NO";
    CCU2C add_7642_3 (.A0(n890), .B0(n30944), .C0(n64_adj_640), .D0(n42827), 
          .A1(n4453), .B1(n30944), .C1(n64_adj_640), .D1(n42823), .CIN(n32706), 
          .COUT(n32707), .S0(n4565), .S1(n4564));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_3.INIT0 = 16'ha9aa;
    defparam add_7642_3.INIT1 = 16'ha9aa;
    defparam add_7642_3.INJECT1_0 = "NO";
    defparam add_7642_3.INJECT1_1 = "NO";
    CCU2C add_7642_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_640), .B1(n30944), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32706));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7642_1.INIT0 = 16'h0000;
    defparam add_7642_1.INIT1 = 16'heee1;
    defparam add_7642_1.INJECT1_0 = "NO";
    defparam add_7642_1.INJECT1_1 = "NO";
    CCU2C add_7641_29 (.A0(n4313), .B0(n42794), .C0(n64_adj_608), .D0(n4352), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32702), 
          .S0(n4427));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_29.INIT0 = 16'ha9aa;
    defparam add_7641_29.INIT1 = 16'h0000;
    defparam add_7641_29.INJECT1_0 = "NO";
    defparam add_7641_29.INJECT1_1 = "NO";
    CCU2C add_7641_27 (.A0(n4315), .B0(n42794), .C0(n64_adj_608), .D0(n4117), 
          .A1(n4314), .B1(n42794), .C1(n64_adj_608), .D1(n4236), .CIN(n32701), 
          .COUT(n32702), .S0(n4429), .S1(n4428));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_27.INIT0 = 16'ha9aa;
    defparam add_7641_27.INIT1 = 16'ha9aa;
    defparam add_7641_27.INJECT1_0 = "NO";
    defparam add_7641_27.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_2993_i59_2_lut (.A(n4540), .B(n106_adj_217), 
         .Z(n39328)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i59_2_lut.init = 16'h9999;
    LUT4 div_4016_LessThan_3137_i15_2_lut_rep_764 (.A(n4775), .B(n126), 
         .Z(n42463)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i15_2_lut_rep_764.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(n110_adj_220), .B(n113_adj_222), 
         .C(n37272), .D(n42811), .Z(n37148)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'hfffe;
    LUT4 i25822_4_lut (.A(n42487), .B(n39328), .C(n42502), .D(n39228), 
         .Z(n39351)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25822_4_lut.init = 16'hbfbb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_47 (.A(n110_adj_220), .B(n113_adj_222), 
         .C(n111), .D(n108), .Z(n37176)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_47.init = 16'hfffe;
    LUT4 i25886_4_lut_4_lut (.A(n42611), .B(n38409), .C(n42602), .D(n42603), 
         .Z(n40092)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25886_4_lut_4_lut.init = 16'hfff4;
    LUT4 i24331_4_lut (.A(n42456), .B(n42457), .C(n29_adj_719), .D(n39576), 
         .Z(n39591)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24331_4_lut.init = 16'h0001;
    LUT4 i1_3_lut_4_lut_adj_48 (.A(n110_adj_220), .B(n113_adj_222), .C(n111), 
         .D(n109_adj_219), .Z(n37242)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_48.init = 16'hfffe;
    IB U_in_pad_480 (.I(U_in[480]), .O(U_in_c_480));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_481 (.I(U_in[481]), .O(U_in_c_481));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_482 (.I(U_in[482]), .O(U_in_c_482));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_483 (.I(U_in[483]), .O(U_in_c_483));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_484 (.I(U_in[484]), .O(U_in_c_484));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_485 (.I(U_in[485]), .O(U_in_c_485));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_486 (.I(U_in[486]), .O(U_in_c_486));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_487 (.I(U_in[487]), .O(U_in_c_487));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_488 (.I(U_in[488]), .O(U_in_c_488));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_489 (.I(U_in[489]), .O(U_in_c_489));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_490 (.I(U_in[490]), .O(U_in_c_490));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_491 (.I(U_in[491]), .O(U_in_c_491));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_492 (.I(U_in[492]), .O(U_in_c_492));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7641_25 (.A0(n4317), .B0(n42794), .C0(n64_adj_608), .D0(n3870), 
          .A1(n4316), .B1(n42794), .C1(n64_adj_608), .D1(n3995), .CIN(n32700), 
          .COUT(n32701), .S0(n4431), .S1(n4430));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_25.INIT0 = 16'ha9aa;
    defparam add_7641_25.INIT1 = 16'ha9aa;
    defparam add_7641_25.INJECT1_0 = "NO";
    defparam add_7641_25.INJECT1_1 = "NO";
    CCU2C add_7641_23 (.A0(n4319), .B0(n42794), .C0(n64_adj_608), .D0(n3611), 
          .A1(n4318), .B1(n42794), .C1(n64_adj_608), .D1(n3871), .CIN(n32699), 
          .COUT(n32700), .S0(n4433), .S1(n4432));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_23.INIT0 = 16'ha9aa;
    defparam add_7641_23.INIT1 = 16'ha9aa;
    defparam add_7641_23.INJECT1_0 = "NO";
    defparam add_7641_23.INJECT1_1 = "NO";
    CCU2C add_7641_21 (.A0(n4321), .B0(n42794), .C0(n64_adj_608), .D0(n3340), 
          .A1(n4320), .B1(n42794), .C1(n64_adj_608), .D1(n3477), .CIN(n32698), 
          .COUT(n32699), .S0(n4435), .S1(n4434));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_21.INIT0 = 16'ha9aa;
    defparam add_7641_21.INIT1 = 16'ha9aa;
    defparam add_7641_21.INJECT1_0 = "NO";
    defparam add_7641_21.INJECT1_1 = "NO";
    CCU2C add_7641_19 (.A0(n4323), .B0(n42794), .C0(n64_adj_608), .D0(n3057), 
          .A1(n4322), .B1(n42794), .C1(n64_adj_608), .D1(n3479), .CIN(n32697), 
          .COUT(n32698), .S0(n4437), .S1(n4436));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_19.INIT0 = 16'ha9aa;
    defparam add_7641_19.INIT1 = 16'ha9aa;
    defparam add_7641_19.INJECT1_0 = "NO";
    defparam add_7641_19.INJECT1_1 = "NO";
    CCU2C add_7641_17 (.A0(n4325), .B0(n42794), .C0(n64_adj_608), .D0(n2762), 
          .A1(n4324), .B1(n42794), .C1(n64_adj_608), .D1(n2911), .CIN(n32696), 
          .COUT(n32697), .S0(n4439), .S1(n4438));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_17.INIT0 = 16'ha9aa;
    defparam add_7641_17.INIT1 = 16'ha9aa;
    defparam add_7641_17.INJECT1_0 = "NO";
    defparam add_7641_17.INJECT1_1 = "NO";
    CCU2C add_7641_15 (.A0(n4327), .B0(n42794), .C0(n64_adj_608), .D0(n2455), 
          .A1(n4326), .B1(n42794), .C1(n64_adj_608), .D1(n3060), .CIN(n32695), 
          .COUT(n32696), .S0(n4441), .S1(n4440));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_15.INIT0 = 16'ha9aa;
    defparam add_7641_15.INIT1 = 16'ha9aa;
    defparam add_7641_15.INJECT1_0 = "NO";
    defparam add_7641_15.INJECT1_1 = "NO";
    CCU2C add_7641_13 (.A0(n4329), .B0(n42794), .C0(n64_adj_608), .D0(n2298), 
          .A1(n4328), .B1(n42794), .C1(n64_adj_608), .D1(n2456), .CIN(n32694), 
          .COUT(n32695), .S0(n4443), .S1(n4442));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_13.INIT0 = 16'ha9aa;
    defparam add_7641_13.INIT1 = 16'ha9aa;
    defparam add_7641_13.INJECT1_0 = "NO";
    defparam add_7641_13.INJECT1_1 = "NO";
    CCU2C add_7641_11 (.A0(n4331), .B0(n42794), .C0(n64_adj_608), .D0(n1805), 
          .A1(n4330), .B1(n42794), .C1(n64_adj_608), .D1(n2137), .CIN(n32693), 
          .COUT(n32694), .S0(n4445), .S1(n4444));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_11.INIT0 = 16'ha9aa;
    defparam add_7641_11.INIT1 = 16'ha9aa;
    defparam add_7641_11.INJECT1_0 = "NO";
    defparam add_7641_11.INJECT1_1 = "NO";
    CCU2C add_7641_9 (.A0(n4333), .B0(n42794), .C0(n64_adj_608), .D0(n1462), 
          .A1(n4332), .B1(n42794), .C1(n64_adj_608), .D1(n1635), .CIN(n32692), 
          .COUT(n32693), .S0(n4447), .S1(n4446));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_9.INIT0 = 16'ha9aa;
    defparam add_7641_9.INIT1 = 16'ha9aa;
    defparam add_7641_9.INJECT1_0 = "NO";
    defparam add_7641_9.INJECT1_1 = "NO";
    CCU2C add_7641_7 (.A0(n4335), .B0(n42794), .C0(n64_adj_608), .D0(n2142), 
          .A1(n4334), .B1(n42794), .C1(n64_adj_608), .D1(n2141), .CIN(n32691), 
          .COUT(n32692), .S0(n4449), .S1(n4448));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_7.INIT0 = 16'ha9aa;
    defparam add_7641_7.INIT1 = 16'ha9aa;
    defparam add_7641_7.INJECT1_0 = "NO";
    defparam add_7641_7.INJECT1_1 = "NO";
    CCU2C add_7641_5 (.A0(n4337), .B0(n42794), .C0(n64_adj_608), .D0(n42824), 
          .A1(n4336), .B1(n42794), .C1(n64_adj_608), .D1(n42822), .CIN(n32690), 
          .COUT(n32691), .S0(n4451), .S1(n4450));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_5.INIT0 = 16'ha9aa;
    defparam add_7641_5.INIT1 = 16'ha9aa;
    defparam add_7641_5.INJECT1_0 = "NO";
    defparam add_7641_5.INJECT1_1 = "NO";
    CCU2C add_7641_3 (.A0(n889), .B0(n42794), .C0(n64_adj_608), .D0(n42827), 
          .A1(n4338), .B1(n42794), .C1(n64_adj_608), .D1(n42823), .CIN(n32689), 
          .COUT(n32690), .S0(n4453), .S1(n4452));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_3.INIT0 = 16'ha9aa;
    defparam add_7641_3.INIT1 = 16'ha9aa;
    defparam add_7641_3.INJECT1_0 = "NO";
    defparam add_7641_3.INJECT1_1 = "NO";
    CCU2C add_7641_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_608), .B1(n42794), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32689));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7641_1.INIT0 = 16'h0000;
    defparam add_7641_1.INIT1 = 16'heee1;
    defparam add_7641_1.INJECT1_0 = "NO";
    defparam add_7641_1.INJECT1_1 = "NO";
    CCU2C add_7640_27 (.A0(n4197), .B0(n30938), .C0(n64_adj_578), .D0(n4117), 
          .A1(n4196), .B1(n30938), .C1(n64_adj_578), .D1(n4236), .CIN(n32684), 
          .S0(n4314), .S1(n4313));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_27.INIT0 = 16'ha9aa;
    defparam add_7640_27.INIT1 = 16'ha9aa;
    defparam add_7640_27.INJECT1_0 = "NO";
    defparam add_7640_27.INJECT1_1 = "NO";
    CCU2C add_7640_25 (.A0(n4199), .B0(n30938), .C0(n64_adj_578), .D0(n3870), 
          .A1(n4198), .B1(n30938), .C1(n64_adj_578), .D1(n3995), .CIN(n32683), 
          .COUT(n32684), .S0(n4316), .S1(n4315));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_25.INIT0 = 16'ha9aa;
    defparam add_7640_25.INIT1 = 16'ha9aa;
    defparam add_7640_25.INJECT1_0 = "NO";
    defparam add_7640_25.INJECT1_1 = "NO";
    CCU2C add_7640_23 (.A0(n4201), .B0(n30938), .C0(n64_adj_578), .D0(n3611), 
          .A1(n4200), .B1(n30938), .C1(n64_adj_578), .D1(n3871), .CIN(n32682), 
          .COUT(n32683), .S0(n4318), .S1(n4317));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_23.INIT0 = 16'ha9aa;
    defparam add_7640_23.INIT1 = 16'ha9aa;
    defparam add_7640_23.INJECT1_0 = "NO";
    defparam add_7640_23.INJECT1_1 = "NO";
    CCU2C add_7640_21 (.A0(n4203), .B0(n30938), .C0(n64_adj_578), .D0(n3340), 
          .A1(n4202), .B1(n30938), .C1(n64_adj_578), .D1(n3477), .CIN(n32681), 
          .COUT(n32682), .S0(n4320), .S1(n4319));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_21.INIT0 = 16'ha9aa;
    defparam add_7640_21.INIT1 = 16'ha9aa;
    defparam add_7640_21.INJECT1_0 = "NO";
    defparam add_7640_21.INJECT1_1 = "NO";
    LUT4 i24316_4_lut (.A(n42459), .B(n42458), .C(n42460), .D(n39557), 
         .Z(n39576)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24316_4_lut.init = 16'h0100;
    LUT4 i24297_4_lut (.A(n21_adj_714), .B(n42461), .C(n17_adj_711), .D(n39544), 
         .Z(n39557)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24297_4_lut.init = 16'h1011;
    LUT4 div_4016_i3325_4_lut (.A(n64_adj_328), .B(n22289), .C(n42786), 
         .D(n30905), .Z(n5508)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3325_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_3066_i27_2_lut_rep_781 (.A(n4664), .B(n121_adj_227), 
         .Z(n42480)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i27_2_lut_rep_781.init = 16'h6666;
    LUT4 i1_4_lut_adj_49 (.A(n37054), .B(n36956), .C(n42797), .D(n42798), 
         .Z(n30905)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_49.init = 16'hfffe;
    LUT4 div_4016_LessThan_1862_i36_4_lut (.A(n132), .B(n131_adj_234), .C(n2875), 
         .D(n878), .Z(n36)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i36_4_lut.init = 16'h0c8e;
    LUT4 i1_2_lut_rep_1111 (.A(n111), .B(n110_adj_220), .Z(n42810)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1111.init = 16'heeee;
    LUT4 i23154_4_lut_4_lut (.A(n42611), .B(n38395), .C(n42614), .D(n42612), 
         .Z(n38414)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23154_4_lut_4_lut.init = 16'h0004;
    LUT4 div_4016_LessThan_2513_i45_2_lut (.A(n3836), .B(n119_adj_226), 
         .Z(n45_adj_483)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i45_2_lut.init = 16'h6666;
    IB U_in_pad_493 (.I(U_in[493]), .O(U_in_c_493));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_494 (.I(U_in[494]), .O(U_in_c_494));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_495 (.I(U_in[495]), .O(U_in_c_495));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_496 (.I(U_in[496]), .O(U_in_c_496));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_497 (.I(U_in[497]), .O(U_in_c_497));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_498 (.I(U_in[498]), .O(U_in_c_498));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_499 (.I(U_in[499]), .O(U_in_c_499));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_500 (.I(U_in[500]), .O(U_in_c_500));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_501 (.I(U_in[501]), .O(U_in_c_501));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_502 (.I(U_in[502]), .O(U_in_c_502));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_503 (.I(U_in[503]), .O(U_in_c_503));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_504 (.I(U_in[504]), .O(U_in_c_504));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    CCU2C add_7640_19 (.A0(n4205), .B0(n30938), .C0(n64_adj_578), .D0(n3057), 
          .A1(n4204), .B1(n30938), .C1(n64_adj_578), .D1(n3479), .CIN(n32680), 
          .COUT(n32681), .S0(n4322), .S1(n4321));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_19.INIT0 = 16'ha9aa;
    defparam add_7640_19.INIT1 = 16'ha9aa;
    defparam add_7640_19.INJECT1_0 = "NO";
    defparam add_7640_19.INJECT1_1 = "NO";
    CCU2C add_7640_17 (.A0(n4207), .B0(n30938), .C0(n64_adj_578), .D0(n2762), 
          .A1(n4206), .B1(n30938), .C1(n64_adj_578), .D1(n2911), .CIN(n32679), 
          .COUT(n32680), .S0(n4324), .S1(n4323));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_17.INIT0 = 16'ha9aa;
    defparam add_7640_17.INIT1 = 16'ha9aa;
    defparam add_7640_17.INJECT1_0 = "NO";
    defparam add_7640_17.INJECT1_1 = "NO";
    CCU2C add_7640_15 (.A0(n4209), .B0(n30938), .C0(n64_adj_578), .D0(n2455), 
          .A1(n4208), .B1(n30938), .C1(n64_adj_578), .D1(n3060), .CIN(n32678), 
          .COUT(n32679), .S0(n4326), .S1(n4325));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_15.INIT0 = 16'ha9aa;
    defparam add_7640_15.INIT1 = 16'ha9aa;
    defparam add_7640_15.INJECT1_0 = "NO";
    defparam add_7640_15.INJECT1_1 = "NO";
    CCU2C add_7640_13 (.A0(n4211), .B0(n30938), .C0(n64_adj_578), .D0(n2298), 
          .A1(n4210), .B1(n30938), .C1(n64_adj_578), .D1(n2456), .CIN(n32677), 
          .COUT(n32678), .S0(n4328), .S1(n4327));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_13.INIT0 = 16'ha9aa;
    defparam add_7640_13.INIT1 = 16'ha9aa;
    defparam add_7640_13.INJECT1_0 = "NO";
    defparam add_7640_13.INJECT1_1 = "NO";
    CCU2C add_7640_11 (.A0(n4213), .B0(n30938), .C0(n64_adj_578), .D0(n1805), 
          .A1(n4212), .B1(n30938), .C1(n64_adj_578), .D1(n2137), .CIN(n32676), 
          .COUT(n32677), .S0(n4330), .S1(n4329));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_11.INIT0 = 16'ha9aa;
    defparam add_7640_11.INIT1 = 16'ha9aa;
    defparam add_7640_11.INJECT1_0 = "NO";
    defparam add_7640_11.INJECT1_1 = "NO";
    CCU2C add_7640_9 (.A0(n4215), .B0(n30938), .C0(n64_adj_578), .D0(n1462), 
          .A1(n4214), .B1(n30938), .C1(n64_adj_578), .D1(n1635), .CIN(n32675), 
          .COUT(n32676), .S0(n4332), .S1(n4331));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_9.INIT0 = 16'ha9aa;
    defparam add_7640_9.INIT1 = 16'ha9aa;
    defparam add_7640_9.INJECT1_0 = "NO";
    defparam add_7640_9.INJECT1_1 = "NO";
    CCU2C add_7640_7 (.A0(n4217), .B0(n30938), .C0(n64_adj_578), .D0(n2142), 
          .A1(n4216), .B1(n30938), .C1(n64_adj_578), .D1(n2141), .CIN(n32674), 
          .COUT(n32675), .S0(n4334), .S1(n4333));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_7.INIT0 = 16'ha9aa;
    defparam add_7640_7.INIT1 = 16'ha9aa;
    defparam add_7640_7.INJECT1_0 = "NO";
    defparam add_7640_7.INJECT1_1 = "NO";
    CCU2C add_7640_5 (.A0(n4219), .B0(n30938), .C0(n64_adj_578), .D0(n42824), 
          .A1(n4218), .B1(n30938), .C1(n64_adj_578), .D1(n42822), .CIN(n32673), 
          .COUT(n32674), .S0(n4336), .S1(n4335));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_5.INIT0 = 16'ha9aa;
    defparam add_7640_5.INIT1 = 16'ha9aa;
    defparam add_7640_5.INJECT1_0 = "NO";
    defparam add_7640_5.INJECT1_1 = "NO";
    CCU2C add_7640_3 (.A0(n888), .B0(n30938), .C0(n64_adj_578), .D0(n42827), 
          .A1(n4220), .B1(n30938), .C1(n64_adj_578), .D1(n42823), .CIN(n32672), 
          .COUT(n32673), .S0(n4338), .S1(n4337));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_3.INIT0 = 16'ha9aa;
    defparam add_7640_3.INIT1 = 16'ha9aa;
    defparam add_7640_3.INJECT1_0 = "NO";
    defparam add_7640_3.INJECT1_1 = "NO";
    CCU2C add_7640_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_578), .B1(n30938), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32672));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7640_1.INIT0 = 16'h0000;
    defparam add_7640_1.INIT1 = 16'heee1;
    defparam add_7640_1.INJECT1_0 = "NO";
    defparam add_7640_1.INJECT1_1 = "NO";
    CCU2C add_7639_27 (.A0(n4076), .B0(n42790), .C0(n64_adj_549), .D0(n4117), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32668), 
          .S0(n4196));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_27.INIT0 = 16'ha9aa;
    defparam add_7639_27.INIT1 = 16'h0000;
    defparam add_7639_27.INJECT1_0 = "NO";
    defparam add_7639_27.INJECT1_1 = "NO";
    CCU2C add_7639_25 (.A0(n4078), .B0(n42790), .C0(n64_adj_549), .D0(n3870), 
          .A1(n4077), .B1(n42790), .C1(n64_adj_549), .D1(n3995), .CIN(n32667), 
          .COUT(n32668), .S0(n4198), .S1(n4197));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_25.INIT0 = 16'ha9aa;
    defparam add_7639_25.INIT1 = 16'ha9aa;
    defparam add_7639_25.INJECT1_0 = "NO";
    defparam add_7639_25.INJECT1_1 = "NO";
    CCU2C add_7639_23 (.A0(n4080), .B0(n42790), .C0(n64_adj_549), .D0(n3611), 
          .A1(n4079), .B1(n42790), .C1(n64_adj_549), .D1(n3871), .CIN(n32666), 
          .COUT(n32667), .S0(n4200), .S1(n4199));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_23.INIT0 = 16'ha9aa;
    defparam add_7639_23.INIT1 = 16'ha9aa;
    defparam add_7639_23.INJECT1_0 = "NO";
    defparam add_7639_23.INJECT1_1 = "NO";
    CCU2C add_7639_21 (.A0(n4082), .B0(n42790), .C0(n64_adj_549), .D0(n3340), 
          .A1(n4081), .B1(n42790), .C1(n64_adj_549), .D1(n3477), .CIN(n32665), 
          .COUT(n32666), .S0(n4202), .S1(n4201));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_21.INIT0 = 16'ha9aa;
    defparam add_7639_21.INIT1 = 16'ha9aa;
    defparam add_7639_21.INJECT1_0 = "NO";
    defparam add_7639_21.INJECT1_1 = "NO";
    CCU2C add_7639_19 (.A0(n4084), .B0(n42790), .C0(n64_adj_549), .D0(n3057), 
          .A1(n4083), .B1(n42790), .C1(n64_adj_549), .D1(n3479), .CIN(n32664), 
          .COUT(n32665), .S0(n4204), .S1(n4203));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_19.INIT0 = 16'ha9aa;
    defparam add_7639_19.INIT1 = 16'ha9aa;
    defparam add_7639_19.INJECT1_0 = "NO";
    defparam add_7639_19.INJECT1_1 = "NO";
    CCU2C add_7639_17 (.A0(n4086), .B0(n42790), .C0(n64_adj_549), .D0(n2762), 
          .A1(n4085), .B1(n42790), .C1(n64_adj_549), .D1(n2911), .CIN(n32663), 
          .COUT(n32664), .S0(n4206), .S1(n4205));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_17.INIT0 = 16'ha9aa;
    defparam add_7639_17.INIT1 = 16'ha9aa;
    defparam add_7639_17.INJECT1_0 = "NO";
    defparam add_7639_17.INJECT1_1 = "NO";
    CCU2C add_7639_15 (.A0(n4088), .B0(n42790), .C0(n64_adj_549), .D0(n2455), 
          .A1(n4087), .B1(n42790), .C1(n64_adj_549), .D1(n3060), .CIN(n32662), 
          .COUT(n32663), .S0(n4208), .S1(n4207));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_15.INIT0 = 16'ha9aa;
    defparam add_7639_15.INIT1 = 16'ha9aa;
    defparam add_7639_15.INJECT1_0 = "NO";
    defparam add_7639_15.INJECT1_1 = "NO";
    CCU2C add_7639_13 (.A0(n4090), .B0(n42790), .C0(n64_adj_549), .D0(n2298), 
          .A1(n4089), .B1(n42790), .C1(n64_adj_549), .D1(n2456), .CIN(n32661), 
          .COUT(n32662), .S0(n4210), .S1(n4209));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_13.INIT0 = 16'ha9aa;
    defparam add_7639_13.INIT1 = 16'ha9aa;
    defparam add_7639_13.INJECT1_0 = "NO";
    defparam add_7639_13.INJECT1_1 = "NO";
    CCU2C add_7639_11 (.A0(n4092), .B0(n42790), .C0(n64_adj_549), .D0(n1805), 
          .A1(n4091), .B1(n42790), .C1(n64_adj_549), .D1(n2137), .CIN(n32660), 
          .COUT(n32661), .S0(n4212), .S1(n4211));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_11.INIT0 = 16'ha9aa;
    defparam add_7639_11.INIT1 = 16'ha9aa;
    defparam add_7639_11.INJECT1_0 = "NO";
    defparam add_7639_11.INJECT1_1 = "NO";
    PFUMX div_4016_LessThan_2058_i58 (.BLUT(n38_adj_365), .ALUT(n40_adj_366), 
          .C0(n37965), .Z(n58_adj_375));
    LUT4 i24284_4_lut (.A(n42463), .B(n42462), .C(n11_adj_707), .D(n39535), 
         .Z(n39544)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24284_4_lut.init = 16'h1011;
    LUT4 i1_4_lut_adj_50 (.A(n163_adj_155), .B(i[0]), .C(done_N_1932), 
         .D(n13381), .Z(n30843)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i1_4_lut_adj_50.init = 16'heca0;
    LUT4 i1_2_lut_adj_51 (.A(done_N_1929), .B(done_N_1934), .Z(n13381)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i1_2_lut_adj_51.init = 16'heeee;
    LUT4 div_4016_LessThan_2513_i33_2_lut (.A(n3842), .B(n125_adj_230), 
         .Z(n33_adj_476)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i33_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i22_3_lut_3_lut (.A(n4664), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n22_adj_680)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i22_3_lut_3_lut.init = 16'hd4d4;
    IB U_in_pad_505 (.I(U_in[505]), .O(U_in_c_505));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_506 (.I(U_in[506]), .O(U_in_c_506));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_507 (.I(U_in[507]), .O(U_in_c_507));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_508 (.I(U_in[508]), .O(U_in_c_508));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_509 (.I(U_in[509]), .O(U_in_c_509));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_510 (.I(U_in[510]), .O(U_in_c_510));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_511 (.I(U_in[511]), .O(U_in_c_511));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB start_pad (.I(start), .O(start_c));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(7[24:29])
    IB rst_pad (.I(rst), .O(rst_c));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    IB clk_pad (.I(clk), .O(clk_c));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(5[24:27])
    OB x_out_pad_0 (.I(x_out_c_0), .O(x_out[0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7639_9 (.A0(n4094), .B0(n42790), .C0(n64_adj_549), .D0(n1462), 
          .A1(n4093), .B1(n42790), .C1(n64_adj_549), .D1(n1635), .CIN(n32659), 
          .COUT(n32660), .S0(n4214), .S1(n4213));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_9.INIT0 = 16'ha9aa;
    defparam add_7639_9.INIT1 = 16'ha9aa;
    defparam add_7639_9.INJECT1_0 = "NO";
    defparam add_7639_9.INJECT1_1 = "NO";
    CCU2C add_7639_7 (.A0(n4096), .B0(n42790), .C0(n64_adj_549), .D0(n2142), 
          .A1(n4095), .B1(n42790), .C1(n64_adj_549), .D1(n2141), .CIN(n32658), 
          .COUT(n32659), .S0(n4216), .S1(n4215));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_7.INIT0 = 16'ha9aa;
    defparam add_7639_7.INIT1 = 16'ha9aa;
    defparam add_7639_7.INJECT1_0 = "NO";
    defparam add_7639_7.INJECT1_1 = "NO";
    CCU2C add_7639_5 (.A0(n4098), .B0(n42790), .C0(n64_adj_549), .D0(n42824), 
          .A1(n4097), .B1(n42790), .C1(n64_adj_549), .D1(n42822), .CIN(n32657), 
          .COUT(n32658), .S0(n4218), .S1(n4217));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_5.INIT0 = 16'ha9aa;
    defparam add_7639_5.INIT1 = 16'ha9aa;
    defparam add_7639_5.INJECT1_0 = "NO";
    defparam add_7639_5.INJECT1_1 = "NO";
    CCU2C add_7639_3 (.A0(n887), .B0(n42790), .C0(n64_adj_549), .D0(n42827), 
          .A1(n4099), .B1(n42790), .C1(n64_adj_549), .D1(n42823), .CIN(n32656), 
          .COUT(n32657), .S0(n4220), .S1(n4219));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_3.INIT0 = 16'ha9aa;
    defparam add_7639_3.INIT1 = 16'ha9aa;
    defparam add_7639_3.INJECT1_0 = "NO";
    defparam add_7639_3.INJECT1_1 = "NO";
    CCU2C add_7639_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_549), .B1(n42790), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32656));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7639_1.INIT0 = 16'h0000;
    defparam add_7639_1.INIT1 = 16'heee1;
    defparam add_7639_1.INJECT1_0 = "NO";
    defparam add_7639_1.INJECT1_1 = "NO";
    CCU2C add_7638_25 (.A0(n3954), .B0(n30932), .C0(n64_adj_520), .D0(n3870), 
          .A1(n3953), .B1(n30932), .C1(n64_adj_520), .D1(n3995), .CIN(n32651), 
          .S0(n4077), .S1(n4076));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_25.INIT0 = 16'ha9aa;
    defparam add_7638_25.INIT1 = 16'ha9aa;
    defparam add_7638_25.INJECT1_0 = "NO";
    defparam add_7638_25.INJECT1_1 = "NO";
    CCU2C add_7638_23 (.A0(n3956), .B0(n30932), .C0(n64_adj_520), .D0(n3611), 
          .A1(n3955), .B1(n30932), .C1(n64_adj_520), .D1(n3871), .CIN(n32650), 
          .COUT(n32651), .S0(n4079), .S1(n4078));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_23.INIT0 = 16'ha9aa;
    defparam add_7638_23.INIT1 = 16'ha9aa;
    defparam add_7638_23.INJECT1_0 = "NO";
    defparam add_7638_23.INJECT1_1 = "NO";
    CCU2C add_7638_21 (.A0(n3958), .B0(n30932), .C0(n64_adj_520), .D0(n3340), 
          .A1(n3957), .B1(n30932), .C1(n64_adj_520), .D1(n3477), .CIN(n32649), 
          .COUT(n32650), .S0(n4081), .S1(n4080));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_21.INIT0 = 16'ha9aa;
    defparam add_7638_21.INIT1 = 16'ha9aa;
    defparam add_7638_21.INJECT1_0 = "NO";
    defparam add_7638_21.INJECT1_1 = "NO";
    CCU2C add_7638_19 (.A0(n3960), .B0(n30932), .C0(n64_adj_520), .D0(n3057), 
          .A1(n3959), .B1(n30932), .C1(n64_adj_520), .D1(n3479), .CIN(n32648), 
          .COUT(n32649), .S0(n4083), .S1(n4082));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_19.INIT0 = 16'ha9aa;
    defparam add_7638_19.INIT1 = 16'ha9aa;
    defparam add_7638_19.INJECT1_0 = "NO";
    defparam add_7638_19.INJECT1_1 = "NO";
    CCU2C add_7638_17 (.A0(n3962), .B0(n30932), .C0(n64_adj_520), .D0(n2762), 
          .A1(n3961), .B1(n30932), .C1(n64_adj_520), .D1(n2911), .CIN(n32647), 
          .COUT(n32648), .S0(n4085), .S1(n4084));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_17.INIT0 = 16'ha9aa;
    defparam add_7638_17.INIT1 = 16'ha9aa;
    defparam add_7638_17.INJECT1_0 = "NO";
    defparam add_7638_17.INJECT1_1 = "NO";
    CCU2C add_7638_15 (.A0(n3964), .B0(n30932), .C0(n64_adj_520), .D0(n2455), 
          .A1(n3963), .B1(n30932), .C1(n64_adj_520), .D1(n3060), .CIN(n32646), 
          .COUT(n32647), .S0(n4087), .S1(n4086));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_15.INIT0 = 16'ha9aa;
    defparam add_7638_15.INIT1 = 16'ha9aa;
    defparam add_7638_15.INJECT1_0 = "NO";
    defparam add_7638_15.INJECT1_1 = "NO";
    CCU2C add_7638_13 (.A0(n3966), .B0(n30932), .C0(n64_adj_520), .D0(n2298), 
          .A1(n3965), .B1(n30932), .C1(n64_adj_520), .D1(n2456), .CIN(n32645), 
          .COUT(n32646), .S0(n4089), .S1(n4088));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_13.INIT0 = 16'ha9aa;
    defparam add_7638_13.INIT1 = 16'ha9aa;
    defparam add_7638_13.INJECT1_0 = "NO";
    defparam add_7638_13.INJECT1_1 = "NO";
    CCU2C add_7638_11 (.A0(n3968), .B0(n30932), .C0(n64_adj_520), .D0(n1805), 
          .A1(n3967), .B1(n30932), .C1(n64_adj_520), .D1(n2137), .CIN(n32644), 
          .COUT(n32645), .S0(n4091), .S1(n4090));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_11.INIT0 = 16'ha9aa;
    defparam add_7638_11.INIT1 = 16'ha9aa;
    defparam add_7638_11.INJECT1_0 = "NO";
    defparam add_7638_11.INJECT1_1 = "NO";
    CCU2C add_7638_9 (.A0(n3970), .B0(n30932), .C0(n64_adj_520), .D0(n1462), 
          .A1(n3969), .B1(n30932), .C1(n64_adj_520), .D1(n1635), .CIN(n32643), 
          .COUT(n32644), .S0(n4093), .S1(n4092));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_9.INIT0 = 16'ha9aa;
    defparam add_7638_9.INIT1 = 16'ha9aa;
    defparam add_7638_9.INJECT1_0 = "NO";
    defparam add_7638_9.INJECT1_1 = "NO";
    CCU2C add_7638_7 (.A0(n3972), .B0(n30932), .C0(n64_adj_520), .D0(n2142), 
          .A1(n3971), .B1(n30932), .C1(n64_adj_520), .D1(n2141), .CIN(n32642), 
          .COUT(n32643), .S0(n4095), .S1(n4094));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_7.INIT0 = 16'ha9aa;
    defparam add_7638_7.INIT1 = 16'ha9aa;
    defparam add_7638_7.INJECT1_0 = "NO";
    defparam add_7638_7.INJECT1_1 = "NO";
    CCU2C add_7638_5 (.A0(n3974), .B0(n30932), .C0(n64_adj_520), .D0(n42824), 
          .A1(n3973), .B1(n30932), .C1(n64_adj_520), .D1(n42822), .CIN(n32641), 
          .COUT(n32642), .S0(n4097), .S1(n4096));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_5.INIT0 = 16'ha9aa;
    defparam add_7638_5.INIT1 = 16'ha9aa;
    defparam add_7638_5.INJECT1_0 = "NO";
    defparam add_7638_5.INJECT1_1 = "NO";
    CCU2C add_7638_3 (.A0(n886), .B0(n30932), .C0(n64_adj_520), .D0(n42827), 
          .A1(n3975), .B1(n30932), .C1(n64_adj_520), .D1(n42823), .CIN(n32640), 
          .COUT(n32641), .S0(n4099), .S1(n4098));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_3.INIT0 = 16'ha9aa;
    defparam add_7638_3.INIT1 = 16'ha9aa;
    defparam add_7638_3.INJECT1_0 = "NO";
    defparam add_7638_3.INJECT1_1 = "NO";
    CCU2C add_7638_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_520), .B1(n30932), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32640));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7638_1.INIT0 = 16'h0000;
    defparam add_7638_1.INIT1 = 16'heee1;
    defparam add_7638_1.INJECT1_0 = "NO";
    defparam add_7638_1.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_2513_i47_2_lut_rep_911 (.A(n3835), .B(n118_adj_225), 
         .Z(n42610)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i47_2_lut_rep_911.init = 16'h6666;
    PFUMX div_4016_LessThan_2058_i52 (.BLUT(n44_adj_368), .ALUT(n50_adj_371), 
          .C0(n37932), .Z(n52_adj_372));
    LUT4 div_4016_LessThan_2513_i32_3_lut_3_lut (.A(n3835), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n32_adj_475)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i32_3_lut_3_lut.init = 16'hd4d4;
    OB x_out_pad_1 (.I(x_out_c_1), .O(x_out[1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_2 (.I(x_out_c_2), .O(x_out[2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_3 (.I(x_out_c_3), .O(x_out[3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_4 (.I(x_out_c_4), .O(x_out[4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_5 (.I(x_out_c_5), .O(x_out[5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_6 (.I(x_out_c_6), .O(x_out[6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_7 (.I(x_out_c_7), .O(x_out[7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_8 (.I(x_out_c_8), .O(x_out[8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_9 (.I(x_out_c_9), .O(x_out[9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_10 (.I(x_out_c_10), .O(x_out[10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7637_25 (.A0(n3827), .B0(n30929), .C0(n64_adj_493), .D0(n3870), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32636), 
          .S0(n3953));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_25.INIT0 = 16'ha9aa;
    defparam add_7637_25.INIT1 = 16'h0000;
    defparam add_7637_25.INJECT1_0 = "NO";
    defparam add_7637_25.INJECT1_1 = "NO";
    CCU2C add_7637_23 (.A0(n3829), .B0(n30929), .C0(n64_adj_493), .D0(n3611), 
          .A1(n3828), .B1(n30929), .C1(n64_adj_493), .D1(n3871), .CIN(n32635), 
          .COUT(n32636), .S0(n3955), .S1(n3954));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_23.INIT0 = 16'ha9aa;
    defparam add_7637_23.INIT1 = 16'ha9aa;
    defparam add_7637_23.INJECT1_0 = "NO";
    defparam add_7637_23.INJECT1_1 = "NO";
    CCU2C add_7637_21 (.A0(n3831), .B0(n30929), .C0(n64_adj_493), .D0(n3340), 
          .A1(n3830), .B1(n30929), .C1(n64_adj_493), .D1(n3477), .CIN(n32634), 
          .COUT(n32635), .S0(n3957), .S1(n3956));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_21.INIT0 = 16'ha9aa;
    defparam add_7637_21.INIT1 = 16'ha9aa;
    defparam add_7637_21.INJECT1_0 = "NO";
    defparam add_7637_21.INJECT1_1 = "NO";
    CCU2C add_7637_19 (.A0(n3833), .B0(n30929), .C0(n64_adj_493), .D0(n3057), 
          .A1(n3832), .B1(n30929), .C1(n64_adj_493), .D1(n3479), .CIN(n32633), 
          .COUT(n32634), .S0(n3959), .S1(n3958));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_19.INIT0 = 16'ha9aa;
    defparam add_7637_19.INIT1 = 16'ha9aa;
    defparam add_7637_19.INJECT1_0 = "NO";
    defparam add_7637_19.INJECT1_1 = "NO";
    CCU2C add_7637_17 (.A0(n3835), .B0(n30929), .C0(n64_adj_493), .D0(n2762), 
          .A1(n3834), .B1(n30929), .C1(n64_adj_493), .D1(n2911), .CIN(n32632), 
          .COUT(n32633), .S0(n3961), .S1(n3960));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_17.INIT0 = 16'ha9aa;
    defparam add_7637_17.INIT1 = 16'ha9aa;
    defparam add_7637_17.INJECT1_0 = "NO";
    defparam add_7637_17.INJECT1_1 = "NO";
    CCU2C add_7637_15 (.A0(n3837), .B0(n30929), .C0(n64_adj_493), .D0(n2455), 
          .A1(n3836), .B1(n30929), .C1(n64_adj_493), .D1(n3060), .CIN(n32631), 
          .COUT(n32632), .S0(n3963), .S1(n3962));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_15.INIT0 = 16'ha9aa;
    defparam add_7637_15.INIT1 = 16'ha9aa;
    defparam add_7637_15.INJECT1_0 = "NO";
    defparam add_7637_15.INJECT1_1 = "NO";
    CCU2C add_7637_13 (.A0(n3839), .B0(n30929), .C0(n64_adj_493), .D0(n2298), 
          .A1(n3838), .B1(n30929), .C1(n64_adj_493), .D1(n2456), .CIN(n32630), 
          .COUT(n32631), .S0(n3965), .S1(n3964));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_13.INIT0 = 16'ha9aa;
    defparam add_7637_13.INIT1 = 16'ha9aa;
    defparam add_7637_13.INJECT1_0 = "NO";
    defparam add_7637_13.INJECT1_1 = "NO";
    CCU2C add_7637_11 (.A0(n3841), .B0(n30929), .C0(n64_adj_493), .D0(n1805), 
          .A1(n3840), .B1(n30929), .C1(n64_adj_493), .D1(n2137), .CIN(n32629), 
          .COUT(n32630), .S0(n3967), .S1(n3966));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_11.INIT0 = 16'ha9aa;
    defparam add_7637_11.INIT1 = 16'ha9aa;
    defparam add_7637_11.INJECT1_0 = "NO";
    defparam add_7637_11.INJECT1_1 = "NO";
    CCU2C add_7637_9 (.A0(n3843), .B0(n30929), .C0(n64_adj_493), .D0(n1462), 
          .A1(n3842), .B1(n30929), .C1(n64_adj_493), .D1(n1635), .CIN(n32628), 
          .COUT(n32629), .S0(n3969), .S1(n3968));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_9.INIT0 = 16'ha9aa;
    defparam add_7637_9.INIT1 = 16'ha9aa;
    defparam add_7637_9.INJECT1_0 = "NO";
    defparam add_7637_9.INJECT1_1 = "NO";
    CCU2C add_7637_7 (.A0(n3845), .B0(n30929), .C0(n64_adj_493), .D0(n2142), 
          .A1(n3844), .B1(n30929), .C1(n64_adj_493), .D1(n2141), .CIN(n32627), 
          .COUT(n32628), .S0(n3971), .S1(n3970));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_7.INIT0 = 16'ha9aa;
    defparam add_7637_7.INIT1 = 16'ha9aa;
    defparam add_7637_7.INJECT1_0 = "NO";
    defparam add_7637_7.INJECT1_1 = "NO";
    CCU2C add_7637_5 (.A0(n3847), .B0(n30929), .C0(n64_adj_493), .D0(n42824), 
          .A1(n3846), .B1(n30929), .C1(n64_adj_493), .D1(n42822), .CIN(n32626), 
          .COUT(n32627), .S0(n3973), .S1(n3972));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_5.INIT0 = 16'ha9aa;
    defparam add_7637_5.INIT1 = 16'ha9aa;
    defparam add_7637_5.INJECT1_0 = "NO";
    defparam add_7637_5.INJECT1_1 = "NO";
    CCU2C add_7637_3 (.A0(n885), .B0(n30929), .C0(n64_adj_493), .D0(n42827), 
          .A1(n3848), .B1(n30929), .C1(n64_adj_493), .D1(n42823), .CIN(n32625), 
          .COUT(n32626), .S0(n3975), .S1(n3974));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_3.INIT0 = 16'ha9aa;
    defparam add_7637_3.INIT1 = 16'ha9aa;
    defparam add_7637_3.INJECT1_0 = "NO";
    defparam add_7637_3.INJECT1_1 = "NO";
    CCU2C add_7637_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_493), .B1(n30929), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32625));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7637_1.INIT0 = 16'h0000;
    defparam add_7637_1.INIT1 = 16'heee1;
    defparam add_7637_1.INJECT1_0 = "NO";
    defparam add_7637_1.INJECT1_1 = "NO";
    CCU2C add_7636_23 (.A0(n3699), .B0(n30926), .C0(n64_adj_469), .D0(n3611), 
          .A1(n3698), .B1(n30926), .C1(n64_adj_469), .D1(n3871), .CIN(n32620), 
          .S0(n3828), .S1(n3827));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_23.INIT0 = 16'ha9aa;
    defparam add_7636_23.INIT1 = 16'ha9aa;
    defparam add_7636_23.INJECT1_0 = "NO";
    defparam add_7636_23.INJECT1_1 = "NO";
    CCU2C add_7636_21 (.A0(n3701), .B0(n30926), .C0(n64_adj_469), .D0(n3340), 
          .A1(n3700), .B1(n30926), .C1(n64_adj_469), .D1(n3477), .CIN(n32619), 
          .COUT(n32620), .S0(n3830), .S1(n3829));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_21.INIT0 = 16'ha9aa;
    defparam add_7636_21.INIT1 = 16'ha9aa;
    defparam add_7636_21.INJECT1_0 = "NO";
    defparam add_7636_21.INJECT1_1 = "NO";
    CCU2C add_7636_19 (.A0(n3703), .B0(n30926), .C0(n64_adj_469), .D0(n3057), 
          .A1(n3702), .B1(n30926), .C1(n64_adj_469), .D1(n3479), .CIN(n32618), 
          .COUT(n32619), .S0(n3832), .S1(n3831));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_19.INIT0 = 16'ha9aa;
    defparam add_7636_19.INIT1 = 16'ha9aa;
    defparam add_7636_19.INJECT1_0 = "NO";
    defparam add_7636_19.INJECT1_1 = "NO";
    CCU2C add_7636_17 (.A0(n3705), .B0(n30926), .C0(n64_adj_469), .D0(n2762), 
          .A1(n3704), .B1(n30926), .C1(n64_adj_469), .D1(n2911), .CIN(n32617), 
          .COUT(n32618), .S0(n3834), .S1(n3833));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_17.INIT0 = 16'ha9aa;
    defparam add_7636_17.INIT1 = 16'ha9aa;
    defparam add_7636_17.INJECT1_0 = "NO";
    defparam add_7636_17.INJECT1_1 = "NO";
    CCU2C add_7636_15 (.A0(n3707), .B0(n30926), .C0(n64_adj_469), .D0(n2455), 
          .A1(n3706), .B1(n30926), .C1(n64_adj_469), .D1(n3060), .CIN(n32616), 
          .COUT(n32617), .S0(n3836), .S1(n3835));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_15.INIT0 = 16'ha9aa;
    defparam add_7636_15.INIT1 = 16'ha9aa;
    defparam add_7636_15.INJECT1_0 = "NO";
    defparam add_7636_15.INJECT1_1 = "NO";
    CCU2C add_7636_13 (.A0(n3709), .B0(n30926), .C0(n64_adj_469), .D0(n2298), 
          .A1(n3708), .B1(n30926), .C1(n64_adj_469), .D1(n2456), .CIN(n32615), 
          .COUT(n32616), .S0(n3838), .S1(n3837));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_13.INIT0 = 16'ha9aa;
    defparam add_7636_13.INIT1 = 16'ha9aa;
    defparam add_7636_13.INJECT1_0 = "NO";
    defparam add_7636_13.INJECT1_1 = "NO";
    CCU2C add_7636_11 (.A0(n3711), .B0(n30926), .C0(n64_adj_469), .D0(n1805), 
          .A1(n3710), .B1(n30926), .C1(n64_adj_469), .D1(n2137), .CIN(n32614), 
          .COUT(n32615), .S0(n3840), .S1(n3839));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_11.INIT0 = 16'ha9aa;
    defparam add_7636_11.INIT1 = 16'ha9aa;
    defparam add_7636_11.INJECT1_0 = "NO";
    defparam add_7636_11.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_3066_i29_2_lut_rep_782 (.A(n4663), .B(n120), 
         .Z(n42481)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i29_2_lut_rep_782.init = 16'h6666;
    LUT4 div_4016_LessThan_2513_i43_2_lut_rep_912 (.A(n3837), .B(n120), 
         .Z(n42611)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i43_2_lut_rep_912.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(n111), .B(n110_adj_220), .C(n42814), 
         .D(n42813), .Z(n36926)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'hfffe;
    FD1P3JX i_i0_i1 (.D(n30845), .SP(clk_c_enable_831), .PD(clk_c_enable_708), 
            .CK(clk_c), .Q(i[1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i_i0_i1.GSR = "ENABLED";
    FD1P3IX x_3___i2 (.D(n5524), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i2.GSR = "ENABLED";
    FD1P3IX x_3___i3 (.D(n5523), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i3.GSR = "ENABLED";
    FD1P3IX x_3___i4 (.D(n5522), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i4.GSR = "ENABLED";
    FD1P3IX x_3___i5 (.D(n5521), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i5.GSR = "ENABLED";
    FD1P3IX x_3___i6 (.D(n5520), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i6.GSR = "ENABLED";
    OB x_out_pad_11 (.I(x_out_c_11), .O(x_out[11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_12 (.I(x_out_c_12), .O(x_out[12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_13 (.I(x_out_c_13), .O(x_out[13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_14 (.I(x_out_c_14), .O(x_out[14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_15 (.I(x_out_c_15), .O(x_out[15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_16 (.I(x_out_c_16), .O(x_out[16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_17 (.I(x_out_c_17), .O(x_out[17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_18 (.I(x_out_c_18), .O(x_out[18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_19 (.I(x_out_c_19), .O(x_out[19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7636_9 (.A0(n3713), .B0(n30926), .C0(n64_adj_469), .D0(n1462), 
          .A1(n3712), .B1(n30926), .C1(n64_adj_469), .D1(n1635), .CIN(n32613), 
          .COUT(n32614), .S0(n3842), .S1(n3841));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_9.INIT0 = 16'ha9aa;
    defparam add_7636_9.INIT1 = 16'ha9aa;
    defparam add_7636_9.INJECT1_0 = "NO";
    defparam add_7636_9.INJECT1_1 = "NO";
    CCU2C add_7636_7 (.A0(n3715), .B0(n30926), .C0(n64_adj_469), .D0(n2142), 
          .A1(n3714), .B1(n30926), .C1(n64_adj_469), .D1(n2141), .CIN(n32612), 
          .COUT(n32613), .S0(n3844), .S1(n3843));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_7.INIT0 = 16'ha9aa;
    defparam add_7636_7.INIT1 = 16'ha9aa;
    defparam add_7636_7.INJECT1_0 = "NO";
    defparam add_7636_7.INJECT1_1 = "NO";
    CCU2C add_7636_5 (.A0(n3717), .B0(n30926), .C0(n64_adj_469), .D0(n42824), 
          .A1(n3716), .B1(n30926), .C1(n64_adj_469), .D1(n42822), .CIN(n32611), 
          .COUT(n32612), .S0(n3846), .S1(n3845));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_5.INIT0 = 16'ha9aa;
    defparam add_7636_5.INIT1 = 16'ha9aa;
    defparam add_7636_5.INJECT1_0 = "NO";
    defparam add_7636_5.INJECT1_1 = "NO";
    CCU2C add_7636_3 (.A0(n884), .B0(n30926), .C0(n64_adj_469), .D0(n42827), 
          .A1(n3718), .B1(n30926), .C1(n64_adj_469), .D1(n42823), .CIN(n32610), 
          .COUT(n32611), .S0(n3848), .S1(n3847));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_3.INIT0 = 16'ha9aa;
    defparam add_7636_3.INIT1 = 16'ha9aa;
    defparam add_7636_3.INJECT1_0 = "NO";
    defparam add_7636_3.INJECT1_1 = "NO";
    CCU2C add_7636_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_469), .B1(n30926), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32610));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7636_1.INIT0 = 16'h0000;
    defparam add_7636_1.INIT1 = 16'heee1;
    defparam add_7636_1.INJECT1_0 = "NO";
    defparam add_7636_1.INJECT1_1 = "NO";
    CCU2C add_7635_23 (.A0(n3566), .B0(n30923), .C0(n64_adj_444), .D0(n3611), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32606), 
          .S0(n3698));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_23.INIT0 = 16'ha9aa;
    defparam add_7635_23.INIT1 = 16'h0000;
    defparam add_7635_23.INJECT1_0 = "NO";
    defparam add_7635_23.INJECT1_1 = "NO";
    CCU2C add_7635_21 (.A0(n3568), .B0(n30923), .C0(n64_adj_444), .D0(n3340), 
          .A1(n3567), .B1(n30923), .C1(n64_adj_444), .D1(n3477), .CIN(n32605), 
          .COUT(n32606), .S0(n3700), .S1(n3699));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_21.INIT0 = 16'ha9aa;
    defparam add_7635_21.INIT1 = 16'ha9aa;
    defparam add_7635_21.INJECT1_0 = "NO";
    defparam add_7635_21.INJECT1_1 = "NO";
    CCU2C add_7635_19 (.A0(n3570), .B0(n30923), .C0(n64_adj_444), .D0(n3057), 
          .A1(n3569), .B1(n30923), .C1(n64_adj_444), .D1(n3479), .CIN(n32604), 
          .COUT(n32605), .S0(n3702), .S1(n3701));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_19.INIT0 = 16'ha9aa;
    defparam add_7635_19.INIT1 = 16'ha9aa;
    defparam add_7635_19.INJECT1_0 = "NO";
    defparam add_7635_19.INJECT1_1 = "NO";
    CCU2C add_7635_17 (.A0(n3572), .B0(n30923), .C0(n64_adj_444), .D0(n2762), 
          .A1(n3571), .B1(n30923), .C1(n64_adj_444), .D1(n2911), .CIN(n32603), 
          .COUT(n32604), .S0(n3704), .S1(n3703));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_17.INIT0 = 16'ha9aa;
    defparam add_7635_17.INIT1 = 16'ha9aa;
    defparam add_7635_17.INJECT1_0 = "NO";
    defparam add_7635_17.INJECT1_1 = "NO";
    CCU2C add_7635_15 (.A0(n3574), .B0(n30923), .C0(n64_adj_444), .D0(n2455), 
          .A1(n3573), .B1(n30923), .C1(n64_adj_444), .D1(n3060), .CIN(n32602), 
          .COUT(n32603), .S0(n3706), .S1(n3705));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_15.INIT0 = 16'ha9aa;
    defparam add_7635_15.INIT1 = 16'ha9aa;
    defparam add_7635_15.INJECT1_0 = "NO";
    defparam add_7635_15.INJECT1_1 = "NO";
    CCU2C add_7635_13 (.A0(n3576), .B0(n30923), .C0(n64_adj_444), .D0(n2298), 
          .A1(n3575), .B1(n30923), .C1(n64_adj_444), .D1(n2456), .CIN(n32601), 
          .COUT(n32602), .S0(n3708), .S1(n3707));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_13.INIT0 = 16'ha9aa;
    defparam add_7635_13.INIT1 = 16'ha9aa;
    defparam add_7635_13.INJECT1_0 = "NO";
    defparam add_7635_13.INJECT1_1 = "NO";
    CCU2C add_7635_11 (.A0(n3578), .B0(n30923), .C0(n64_adj_444), .D0(n1805), 
          .A1(n3577), .B1(n30923), .C1(n64_adj_444), .D1(n2137), .CIN(n32600), 
          .COUT(n32601), .S0(n3710), .S1(n3709));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_11.INIT0 = 16'ha9aa;
    defparam add_7635_11.INIT1 = 16'ha9aa;
    defparam add_7635_11.INJECT1_0 = "NO";
    defparam add_7635_11.INJECT1_1 = "NO";
    CCU2C add_7635_9 (.A0(n3580), .B0(n30923), .C0(n64_adj_444), .D0(n1462), 
          .A1(n3579), .B1(n30923), .C1(n64_adj_444), .D1(n1635), .CIN(n32599), 
          .COUT(n32600), .S0(n3712), .S1(n3711));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_9.INIT0 = 16'ha9aa;
    defparam add_7635_9.INIT1 = 16'ha9aa;
    defparam add_7635_9.INJECT1_0 = "NO";
    defparam add_7635_9.INJECT1_1 = "NO";
    CCU2C add_7635_7 (.A0(n3582), .B0(n30923), .C0(n64_adj_444), .D0(n2142), 
          .A1(n3581), .B1(n30923), .C1(n64_adj_444), .D1(n2141), .CIN(n32598), 
          .COUT(n32599), .S0(n3714), .S1(n3713));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_7.INIT0 = 16'ha9aa;
    defparam add_7635_7.INIT1 = 16'ha9aa;
    defparam add_7635_7.INJECT1_0 = "NO";
    defparam add_7635_7.INJECT1_1 = "NO";
    CCU2C add_7635_5 (.A0(n3584), .B0(n30923), .C0(n64_adj_444), .D0(n42824), 
          .A1(n3583), .B1(n30923), .C1(n64_adj_444), .D1(n42822), .CIN(n32597), 
          .COUT(n32598), .S0(n3716), .S1(n3715));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_5.INIT0 = 16'ha9aa;
    defparam add_7635_5.INIT1 = 16'ha9aa;
    defparam add_7635_5.INJECT1_0 = "NO";
    defparam add_7635_5.INJECT1_1 = "NO";
    CCU2C add_7635_3 (.A0(n883), .B0(n30923), .C0(n64_adj_444), .D0(n42827), 
          .A1(n3585), .B1(n30923), .C1(n64_adj_444), .D1(n42823), .CIN(n32596), 
          .COUT(n32597), .S0(n3718), .S1(n3717));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_3.INIT0 = 16'ha9aa;
    defparam add_7635_3.INIT1 = 16'ha9aa;
    defparam add_7635_3.INJECT1_0 = "NO";
    defparam add_7635_3.INJECT1_1 = "NO";
    CCU2C add_7635_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_444), .B1(n30923), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32596));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7635_1.INIT0 = 16'h0000;
    defparam add_7635_1.INIT1 = 16'heee1;
    defparam add_7635_1.INJECT1_0 = "NO";
    defparam add_7635_1.INJECT1_1 = "NO";
    CCU2C add_7634_21 (.A0(n3432), .B0(n30920), .C0(n64_adj_421), .D0(n3340), 
          .A1(n3431), .B1(n30920), .C1(n64_adj_421), .D1(n3477), .CIN(n32591), 
          .S0(n3567), .S1(n3566));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_21.INIT0 = 16'ha9aa;
    defparam add_7634_21.INIT1 = 16'ha9aa;
    defparam add_7634_21.INJECT1_0 = "NO";
    defparam add_7634_21.INJECT1_1 = "NO";
    CCU2C add_7634_19 (.A0(n3434), .B0(n30920), .C0(n64_adj_421), .D0(n3057), 
          .A1(n3433), .B1(n30920), .C1(n64_adj_421), .D1(n3479), .CIN(n32590), 
          .COUT(n32591), .S0(n3569), .S1(n3568));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_19.INIT0 = 16'ha9aa;
    defparam add_7634_19.INIT1 = 16'ha9aa;
    defparam add_7634_19.INJECT1_0 = "NO";
    defparam add_7634_19.INJECT1_1 = "NO";
    CCU2C add_7634_17 (.A0(n3436), .B0(n30920), .C0(n64_adj_421), .D0(n2762), 
          .A1(n3435), .B1(n30920), .C1(n64_adj_421), .D1(n2911), .CIN(n32589), 
          .COUT(n32590), .S0(n3571), .S1(n3570));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_17.INIT0 = 16'ha9aa;
    defparam add_7634_17.INIT1 = 16'ha9aa;
    defparam add_7634_17.INJECT1_0 = "NO";
    defparam add_7634_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1103_3_lut_4_lut (.A(n111), .B(n110_adj_220), .C(n108), 
         .D(n109_adj_219), .Z(n42802)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1103_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX x_3___i7 (.D(n5519), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i7.GSR = "ENABLED";
    FD1P3IX x_3___i8 (.D(n5518), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i8.GSR = "ENABLED";
    FD1P3IX x_3___i9 (.D(n5517), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i9.GSR = "ENABLED";
    FD1P3IX x_3___i10 (.D(n5516), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i10.GSR = "ENABLED";
    FD1P3IX x_3___i11 (.D(n5515), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i11.GSR = "ENABLED";
    FD1P3IX x_3___i12 (.D(n5514), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i12.GSR = "ENABLED";
    FD1P3IX x_3___i13 (.D(n5513), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i13.GSR = "ENABLED";
    FD1P3IX x_3___i14 (.D(n5512), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i14.GSR = "ENABLED";
    FD1P3IX x_3___i15 (.D(n5511), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i15.GSR = "ENABLED";
    FD1P3IX x_3___i16 (.D(n5510), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i16.GSR = "ENABLED";
    FD1P3IX x_3___i17 (.D(n5509), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i17.GSR = "ENABLED";
    FD1P3IX x_3___i18 (.D(n5508), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i18.GSR = "ENABLED";
    FD1P3IX x_3___i19 (.D(n5507), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i19.GSR = "ENABLED";
    FD1P3IX x_3___i20 (.D(n5506), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i20.GSR = "ENABLED";
    FD1P3IX x_3___i21 (.D(n5505), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i21.GSR = "ENABLED";
    FD1P3IX x_3___i22 (.D(n5504), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i22.GSR = "ENABLED";
    FD1P3IX x_3___i23 (.D(n5503), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i23.GSR = "ENABLED";
    FD1P3IX x_3___i24 (.D(n5502), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i24.GSR = "ENABLED";
    FD1P3IX x_3___i25 (.D(n5501), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i25.GSR = "ENABLED";
    FD1P3IX x_3___i26 (.D(n5500), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i26.GSR = "ENABLED";
    FD1P3IX x_3___i27 (.D(n5499), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i27.GSR = "ENABLED";
    FD1P3IX x_3___i28 (.D(n5498), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i28.GSR = "ENABLED";
    FD1P3IX x_3___i29 (.D(n5497), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i29.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_1112 (.A(n112_adj_221), .B(n115_adj_223), .Z(n42811)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1112.init = 16'heeee;
    OB x_out_pad_20 (.I(x_out_c_20), .O(x_out[20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_21 (.I(x_out_c_21), .O(x_out[21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_22 (.I(x_out_c_22), .O(x_out[22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_23 (.I(x_out_c_23), .O(x_out[23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_24 (.I(x_out_c_24), .O(x_out[24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_25 (.I(x_out_c_25), .O(x_out[25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_26 (.I(x_out_c_26), .O(x_out[26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_27 (.I(x_out_c_27), .O(x_out[27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7634_15 (.A0(n3438), .B0(n30920), .C0(n64_adj_421), .D0(n2455), 
          .A1(n3437), .B1(n30920), .C1(n64_adj_421), .D1(n3060), .CIN(n32588), 
          .COUT(n32589), .S0(n3573), .S1(n3572));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_15.INIT0 = 16'ha9aa;
    defparam add_7634_15.INIT1 = 16'ha9aa;
    defparam add_7634_15.INJECT1_0 = "NO";
    defparam add_7634_15.INJECT1_1 = "NO";
    CCU2C add_7634_13 (.A0(n3440), .B0(n30920), .C0(n64_adj_421), .D0(n2298), 
          .A1(n3439), .B1(n30920), .C1(n64_adj_421), .D1(n2456), .CIN(n32587), 
          .COUT(n32588), .S0(n3575), .S1(n3574));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_13.INIT0 = 16'ha9aa;
    defparam add_7634_13.INIT1 = 16'ha9aa;
    defparam add_7634_13.INJECT1_0 = "NO";
    defparam add_7634_13.INJECT1_1 = "NO";
    CCU2C add_7634_11 (.A0(n3442), .B0(n30920), .C0(n64_adj_421), .D0(n1805), 
          .A1(n3441), .B1(n30920), .C1(n64_adj_421), .D1(n2137), .CIN(n32586), 
          .COUT(n32587), .S0(n3577), .S1(n3576));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_11.INIT0 = 16'ha9aa;
    defparam add_7634_11.INIT1 = 16'ha9aa;
    defparam add_7634_11.INJECT1_0 = "NO";
    defparam add_7634_11.INJECT1_1 = "NO";
    CCU2C add_7634_9 (.A0(n3444), .B0(n30920), .C0(n64_adj_421), .D0(n1462), 
          .A1(n3443), .B1(n30920), .C1(n64_adj_421), .D1(n1635), .CIN(n32585), 
          .COUT(n32586), .S0(n3579), .S1(n3578));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_9.INIT0 = 16'ha9aa;
    defparam add_7634_9.INIT1 = 16'ha9aa;
    defparam add_7634_9.INJECT1_0 = "NO";
    defparam add_7634_9.INJECT1_1 = "NO";
    CCU2C add_7634_7 (.A0(n3446), .B0(n30920), .C0(n64_adj_421), .D0(n2142), 
          .A1(n3445), .B1(n30920), .C1(n64_adj_421), .D1(n2141), .CIN(n32584), 
          .COUT(n32585), .S0(n3581), .S1(n3580));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_7.INIT0 = 16'ha9aa;
    defparam add_7634_7.INIT1 = 16'ha9aa;
    defparam add_7634_7.INJECT1_0 = "NO";
    defparam add_7634_7.INJECT1_1 = "NO";
    CCU2C add_7634_5 (.A0(n3448), .B0(n30920), .C0(n64_adj_421), .D0(n42824), 
          .A1(n3447), .B1(n30920), .C1(n64_adj_421), .D1(n42822), .CIN(n32583), 
          .COUT(n32584), .S0(n3583), .S1(n3582));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_5.INIT0 = 16'ha9aa;
    defparam add_7634_5.INIT1 = 16'ha9aa;
    defparam add_7634_5.INJECT1_0 = "NO";
    defparam add_7634_5.INJECT1_1 = "NO";
    CCU2C add_7634_3 (.A0(n882), .B0(n30920), .C0(n64_adj_421), .D0(n42827), 
          .A1(n3449), .B1(n30920), .C1(n64_adj_421), .D1(n42823), .CIN(n32582), 
          .COUT(n32583), .S0(n3585), .S1(n3584));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_3.INIT0 = 16'ha9aa;
    defparam add_7634_3.INIT1 = 16'ha9aa;
    defparam add_7634_3.INJECT1_0 = "NO";
    defparam add_7634_3.INJECT1_1 = "NO";
    CCU2C add_7634_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_421), .B1(n30920), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32582));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7634_1.INIT0 = 16'h0000;
    defparam add_7634_1.INIT1 = 16'heee1;
    defparam add_7634_1.INJECT1_0 = "NO";
    defparam add_7634_1.INJECT1_1 = "NO";
    CCU2C add_7633_21 (.A0(n3293), .B0(n30917), .C0(n64_adj_399), .D0(n3340), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32578), 
          .S0(n3431));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_21.INIT0 = 16'ha9aa;
    defparam add_7633_21.INIT1 = 16'h0000;
    defparam add_7633_21.INJECT1_0 = "NO";
    defparam add_7633_21.INJECT1_1 = "NO";
    CCU2C add_7633_19 (.A0(n3295), .B0(n30917), .C0(n64_adj_399), .D0(n3057), 
          .A1(n3294), .B1(n30917), .C1(n64_adj_399), .D1(n3479), .CIN(n32577), 
          .COUT(n32578), .S0(n3433), .S1(n3432));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_19.INIT0 = 16'ha9aa;
    defparam add_7633_19.INIT1 = 16'ha9aa;
    defparam add_7633_19.INJECT1_0 = "NO";
    defparam add_7633_19.INJECT1_1 = "NO";
    CCU2C add_7633_17 (.A0(n3297), .B0(n30917), .C0(n64_adj_399), .D0(n2762), 
          .A1(n3296), .B1(n30917), .C1(n64_adj_399), .D1(n2911), .CIN(n32576), 
          .COUT(n32577), .S0(n3435), .S1(n3434));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_17.INIT0 = 16'ha9aa;
    defparam add_7633_17.INIT1 = 16'ha9aa;
    defparam add_7633_17.INJECT1_0 = "NO";
    defparam add_7633_17.INJECT1_1 = "NO";
    CCU2C add_7633_15 (.A0(n3299), .B0(n30917), .C0(n64_adj_399), .D0(n2455), 
          .A1(n3298), .B1(n30917), .C1(n64_adj_399), .D1(n3060), .CIN(n32575), 
          .COUT(n32576), .S0(n3437), .S1(n3436));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_15.INIT0 = 16'ha9aa;
    defparam add_7633_15.INIT1 = 16'ha9aa;
    defparam add_7633_15.INJECT1_0 = "NO";
    defparam add_7633_15.INJECT1_1 = "NO";
    CCU2C add_7633_13 (.A0(n3301), .B0(n30917), .C0(n64_adj_399), .D0(n2298), 
          .A1(n3300), .B1(n30917), .C1(n64_adj_399), .D1(n2456), .CIN(n32574), 
          .COUT(n32575), .S0(n3439), .S1(n3438));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_13.INIT0 = 16'ha9aa;
    defparam add_7633_13.INIT1 = 16'ha9aa;
    defparam add_7633_13.INJECT1_0 = "NO";
    defparam add_7633_13.INJECT1_1 = "NO";
    CCU2C add_7633_11 (.A0(n3303), .B0(n30917), .C0(n64_adj_399), .D0(n1805), 
          .A1(n3302), .B1(n30917), .C1(n64_adj_399), .D1(n2137), .CIN(n32573), 
          .COUT(n32574), .S0(n3441), .S1(n3440));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_11.INIT0 = 16'ha9aa;
    defparam add_7633_11.INIT1 = 16'ha9aa;
    defparam add_7633_11.INJECT1_0 = "NO";
    defparam add_7633_11.INJECT1_1 = "NO";
    CCU2C add_7633_9 (.A0(n3305), .B0(n30917), .C0(n64_adj_399), .D0(n1462), 
          .A1(n3304), .B1(n30917), .C1(n64_adj_399), .D1(n1635), .CIN(n32572), 
          .COUT(n32573), .S0(n3443), .S1(n3442));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_9.INIT0 = 16'ha9aa;
    defparam add_7633_9.INIT1 = 16'ha9aa;
    defparam add_7633_9.INJECT1_0 = "NO";
    defparam add_7633_9.INJECT1_1 = "NO";
    CCU2C add_7633_7 (.A0(n3307), .B0(n30917), .C0(n64_adj_399), .D0(n2142), 
          .A1(n3306), .B1(n30917), .C1(n64_adj_399), .D1(n2141), .CIN(n32571), 
          .COUT(n32572), .S0(n3445), .S1(n3444));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_7.INIT0 = 16'ha9aa;
    defparam add_7633_7.INIT1 = 16'ha9aa;
    defparam add_7633_7.INJECT1_0 = "NO";
    defparam add_7633_7.INJECT1_1 = "NO";
    CCU2C add_7633_5 (.A0(n3309), .B0(n30917), .C0(n64_adj_399), .D0(n42824), 
          .A1(n3308), .B1(n30917), .C1(n64_adj_399), .D1(n42822), .CIN(n32570), 
          .COUT(n32571), .S0(n3447), .S1(n3446));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_5.INIT0 = 16'ha9aa;
    defparam add_7633_5.INIT1 = 16'ha9aa;
    defparam add_7633_5.INJECT1_0 = "NO";
    defparam add_7633_5.INJECT1_1 = "NO";
    CCU2C add_7633_3 (.A0(n881), .B0(n30917), .C0(n64_adj_399), .D0(n42827), 
          .A1(n3310), .B1(n30917), .C1(n64_adj_399), .D1(n42823), .CIN(n32569), 
          .COUT(n32570), .S0(n3449), .S1(n3448));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_3.INIT0 = 16'ha9aa;
    defparam add_7633_3.INIT1 = 16'ha9aa;
    defparam add_7633_3.INJECT1_0 = "NO";
    defparam add_7633_3.INJECT1_1 = "NO";
    CCU2C add_7633_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_399), .B1(n30917), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32569));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7633_1.INIT0 = 16'h0000;
    defparam add_7633_1.INIT1 = 16'heee1;
    defparam add_7633_1.INJECT1_0 = "NO";
    defparam add_7633_1.INJECT1_1 = "NO";
    CCU2C add_7632_19 (.A0(n3153), .B0(n30914), .C0(n64_adj_378), .D0(n3057), 
          .A1(n3152), .B1(n30914), .C1(n64_adj_378), .D1(n3479), .CIN(n32564), 
          .S0(n3294), .S1(n3293));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_19.INIT0 = 16'ha9aa;
    defparam add_7632_19.INIT1 = 16'ha9aa;
    defparam add_7632_19.INJECT1_0 = "NO";
    defparam add_7632_19.INJECT1_1 = "NO";
    CCU2C add_7632_17 (.A0(n3155), .B0(n30914), .C0(n64_adj_378), .D0(n2762), 
          .A1(n3154), .B1(n30914), .C1(n64_adj_378), .D1(n2911), .CIN(n32563), 
          .COUT(n32564), .S0(n3296), .S1(n3295));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_17.INIT0 = 16'ha9aa;
    defparam add_7632_17.INIT1 = 16'ha9aa;
    defparam add_7632_17.INJECT1_0 = "NO";
    defparam add_7632_17.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_53 (.A(n112_adj_221), .B(n115_adj_223), .C(n113_adj_222), 
         .D(n111), .Z(n37274)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_53.init = 16'hfffe;
    FD1P3IX x_3___i30 (.D(n5496), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i30.GSR = "ENABLED";
    FD1P3IX x_3___i31 (.D(n5495), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i31.GSR = "ENABLED";
    FD1P3IX x_3___i32 (.D(n5494), .SP(clk_c_enable_829), .CD(n31084), 
            .CK(clk_c), .Q(\x[3] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i32.GSR = "ENABLED";
    FD1P3IX x_3___i33 (.D(n5525), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i33.GSR = "ENABLED";
    FD1P3IX x_3___i34 (.D(n5524), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i34.GSR = "ENABLED";
    FD1P3IX x_3___i35 (.D(n5523), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i35.GSR = "ENABLED";
    FD1P3IX x_3___i36 (.D(n5522), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i36.GSR = "ENABLED";
    FD1P3IX x_3___i37 (.D(n5521), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i37.GSR = "ENABLED";
    FD1P3IX x_3___i38 (.D(n5520), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i38.GSR = "ENABLED";
    FD1P3IX x_3___i39 (.D(n5519), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i39.GSR = "ENABLED";
    FD1P3IX x_3___i40 (.D(n5518), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i40.GSR = "ENABLED";
    FD1P3IX x_3___i41 (.D(n5517), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i41.GSR = "ENABLED";
    FD1P3IX x_3___i42 (.D(n5516), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i42.GSR = "ENABLED";
    FD1P3IX x_3___i43 (.D(n5515), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i43.GSR = "ENABLED";
    FD1P3IX x_3___i44 (.D(n5514), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i44.GSR = "ENABLED";
    FD1P3IX x_3___i45 (.D(n5513), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i45.GSR = "ENABLED";
    FD1P3IX x_3___i46 (.D(n5512), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i46.GSR = "ENABLED";
    FD1P3IX x_3___i47 (.D(n5511), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i47.GSR = "ENABLED";
    FD1P3IX x_3___i48 (.D(n5510), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i48.GSR = "ENABLED";
    FD1P3IX x_3___i49 (.D(n5509), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i49.GSR = "ENABLED";
    FD1P3IX x_3___i50 (.D(n5508), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i50.GSR = "ENABLED";
    FD1P3IX x_3___i51 (.D(n5507), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i51.GSR = "ENABLED";
    FD1P3IX x_3___i52 (.D(n5506), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i52.GSR = "ENABLED";
    FD1P3IX x_3___i53 (.D(n5505), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i53.GSR = "ENABLED";
    FD1P3IX x_3___i54 (.D(n5504), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i54.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_54 (.A(n112_adj_221), .B(n115_adj_223), .C(n116_adj_224), 
         .D(n114), .Z(n37240)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_54.init = 16'hfffe;
    OB x_out_pad_28 (.I(x_out_c_28), .O(x_out[28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_29 (.I(x_out_c_29), .O(x_out[29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_30 (.I(x_out_c_30), .O(x_out[30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_31 (.I(x_out_c_31), .O(x_out[31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_32 (.I(x_out_c_32), .O(x_out[32]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_33 (.I(x_out_c_33), .O(x_out[33]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_34 (.I(x_out_c_34), .O(x_out[34]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7632_15 (.A0(n3157), .B0(n30914), .C0(n64_adj_378), .D0(n2455), 
          .A1(n3156), .B1(n30914), .C1(n64_adj_378), .D1(n3060), .CIN(n32562), 
          .COUT(n32563), .S0(n3298), .S1(n3297));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_15.INIT0 = 16'ha9aa;
    defparam add_7632_15.INIT1 = 16'ha9aa;
    defparam add_7632_15.INJECT1_0 = "NO";
    defparam add_7632_15.INJECT1_1 = "NO";
    CCU2C add_7632_13 (.A0(n3159), .B0(n30914), .C0(n64_adj_378), .D0(n2298), 
          .A1(n3158), .B1(n30914), .C1(n64_adj_378), .D1(n2456), .CIN(n32561), 
          .COUT(n32562), .S0(n3300), .S1(n3299));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_13.INIT0 = 16'ha9aa;
    defparam add_7632_13.INIT1 = 16'ha9aa;
    defparam add_7632_13.INJECT1_0 = "NO";
    defparam add_7632_13.INJECT1_1 = "NO";
    CCU2C add_7632_11 (.A0(n3161), .B0(n30914), .C0(n64_adj_378), .D0(n1805), 
          .A1(n3160), .B1(n30914), .C1(n64_adj_378), .D1(n2137), .CIN(n32560), 
          .COUT(n32561), .S0(n3302), .S1(n3301));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_11.INIT0 = 16'ha9aa;
    defparam add_7632_11.INIT1 = 16'ha9aa;
    defparam add_7632_11.INJECT1_0 = "NO";
    defparam add_7632_11.INJECT1_1 = "NO";
    CCU2C add_7632_9 (.A0(n3163), .B0(n30914), .C0(n64_adj_378), .D0(n1462), 
          .A1(n3162), .B1(n30914), .C1(n64_adj_378), .D1(n1635), .CIN(n32559), 
          .COUT(n32560), .S0(n3304), .S1(n3303));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_9.INIT0 = 16'ha9aa;
    defparam add_7632_9.INIT1 = 16'ha9aa;
    defparam add_7632_9.INJECT1_0 = "NO";
    defparam add_7632_9.INJECT1_1 = "NO";
    CCU2C add_7632_7 (.A0(n3165), .B0(n30914), .C0(n64_adj_378), .D0(n2142), 
          .A1(n3164), .B1(n30914), .C1(n64_adj_378), .D1(n2141), .CIN(n32558), 
          .COUT(n32559), .S0(n3306), .S1(n3305));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_7.INIT0 = 16'ha9aa;
    defparam add_7632_7.INIT1 = 16'ha9aa;
    defparam add_7632_7.INJECT1_0 = "NO";
    defparam add_7632_7.INJECT1_1 = "NO";
    CCU2C add_7632_5 (.A0(n3167), .B0(n30914), .C0(n64_adj_378), .D0(n42824), 
          .A1(n3166), .B1(n30914), .C1(n64_adj_378), .D1(n42822), .CIN(n32557), 
          .COUT(n32558), .S0(n3308), .S1(n3307));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_5.INIT0 = 16'ha9aa;
    defparam add_7632_5.INIT1 = 16'ha9aa;
    defparam add_7632_5.INJECT1_0 = "NO";
    defparam add_7632_5.INJECT1_1 = "NO";
    CCU2C add_7632_3 (.A0(n880), .B0(n30914), .C0(n64_adj_378), .D0(n42827), 
          .A1(n3168), .B1(n30914), .C1(n64_adj_378), .D1(n42823), .CIN(n32556), 
          .COUT(n32557), .S0(n3310), .S1(n3309));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_3.INIT0 = 16'ha9aa;
    defparam add_7632_3.INIT1 = 16'ha9aa;
    defparam add_7632_3.INJECT1_0 = "NO";
    defparam add_7632_3.INJECT1_1 = "NO";
    CCU2C add_7632_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_378), .B1(n30914), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32556));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7632_1.INIT0 = 16'h0000;
    defparam add_7632_1.INIT1 = 16'heee1;
    defparam add_7632_1.INJECT1_0 = "NO";
    defparam add_7632_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1106_3_lut_4_lut (.A(n112_adj_221), .B(n115_adj_223), 
         .C(n113_adj_222), .D(n110_adj_220), .Z(n42805)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1106_3_lut_4_lut.init = 16'hfffe;
    CCU2C add_7631_19 (.A0(n3008), .B0(n30911), .C0(n64_adj_360), .D0(n3057), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32552), 
          .S0(n3152));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_19.INIT0 = 16'ha9aa;
    defparam add_7631_19.INIT1 = 16'h0000;
    defparam add_7631_19.INJECT1_0 = "NO";
    defparam add_7631_19.INJECT1_1 = "NO";
    CCU2C add_7631_17 (.A0(n3010), .B0(n30911), .C0(n64_adj_360), .D0(n2762), 
          .A1(n3009), .B1(n30911), .C1(n64_adj_360), .D1(n2911), .CIN(n32551), 
          .COUT(n32552), .S0(n3154), .S1(n3153));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_17.INIT0 = 16'ha9aa;
    defparam add_7631_17.INIT1 = 16'ha9aa;
    defparam add_7631_17.INJECT1_0 = "NO";
    defparam add_7631_17.INJECT1_1 = "NO";
    CCU2C add_7631_15 (.A0(n3012), .B0(n30911), .C0(n64_adj_360), .D0(n2455), 
          .A1(n3011), .B1(n30911), .C1(n64_adj_360), .D1(n3060), .CIN(n32550), 
          .COUT(n32551), .S0(n3156), .S1(n3155));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_15.INIT0 = 16'ha9aa;
    defparam add_7631_15.INIT1 = 16'ha9aa;
    defparam add_7631_15.INJECT1_0 = "NO";
    defparam add_7631_15.INJECT1_1 = "NO";
    CCU2C add_7631_13 (.A0(n3014), .B0(n30911), .C0(n64_adj_360), .D0(n2298), 
          .A1(n3013), .B1(n30911), .C1(n64_adj_360), .D1(n2456), .CIN(n32549), 
          .COUT(n32550), .S0(n3158), .S1(n3157));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_13.INIT0 = 16'ha9aa;
    defparam add_7631_13.INIT1 = 16'ha9aa;
    defparam add_7631_13.INJECT1_0 = "NO";
    defparam add_7631_13.INJECT1_1 = "NO";
    CCU2C add_7631_11 (.A0(n3016), .B0(n30911), .C0(n64_adj_360), .D0(n1805), 
          .A1(n3015), .B1(n30911), .C1(n64_adj_360), .D1(n2137), .CIN(n32548), 
          .COUT(n32549), .S0(n3160), .S1(n3159));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_11.INIT0 = 16'ha9aa;
    defparam add_7631_11.INIT1 = 16'ha9aa;
    defparam add_7631_11.INJECT1_0 = "NO";
    defparam add_7631_11.INJECT1_1 = "NO";
    CCU2C add_7631_9 (.A0(n3018), .B0(n30911), .C0(n64_adj_360), .D0(n1462), 
          .A1(n3017), .B1(n30911), .C1(n64_adj_360), .D1(n1635), .CIN(n32547), 
          .COUT(n32548), .S0(n3162), .S1(n3161));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_9.INIT0 = 16'ha9aa;
    defparam add_7631_9.INIT1 = 16'ha9aa;
    defparam add_7631_9.INJECT1_0 = "NO";
    defparam add_7631_9.INJECT1_1 = "NO";
    CCU2C add_7631_7 (.A0(n3020), .B0(n30911), .C0(n64_adj_360), .D0(n2142), 
          .A1(n3019), .B1(n30911), .C1(n64_adj_360), .D1(n2141), .CIN(n32546), 
          .COUT(n32547), .S0(n3164), .S1(n3163));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_7.INIT0 = 16'ha9aa;
    defparam add_7631_7.INIT1 = 16'ha9aa;
    defparam add_7631_7.INJECT1_0 = "NO";
    defparam add_7631_7.INJECT1_1 = "NO";
    CCU2C add_7631_5 (.A0(n3022), .B0(n30911), .C0(n64_adj_360), .D0(n42824), 
          .A1(n3021), .B1(n30911), .C1(n64_adj_360), .D1(n42822), .CIN(n32545), 
          .COUT(n32546), .S0(n3166), .S1(n3165));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_5.INIT0 = 16'ha9aa;
    defparam add_7631_5.INIT1 = 16'ha9aa;
    defparam add_7631_5.INJECT1_0 = "NO";
    defparam add_7631_5.INJECT1_1 = "NO";
    CCU2C add_7631_3 (.A0(n879), .B0(n30911), .C0(n64_adj_360), .D0(n42827), 
          .A1(n3023), .B1(n30911), .C1(n64_adj_360), .D1(n42823), .CIN(n32544), 
          .COUT(n32545), .S0(n3168), .S1(n3167));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_3.INIT0 = 16'ha9aa;
    defparam add_7631_3.INIT1 = 16'ha9aa;
    defparam add_7631_3.INJECT1_0 = "NO";
    defparam add_7631_3.INJECT1_1 = "NO";
    CCU2C add_7631_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_360), .B1(n30911), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32544));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7631_1.INIT0 = 16'h0000;
    defparam add_7631_1.INIT1 = 16'heee1;
    defparam add_7631_1.INJECT1_0 = "NO";
    defparam add_7631_1.INJECT1_1 = "NO";
    CCU2C add_7630_17 (.A0(n2862), .B0(n30908), .C0(n64_adj_343), .D0(n2762), 
          .A1(n2861), .B1(n30908), .C1(n64_adj_343), .D1(n2911), .CIN(n32539), 
          .S0(n3009), .S1(n3008));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_17.INIT0 = 16'ha9aa;
    defparam add_7630_17.INIT1 = 16'ha9aa;
    defparam add_7630_17.INJECT1_0 = "NO";
    defparam add_7630_17.INJECT1_1 = "NO";
    CCU2C add_7630_15 (.A0(n2864), .B0(n30908), .C0(n64_adj_343), .D0(n2455), 
          .A1(n2863), .B1(n30908), .C1(n64_adj_343), .D1(n3060), .CIN(n32538), 
          .COUT(n32539), .S0(n3011), .S1(n3010));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_15.INIT0 = 16'ha9aa;
    defparam add_7630_15.INIT1 = 16'ha9aa;
    defparam add_7630_15.INJECT1_0 = "NO";
    defparam add_7630_15.INJECT1_1 = "NO";
    CCU2C add_7630_13 (.A0(n2866), .B0(n30908), .C0(n64_adj_343), .D0(n2298), 
          .A1(n2865), .B1(n30908), .C1(n64_adj_343), .D1(n2456), .CIN(n32537), 
          .COUT(n32538), .S0(n3013), .S1(n3012));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_13.INIT0 = 16'ha9aa;
    defparam add_7630_13.INIT1 = 16'ha9aa;
    defparam add_7630_13.INJECT1_0 = "NO";
    defparam add_7630_13.INJECT1_1 = "NO";
    CCU2C add_7630_11 (.A0(n2868), .B0(n30908), .C0(n64_adj_343), .D0(n1805), 
          .A1(n2867), .B1(n30908), .C1(n64_adj_343), .D1(n2137), .CIN(n32536), 
          .COUT(n32537), .S0(n3015), .S1(n3014));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_11.INIT0 = 16'ha9aa;
    defparam add_7630_11.INIT1 = 16'ha9aa;
    defparam add_7630_11.INJECT1_0 = "NO";
    defparam add_7630_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1113 (.A(n112_adj_221), .B(n114), .Z(n42812)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1113.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_55 (.A(n112_adj_221), .B(n114), .C(n113_adj_222), 
         .D(n110_adj_220), .Z(n37082)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_55.init = 16'hfffe;
    FD1P3IX x_3___i55 (.D(n5503), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i55.GSR = "ENABLED";
    FD1P3IX x_3___i56 (.D(n5502), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i56.GSR = "ENABLED";
    FD1P3IX x_3___i57 (.D(n5501), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i57.GSR = "ENABLED";
    FD1P3IX x_3___i58 (.D(n5500), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i58.GSR = "ENABLED";
    FD1P3IX x_3___i59 (.D(n5499), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i59.GSR = "ENABLED";
    FD1P3IX x_3___i60 (.D(n5498), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i60.GSR = "ENABLED";
    FD1P3IX x_3___i61 (.D(n5497), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i61.GSR = "ENABLED";
    FD1P3IX x_3___i62 (.D(n5496), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i62.GSR = "ENABLED";
    FD1P3IX x_3___i63 (.D(n5495), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i63.GSR = "ENABLED";
    FD1P3IX x_3___i64 (.D(n5494), .SP(clk_c_enable_780), .CD(n31054), 
            .CK(clk_c), .Q(\x[2] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i64.GSR = "ENABLED";
    FD1P3IX x_3___i65 (.D(n5525), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i65.GSR = "ENABLED";
    FD1P3IX x_3___i66 (.D(n5524), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i66.GSR = "ENABLED";
    FD1P3IX x_3___i67 (.D(n5523), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i67.GSR = "ENABLED";
    FD1P3IX x_3___i68 (.D(n5522), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i68.GSR = "ENABLED";
    FD1P3IX x_3___i69 (.D(n5521), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i69.GSR = "ENABLED";
    FD1P3IX x_3___i70 (.D(n5520), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i70.GSR = "ENABLED";
    FD1P3IX x_3___i71 (.D(n5519), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i71.GSR = "ENABLED";
    FD1P3IX x_3___i72 (.D(n5518), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i72.GSR = "ENABLED";
    FD1P3IX x_3___i73 (.D(n5517), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i73.GSR = "ENABLED";
    FD1P3IX x_3___i74 (.D(n5516), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i74.GSR = "ENABLED";
    FD1P3IX x_3___i75 (.D(n5515), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [10]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i75.GSR = "ENABLED";
    FD1P3IX x_3___i76 (.D(n5514), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [11]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i76.GSR = "ENABLED";
    FD1P3IX x_3___i77 (.D(n5513), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [12]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i77.GSR = "ENABLED";
    FD1P3IX x_3___i78 (.D(n5512), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [13]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i78.GSR = "ENABLED";
    OB x_out_pad_35 (.I(x_out_c_35), .O(x_out[35]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_36 (.I(x_out_c_36), .O(x_out[36]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_37 (.I(x_out_c_37), .O(x_out[37]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_38 (.I(x_out_c_38), .O(x_out[38]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_39 (.I(x_out_c_39), .O(x_out[39]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_40 (.I(x_out_c_40), .O(x_out[40]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7630_9 (.A0(n2870), .B0(n30908), .C0(n64_adj_343), .D0(n1462), 
          .A1(n2869), .B1(n30908), .C1(n64_adj_343), .D1(n1635), .CIN(n32535), 
          .COUT(n32536), .S0(n3017), .S1(n3016));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_9.INIT0 = 16'ha9aa;
    defparam add_7630_9.INIT1 = 16'ha9aa;
    defparam add_7630_9.INJECT1_0 = "NO";
    defparam add_7630_9.INJECT1_1 = "NO";
    CCU2C add_7630_7 (.A0(n2872), .B0(n30908), .C0(n64_adj_343), .D0(n2142), 
          .A1(n2871), .B1(n30908), .C1(n64_adj_343), .D1(n2141), .CIN(n32534), 
          .COUT(n32535), .S0(n3019), .S1(n3018));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_7.INIT0 = 16'ha9aa;
    defparam add_7630_7.INIT1 = 16'ha9aa;
    defparam add_7630_7.INJECT1_0 = "NO";
    defparam add_7630_7.INJECT1_1 = "NO";
    CCU2C add_7630_5 (.A0(n2874), .B0(n30908), .C0(n64_adj_343), .D0(n42824), 
          .A1(n2873), .B1(n30908), .C1(n64_adj_343), .D1(n42822), .CIN(n32533), 
          .COUT(n32534), .S0(n3021), .S1(n3020));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_5.INIT0 = 16'ha9aa;
    defparam add_7630_5.INIT1 = 16'ha9aa;
    defparam add_7630_5.INJECT1_0 = "NO";
    defparam add_7630_5.INJECT1_1 = "NO";
    CCU2C add_7630_3 (.A0(n878), .B0(n30908), .C0(n64_adj_343), .D0(n42827), 
          .A1(n2875), .B1(n30908), .C1(n64_adj_343), .D1(n42823), .CIN(n32532), 
          .COUT(n32533), .S0(n3023), .S1(n3022));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_3.INIT0 = 16'ha9aa;
    defparam add_7630_3.INIT1 = 16'ha9aa;
    defparam add_7630_3.INJECT1_0 = "NO";
    defparam add_7630_3.INJECT1_1 = "NO";
    CCU2C add_7630_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_343), .B1(n30908), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32532));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7630_1.INIT0 = 16'h0000;
    defparam add_7630_1.INIT1 = 16'heee1;
    defparam add_7630_1.INJECT1_0 = "NO";
    defparam add_7630_1.INJECT1_1 = "NO";
    CCU2C add_7629_17 (.A0(n2711), .B0(n30905), .C0(n64_adj_328), .D0(n2762), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32528), 
          .S0(n2861));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_17.INIT0 = 16'ha9aa;
    defparam add_7629_17.INIT1 = 16'h0000;
    defparam add_7629_17.INJECT1_0 = "NO";
    defparam add_7629_17.INJECT1_1 = "NO";
    CCU2C add_7629_15 (.A0(n2713), .B0(n30905), .C0(n64_adj_328), .D0(n2455), 
          .A1(n2712), .B1(n30905), .C1(n64_adj_328), .D1(n3060), .CIN(n32527), 
          .COUT(n32528), .S0(n2863), .S1(n2862));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_15.INIT0 = 16'ha9aa;
    defparam add_7629_15.INIT1 = 16'ha9aa;
    defparam add_7629_15.INJECT1_0 = "NO";
    defparam add_7629_15.INJECT1_1 = "NO";
    CCU2C add_7629_13 (.A0(n2715), .B0(n30905), .C0(n64_adj_328), .D0(n2298), 
          .A1(n2714), .B1(n30905), .C1(n64_adj_328), .D1(n2456), .CIN(n32526), 
          .COUT(n32527), .S0(n2865), .S1(n2864));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_13.INIT0 = 16'ha9aa;
    defparam add_7629_13.INIT1 = 16'ha9aa;
    defparam add_7629_13.INJECT1_0 = "NO";
    defparam add_7629_13.INJECT1_1 = "NO";
    CCU2C add_7629_11 (.A0(n2717), .B0(n30905), .C0(n64_adj_328), .D0(n1805), 
          .A1(n2716), .B1(n30905), .C1(n64_adj_328), .D1(n2137), .CIN(n32525), 
          .COUT(n32526), .S0(n2867), .S1(n2866));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_11.INIT0 = 16'ha9aa;
    defparam add_7629_11.INIT1 = 16'ha9aa;
    defparam add_7629_11.INJECT1_0 = "NO";
    defparam add_7629_11.INJECT1_1 = "NO";
    CCU2C add_7629_9 (.A0(n2719), .B0(n30905), .C0(n64_adj_328), .D0(n1462), 
          .A1(n2718), .B1(n30905), .C1(n64_adj_328), .D1(n1635), .CIN(n32524), 
          .COUT(n32525), .S0(n2869), .S1(n2868));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_9.INIT0 = 16'ha9aa;
    defparam add_7629_9.INIT1 = 16'ha9aa;
    defparam add_7629_9.INJECT1_0 = "NO";
    defparam add_7629_9.INJECT1_1 = "NO";
    CCU2C add_7629_7 (.A0(n2721), .B0(n30905), .C0(n64_adj_328), .D0(n2142), 
          .A1(n2720), .B1(n30905), .C1(n64_adj_328), .D1(n2141), .CIN(n32523), 
          .COUT(n32524), .S0(n2871), .S1(n2870));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_7.INIT0 = 16'ha9aa;
    defparam add_7629_7.INIT1 = 16'ha9aa;
    defparam add_7629_7.INJECT1_0 = "NO";
    defparam add_7629_7.INJECT1_1 = "NO";
    CCU2C add_7629_5 (.A0(n2723), .B0(n30905), .C0(n64_adj_328), .D0(n42824), 
          .A1(n2722), .B1(n30905), .C1(n64_adj_328), .D1(n42822), .CIN(n32522), 
          .COUT(n32523), .S0(n2873), .S1(n2872));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_5.INIT0 = 16'ha9aa;
    defparam add_7629_5.INIT1 = 16'ha9aa;
    defparam add_7629_5.INJECT1_0 = "NO";
    defparam add_7629_5.INJECT1_1 = "NO";
    CCU2C add_7629_3 (.A0(n877), .B0(n30905), .C0(n64_adj_328), .D0(n42827), 
          .A1(n2724), .B1(n30905), .C1(n64_adj_328), .D1(n42823), .CIN(n32521), 
          .COUT(n32522), .S0(n2875), .S1(n2874));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_3.INIT0 = 16'ha9aa;
    defparam add_7629_3.INIT1 = 16'ha9aa;
    defparam add_7629_3.INJECT1_0 = "NO";
    defparam add_7629_3.INJECT1_1 = "NO";
    CCU2C add_7629_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_328), .B1(n30905), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32521));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7629_1.INIT0 = 16'h0000;
    defparam add_7629_1.INIT1 = 16'heee1;
    defparam add_7629_1.INJECT1_0 = "NO";
    defparam add_7629_1.INJECT1_1 = "NO";
    CCU2C add_7628_15 (.A0(n2559), .B0(n30902), .C0(n64_adj_315), .D0(n2455), 
          .A1(n2558), .B1(n30902), .C1(n64_adj_315), .D1(n3060), .CIN(n32516), 
          .S0(n2712), .S1(n2711));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_15.INIT0 = 16'ha9aa;
    defparam add_7628_15.INIT1 = 16'ha9aa;
    defparam add_7628_15.INJECT1_0 = "NO";
    defparam add_7628_15.INJECT1_1 = "NO";
    CCU2C add_7628_13 (.A0(n2561), .B0(n30902), .C0(n64_adj_315), .D0(n2298), 
          .A1(n2560), .B1(n30902), .C1(n64_adj_315), .D1(n2456), .CIN(n32515), 
          .COUT(n32516), .S0(n2714), .S1(n2713));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_13.INIT0 = 16'ha9aa;
    defparam add_7628_13.INIT1 = 16'ha9aa;
    defparam add_7628_13.INJECT1_0 = "NO";
    defparam add_7628_13.INJECT1_1 = "NO";
    CCU2C add_7628_11 (.A0(n2563), .B0(n30902), .C0(n64_adj_315), .D0(n1805), 
          .A1(n2562), .B1(n30902), .C1(n64_adj_315), .D1(n2137), .CIN(n32514), 
          .COUT(n32515), .S0(n2716), .S1(n2715));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_11.INIT0 = 16'ha9aa;
    defparam add_7628_11.INIT1 = 16'ha9aa;
    defparam add_7628_11.INJECT1_0 = "NO";
    defparam add_7628_11.INJECT1_1 = "NO";
    CCU2C add_7628_9 (.A0(n2565), .B0(n30902), .C0(n64_adj_315), .D0(n1462), 
          .A1(n2564), .B1(n30902), .C1(n64_adj_315), .D1(n1635), .CIN(n32513), 
          .COUT(n32514), .S0(n2718), .S1(n2717));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_9.INIT0 = 16'ha9aa;
    defparam add_7628_9.INIT1 = 16'ha9aa;
    defparam add_7628_9.INJECT1_0 = "NO";
    defparam add_7628_9.INJECT1_1 = "NO";
    CCU2C add_7628_7 (.A0(n2567), .B0(n30902), .C0(n64_adj_315), .D0(n2142), 
          .A1(n2566), .B1(n30902), .C1(n64_adj_315), .D1(n2141), .CIN(n32512), 
          .COUT(n32513), .S0(n2720), .S1(n2719));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_7.INIT0 = 16'ha9aa;
    defparam add_7628_7.INIT1 = 16'ha9aa;
    defparam add_7628_7.INJECT1_0 = "NO";
    defparam add_7628_7.INJECT1_1 = "NO";
    CCU2C add_7628_5 (.A0(n2569), .B0(n30902), .C0(n64_adj_315), .D0(n42824), 
          .A1(n2568), .B1(n30902), .C1(n64_adj_315), .D1(n42822), .CIN(n32511), 
          .COUT(n32512), .S0(n2722), .S1(n2721));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_5.INIT0 = 16'ha9aa;
    defparam add_7628_5.INIT1 = 16'ha9aa;
    defparam add_7628_5.INJECT1_0 = "NO";
    defparam add_7628_5.INJECT1_1 = "NO";
    CCU2C add_7628_3 (.A0(n876), .B0(n30902), .C0(n64_adj_315), .D0(n42827), 
          .A1(n2570), .B1(n30902), .C1(n64_adj_315), .D1(n42823), .CIN(n32510), 
          .COUT(n32511), .S0(n2724), .S1(n2723));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_3.INIT0 = 16'ha9aa;
    defparam add_7628_3.INIT1 = 16'ha9aa;
    defparam add_7628_3.INJECT1_0 = "NO";
    defparam add_7628_3.INJECT1_1 = "NO";
    CCU2C add_7628_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_315), .B1(n30902), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32510));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7628_1.INIT0 = 16'h0000;
    defparam add_7628_1.INIT1 = 16'heee1;
    defparam add_7628_1.INJECT1_0 = "NO";
    defparam add_7628_1.INJECT1_1 = "NO";
    PFUMX div_4016_LessThan_1961_i62 (.BLUT(n58_adj_357), .ALUT(n60_adj_358), 
          .C0(n37885), .Z(n62_adj_359));
    FD1P3IX x_3___i79 (.D(n5511), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [14]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i79.GSR = "ENABLED";
    FD1P3IX x_3___i80 (.D(n5510), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [15]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i80.GSR = "ENABLED";
    FD1P3IX x_3___i81 (.D(n5509), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [16]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i81.GSR = "ENABLED";
    FD1P3IX x_3___i82 (.D(n5508), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [17]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i82.GSR = "ENABLED";
    FD1P3IX x_3___i83 (.D(n5507), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [18]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i83.GSR = "ENABLED";
    FD1P3IX x_3___i84 (.D(n5506), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [19]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i84.GSR = "ENABLED";
    FD1P3IX x_3___i85 (.D(n5505), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [20]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i85.GSR = "ENABLED";
    FD1P3IX x_3___i86 (.D(n5504), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [21]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i86.GSR = "ENABLED";
    FD1P3IX x_3___i87 (.D(n5503), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [22]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i87.GSR = "ENABLED";
    FD1P3IX x_3___i88 (.D(n5502), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [23]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i88.GSR = "ENABLED";
    FD1P3IX x_3___i89 (.D(n5501), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [24]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i89.GSR = "ENABLED";
    FD1P3IX x_3___i90 (.D(n5500), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [25]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i90.GSR = "ENABLED";
    FD1P3IX x_3___i91 (.D(n5499), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i91.GSR = "ENABLED";
    FD1P3IX x_3___i92 (.D(n5498), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i92.GSR = "ENABLED";
    FD1P3IX x_3___i93 (.D(n5497), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i93.GSR = "ENABLED";
    FD1P3IX x_3___i94 (.D(n5496), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i94.GSR = "ENABLED";
    FD1P3IX x_3___i95 (.D(n5495), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i95.GSR = "ENABLED";
    FD1P3IX x_3___i96 (.D(n5494), .SP(clk_c_enable_812), .CD(n31021), 
            .CK(clk_c), .Q(\x[1] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i96.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_1114 (.A(n113_adj_222), .B(n112_adj_221), .Z(n42813)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1114.init = 16'heeee;
    FD1P3IX x_3___i97 (.D(n5525), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i97.GSR = "ENABLED";
    FD1P3IX x_3___i98 (.D(n5524), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [1]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i98.GSR = "ENABLED";
    FD1P3IX x_3___i99 (.D(n5523), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [2]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i99.GSR = "ENABLED";
    FD1P3IX x_3___i100 (.D(n5522), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [3]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i100.GSR = "ENABLED";
    FD1P3IX x_3___i101 (.D(n5521), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [4]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i101.GSR = "ENABLED";
    FD1P3IX x_3___i102 (.D(n5520), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [5]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i102.GSR = "ENABLED";
    OB x_out_pad_41 (.I(x_out_c_41), .O(x_out[41]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_42 (.I(x_out_c_42), .O(x_out[42]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_43 (.I(x_out_c_43), .O(x_out[43]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_44 (.I(x_out_c_44), .O(x_out[44]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_45 (.I(x_out_c_45), .O(x_out[45]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7627_15 (.A0(n2402), .B0(n42789), .C0(n64_adj_301), .D0(n2455), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32506), 
          .S0(n2558));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_15.INIT0 = 16'ha9aa;
    defparam add_7627_15.INIT1 = 16'h0000;
    defparam add_7627_15.INJECT1_0 = "NO";
    defparam add_7627_15.INJECT1_1 = "NO";
    CCU2C add_7627_13 (.A0(n2404), .B0(n42789), .C0(n64_adj_301), .D0(n2298), 
          .A1(n2403), .B1(n42789), .C1(n64_adj_301), .D1(n2456), .CIN(n32505), 
          .COUT(n32506), .S0(n2560), .S1(n2559));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_13.INIT0 = 16'ha9aa;
    defparam add_7627_13.INIT1 = 16'ha9aa;
    defparam add_7627_13.INJECT1_0 = "NO";
    defparam add_7627_13.INJECT1_1 = "NO";
    CCU2C add_7627_11 (.A0(n2406), .B0(n42789), .C0(n64_adj_301), .D0(n1805), 
          .A1(n2405), .B1(n42789), .C1(n64_adj_301), .D1(n2137), .CIN(n32504), 
          .COUT(n32505), .S0(n2562), .S1(n2561));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_11.INIT0 = 16'ha9aa;
    defparam add_7627_11.INIT1 = 16'ha9aa;
    defparam add_7627_11.INJECT1_0 = "NO";
    defparam add_7627_11.INJECT1_1 = "NO";
    CCU2C add_7627_9 (.A0(n2408), .B0(n42789), .C0(n64_adj_301), .D0(n1462), 
          .A1(n2407), .B1(n42789), .C1(n64_adj_301), .D1(n1635), .CIN(n32503), 
          .COUT(n32504), .S0(n2564), .S1(n2563));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_9.INIT0 = 16'ha9aa;
    defparam add_7627_9.INIT1 = 16'ha9aa;
    defparam add_7627_9.INJECT1_0 = "NO";
    defparam add_7627_9.INJECT1_1 = "NO";
    CCU2C add_7627_7 (.A0(n2410), .B0(n42789), .C0(n64_adj_301), .D0(n2142), 
          .A1(n2409), .B1(n42789), .C1(n64_adj_301), .D1(n2141), .CIN(n32502), 
          .COUT(n32503), .S0(n2566), .S1(n2565));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_7.INIT0 = 16'ha9aa;
    defparam add_7627_7.INIT1 = 16'ha9aa;
    defparam add_7627_7.INJECT1_0 = "NO";
    defparam add_7627_7.INJECT1_1 = "NO";
    CCU2C add_7627_5 (.A0(n2412), .B0(n42789), .C0(n64_adj_301), .D0(n42824), 
          .A1(n2411), .B1(n42789), .C1(n64_adj_301), .D1(n42822), .CIN(n32501), 
          .COUT(n32502), .S0(n2568), .S1(n2567));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_5.INIT0 = 16'ha9aa;
    defparam add_7627_5.INIT1 = 16'ha9aa;
    defparam add_7627_5.INJECT1_0 = "NO";
    defparam add_7627_5.INJECT1_1 = "NO";
    CCU2C add_7627_3 (.A0(n875), .B0(n42789), .C0(n64_adj_301), .D0(n42827), 
          .A1(n2413), .B1(n42789), .C1(n64_adj_301), .D1(n42823), .CIN(n32500), 
          .COUT(n32501), .S0(n2570), .S1(n2569));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_3.INIT0 = 16'ha9aa;
    defparam add_7627_3.INIT1 = 16'ha9aa;
    defparam add_7627_3.INJECT1_0 = "NO";
    defparam add_7627_3.INJECT1_1 = "NO";
    CCU2C add_7627_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_301), .B1(n42789), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32500));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7627_1.INIT0 = 16'h0000;
    defparam add_7627_1.INIT1 = 16'heee1;
    defparam add_7627_1.INJECT1_0 = "NO";
    defparam add_7627_1.INJECT1_1 = "NO";
    CCU2C add_7626_13 (.A0(n2244), .B0(n30896), .C0(n64_adj_289), .D0(n2298), 
          .A1(n2243), .B1(n30896), .C1(n64_adj_289), .D1(n2456), .CIN(n32495), 
          .S0(n2403), .S1(n2402));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_13.INIT0 = 16'ha9aa;
    defparam add_7626_13.INIT1 = 16'ha9aa;
    defparam add_7626_13.INJECT1_0 = "NO";
    defparam add_7626_13.INJECT1_1 = "NO";
    CCU2C add_7626_11 (.A0(n2246), .B0(n30896), .C0(n64_adj_289), .D0(n1805), 
          .A1(n2245), .B1(n30896), .C1(n64_adj_289), .D1(n2137), .CIN(n32494), 
          .COUT(n32495), .S0(n2405), .S1(n2404));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_11.INIT0 = 16'ha9aa;
    defparam add_7626_11.INIT1 = 16'ha9aa;
    defparam add_7626_11.INJECT1_0 = "NO";
    defparam add_7626_11.INJECT1_1 = "NO";
    CCU2C add_7626_9 (.A0(n2248), .B0(n30896), .C0(n64_adj_289), .D0(n1462), 
          .A1(n2247), .B1(n30896), .C1(n64_adj_289), .D1(n1635), .CIN(n32493), 
          .COUT(n32494), .S0(n2407), .S1(n2406));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_9.INIT0 = 16'ha9aa;
    defparam add_7626_9.INIT1 = 16'ha9aa;
    defparam add_7626_9.INJECT1_0 = "NO";
    defparam add_7626_9.INJECT1_1 = "NO";
    CCU2C add_7626_7 (.A0(n2250), .B0(n30896), .C0(n64_adj_289), .D0(n2142), 
          .A1(n2249), .B1(n30896), .C1(n64_adj_289), .D1(n2141), .CIN(n32492), 
          .COUT(n32493), .S0(n2409), .S1(n2408));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_7.INIT0 = 16'ha9aa;
    defparam add_7626_7.INIT1 = 16'ha9aa;
    defparam add_7626_7.INJECT1_0 = "NO";
    defparam add_7626_7.INJECT1_1 = "NO";
    CCU2C add_7626_5 (.A0(n2252), .B0(n30896), .C0(n64_adj_289), .D0(n42824), 
          .A1(n2251), .B1(n30896), .C1(n64_adj_289), .D1(n42822), .CIN(n32491), 
          .COUT(n32492), .S0(n2411), .S1(n2410));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_5.INIT0 = 16'ha9aa;
    defparam add_7626_5.INIT1 = 16'ha9aa;
    defparam add_7626_5.INJECT1_0 = "NO";
    defparam add_7626_5.INJECT1_1 = "NO";
    CCU2C add_7626_3 (.A0(n874), .B0(n30896), .C0(n64_adj_289), .D0(n42827), 
          .A1(n2253), .B1(n30896), .C1(n64_adj_289), .D1(n42823), .CIN(n32490), 
          .COUT(n32491), .S0(n2413), .S1(n2412));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_3.INIT0 = 16'ha9aa;
    defparam add_7626_3.INIT1 = 16'ha9aa;
    defparam add_7626_3.INJECT1_0 = "NO";
    defparam add_7626_3.INJECT1_1 = "NO";
    CCU2C add_7626_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_289), .B1(n30896), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32490));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7626_1.INIT0 = 16'h0000;
    defparam add_7626_1.INIT1 = 16'heee1;
    defparam add_7626_1.INJECT1_0 = "NO";
    defparam add_7626_1.INJECT1_1 = "NO";
    CCU2C add_7625_13 (.A0(n2081), .B0(n30893), .C0(n64_adj_278), .D0(n2298), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32486), 
          .S0(n2243));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_13.INIT0 = 16'ha9aa;
    defparam add_7625_13.INIT1 = 16'h0000;
    defparam add_7625_13.INJECT1_0 = "NO";
    defparam add_7625_13.INJECT1_1 = "NO";
    CCU2C add_7625_11 (.A0(n2083), .B0(n30893), .C0(n64_adj_278), .D0(n1805), 
          .A1(n2082), .B1(n30893), .C1(n64_adj_278), .D1(n2137), .CIN(n32485), 
          .COUT(n32486), .S0(n2245), .S1(n2244));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_11.INIT0 = 16'ha9aa;
    defparam add_7625_11.INIT1 = 16'ha9aa;
    defparam add_7625_11.INJECT1_0 = "NO";
    defparam add_7625_11.INJECT1_1 = "NO";
    CCU2C add_7625_9 (.A0(n2085), .B0(n30893), .C0(n64_adj_278), .D0(n1462), 
          .A1(n2084), .B1(n30893), .C1(n64_adj_278), .D1(n1635), .CIN(n32484), 
          .COUT(n32485), .S0(n2247), .S1(n2246));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_9.INIT0 = 16'ha9aa;
    defparam add_7625_9.INIT1 = 16'ha9aa;
    defparam add_7625_9.INJECT1_0 = "NO";
    defparam add_7625_9.INJECT1_1 = "NO";
    CCU2C add_7625_7 (.A0(n2087), .B0(n30893), .C0(n64_adj_278), .D0(n2142), 
          .A1(n2086), .B1(n30893), .C1(n64_adj_278), .D1(n2141), .CIN(n32483), 
          .COUT(n32484), .S0(n2249), .S1(n2248));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_7.INIT0 = 16'ha9aa;
    defparam add_7625_7.INIT1 = 16'ha9aa;
    defparam add_7625_7.INJECT1_0 = "NO";
    defparam add_7625_7.INJECT1_1 = "NO";
    CCU2C add_7625_5 (.A0(n2089), .B0(n30893), .C0(n64_adj_278), .D0(n42824), 
          .A1(n2088), .B1(n30893), .C1(n64_adj_278), .D1(n42822), .CIN(n32482), 
          .COUT(n32483), .S0(n2251), .S1(n2250));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_5.INIT0 = 16'ha9aa;
    defparam add_7625_5.INIT1 = 16'ha9aa;
    defparam add_7625_5.INJECT1_0 = "NO";
    defparam add_7625_5.INJECT1_1 = "NO";
    CCU2C add_7625_3 (.A0(n873), .B0(n30893), .C0(n64_adj_278), .D0(n42827), 
          .A1(n2090), .B1(n30893), .C1(n64_adj_278), .D1(n42823), .CIN(n32481), 
          .COUT(n32482), .S0(n2253), .S1(n2252));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_3.INIT0 = 16'ha9aa;
    defparam add_7625_3.INIT1 = 16'ha9aa;
    defparam add_7625_3.INJECT1_0 = "NO";
    defparam add_7625_3.INJECT1_1 = "NO";
    CCU2C add_7625_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_278), .B1(n30893), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32481));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7625_1.INIT0 = 16'h0000;
    defparam add_7625_1.INIT1 = 16'heee1;
    defparam add_7625_1.INJECT1_0 = "NO";
    defparam add_7625_1.INJECT1_1 = "NO";
    LUT4 div_4016_LessThan_1961_i34_4_lut (.A(n132), .B(n131_adj_234), .C(n3023), 
         .D(n879), .Z(n34)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i34_4_lut.init = 16'h0c8e;
    LUT4 i1_2_lut_3_lut_4_lut_adj_56 (.A(n113_adj_222), .B(n112_adj_221), 
         .C(n36948), .D(n42816), .Z(n36882)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_56.init = 16'hfffe;
    FD1P3IX x_3___i103 (.D(n5519), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [6]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i103.GSR = "ENABLED";
    FD1P3IX x_3___i104 (.D(n5518), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [7]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i104.GSR = "ENABLED";
    FD1P3IX x_3___i105 (.D(n5517), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [8]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i105.GSR = "ENABLED";
    FD1P3IX x_3___i106 (.D(n5516), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [9]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i106.GSR = "ENABLED";
    FD1P3IX x_3___i123 (.D(n5499), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [26]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i123.GSR = "ENABLED";
    FD1P3IX x_3___i124 (.D(n5498), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [27]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i124.GSR = "ENABLED";
    FD1P3AX U_15___i509 (.D(\U[0] [28]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i509.GSR = "ENABLED";
    LUT4 div_4016_LessThan_2513_i38_3_lut_3_lut (.A(n3837), .B(n120), .C(n36_adj_478), 
         .Z(n38_adj_479)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_rep_1107_3_lut_4_lut (.A(n113_adj_222), .B(n112_adj_221), 
         .C(n110_adj_220), .D(n111), .Z(n42806)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1107_3_lut_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i24_3_lut_3_lut (.A(n4663), .B(n120), .C(n22_adj_680), 
         .Z(n24_adj_681)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3137_i21_2_lut (.A(n4772), .B(n123), .Z(n21_adj_714)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i21_2_lut.init = 16'h6666;
    OB x_out_pad_46 (.I(x_out_c_46), .O(x_out[46]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_47 (.I(x_out_c_47), .O(x_out[47]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_48 (.I(x_out_c_48), .O(x_out[48]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_49 (.I(x_out_c_49), .O(x_out[49]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7624_11 (.A0(n1917), .B0(n30890), .C0(n64_adj_269), .D0(n1805), 
          .A1(n1916), .B1(n30890), .C1(n64_adj_269), .D1(n2137), .CIN(n32476), 
          .S0(n2082), .S1(n2081));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7624_11.INIT0 = 16'ha9aa;
    defparam add_7624_11.INIT1 = 16'ha9aa;
    defparam add_7624_11.INJECT1_0 = "NO";
    defparam add_7624_11.INJECT1_1 = "NO";
    CCU2C add_7624_9 (.A0(n1919), .B0(n30890), .C0(n64_adj_269), .D0(n1462), 
          .A1(n1918), .B1(n30890), .C1(n64_adj_269), .D1(n1635), .CIN(n32475), 
          .COUT(n32476), .S0(n2084), .S1(n2083));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7624_9.INIT0 = 16'ha9aa;
    defparam add_7624_9.INIT1 = 16'ha9aa;
    defparam add_7624_9.INJECT1_0 = "NO";
    defparam add_7624_9.INJECT1_1 = "NO";
    CCU2C add_7624_7 (.A0(n1921), .B0(n30890), .C0(n64_adj_269), .D0(n2142), 
          .A1(n1920), .B1(n30890), .C1(n64_adj_269), .D1(n2141), .CIN(n32474), 
          .COUT(n32475), .S0(n2086), .S1(n2085));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7624_7.INIT0 = 16'ha9aa;
    defparam add_7624_7.INIT1 = 16'ha9aa;
    defparam add_7624_7.INJECT1_0 = "NO";
    defparam add_7624_7.INJECT1_1 = "NO";
    CCU2C add_7624_5 (.A0(n1923), .B0(n30890), .C0(n64_adj_269), .D0(n42824), 
          .A1(n1922), .B1(n30890), .C1(n64_adj_269), .D1(n42822), .CIN(n32473), 
          .COUT(n32474), .S0(n2088), .S1(n2087));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7624_5.INIT0 = 16'ha9aa;
    defparam add_7624_5.INIT1 = 16'ha9aa;
    defparam add_7624_5.INJECT1_0 = "NO";
    defparam add_7624_5.INJECT1_1 = "NO";
    CCU2C add_7624_3 (.A0(n872), .B0(n30890), .C0(n64_adj_269), .D0(n42827), 
          .A1(n1924), .B1(n30890), .C1(n64_adj_269), .D1(n42823), .CIN(n32472), 
          .COUT(n32473), .S0(n2090), .S1(n2089));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7624_3.INIT0 = 16'ha9aa;
    defparam add_7624_3.INIT1 = 16'ha9aa;
    defparam add_7624_3.INJECT1_0 = "NO";
    defparam add_7624_3.INJECT1_1 = "NO";
    CCU2C add_7624_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_269), .B1(n30890), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32472));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7624_1.INIT0 = 16'h0000;
    defparam add_7624_1.INIT1 = 16'heee1;
    defparam add_7624_1.INJECT1_0 = "NO";
    defparam add_7624_1.INJECT1_1 = "NO";
    CCU2C add_7623_11 (.A0(n1748), .B0(n30887), .C0(n64_adj_260), .D0(n1805), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32468), 
          .S0(n1916));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7623_11.INIT0 = 16'ha9aa;
    defparam add_7623_11.INIT1 = 16'h0000;
    defparam add_7623_11.INJECT1_0 = "NO";
    defparam add_7623_11.INJECT1_1 = "NO";
    CCU2C add_7623_9 (.A0(n1750), .B0(n30887), .C0(n64_adj_260), .D0(n1462), 
          .A1(n1749), .B1(n30887), .C1(n64_adj_260), .D1(n1635), .CIN(n32467), 
          .COUT(n32468), .S0(n1918), .S1(n1917));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7623_9.INIT0 = 16'ha9aa;
    defparam add_7623_9.INIT1 = 16'ha9aa;
    defparam add_7623_9.INJECT1_0 = "NO";
    defparam add_7623_9.INJECT1_1 = "NO";
    CCU2C add_7623_7 (.A0(n1752), .B0(n30887), .C0(n64_adj_260), .D0(n2142), 
          .A1(n1751), .B1(n30887), .C1(n64_adj_260), .D1(n2141), .CIN(n32466), 
          .COUT(n32467), .S0(n1920), .S1(n1919));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7623_7.INIT0 = 16'ha9aa;
    defparam add_7623_7.INIT1 = 16'ha9aa;
    defparam add_7623_7.INJECT1_0 = "NO";
    defparam add_7623_7.INJECT1_1 = "NO";
    CCU2C add_7623_5 (.A0(n1754), .B0(n30887), .C0(n64_adj_260), .D0(n42824), 
          .A1(n1753), .B1(n30887), .C1(n64_adj_260), .D1(n42822), .CIN(n32465), 
          .COUT(n32466), .S0(n1922), .S1(n1921));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7623_5.INIT0 = 16'ha9aa;
    defparam add_7623_5.INIT1 = 16'ha9aa;
    defparam add_7623_5.INJECT1_0 = "NO";
    defparam add_7623_5.INJECT1_1 = "NO";
    CCU2C add_7623_3 (.A0(n685), .B0(n30887), .C0(n64_adj_260), .D0(n42827), 
          .A1(n1755), .B1(n30887), .C1(n64_adj_260), .D1(n42823), .CIN(n32464), 
          .COUT(n32465), .S0(n1924), .S1(n1923));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7623_3.INIT0 = 16'ha9aa;
    defparam add_7623_3.INIT1 = 16'ha9aa;
    defparam add_7623_3.INJECT1_0 = "NO";
    defparam add_7623_3.INJECT1_1 = "NO";
    CCU2C add_7623_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_260), .B1(n30887), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32464));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7623_1.INIT0 = 16'h0000;
    defparam add_7623_1.INIT1 = 16'heee1;
    defparam add_7623_1.INJECT1_0 = "NO";
    defparam add_7623_1.INJECT1_1 = "NO";
    CCU2C add_7622_9 (.A0(n1578), .B0(n30884), .C0(n64_adj_252), .D0(n1462), 
          .A1(n1577), .B1(n30884), .C1(n64_adj_252), .D1(n1635), .CIN(n32459), 
          .S0(n1749), .S1(n1748));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7622_9.INIT0 = 16'ha9aa;
    defparam add_7622_9.INIT1 = 16'ha9aa;
    defparam add_7622_9.INJECT1_0 = "NO";
    defparam add_7622_9.INJECT1_1 = "NO";
    CCU2C add_7622_7 (.A0(n1580), .B0(n30884), .C0(n64_adj_252), .D0(n2142), 
          .A1(n1579), .B1(n30884), .C1(n64_adj_252), .D1(n2141), .CIN(n32458), 
          .COUT(n32459), .S0(n1751), .S1(n1750));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7622_7.INIT0 = 16'ha9aa;
    defparam add_7622_7.INIT1 = 16'ha9aa;
    defparam add_7622_7.INJECT1_0 = "NO";
    defparam add_7622_7.INJECT1_1 = "NO";
    CCU2C add_7622_5 (.A0(n1582), .B0(n30884), .C0(n64_adj_252), .D0(n42824), 
          .A1(n1581), .B1(n30884), .C1(n64_adj_252), .D1(n42822), .CIN(n32457), 
          .COUT(n32458), .S0(n1753), .S1(n1752));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7622_5.INIT0 = 16'ha9aa;
    defparam add_7622_5.INIT1 = 16'ha9aa;
    defparam add_7622_5.INJECT1_0 = "NO";
    defparam add_7622_5.INJECT1_1 = "NO";
    CCU2C add_7622_3 (.A0(n684), .B0(n30884), .C0(n64_adj_252), .D0(n42827), 
          .A1(n1583), .B1(n30884), .C1(n64_adj_252), .D1(n42823), .CIN(n32456), 
          .COUT(n32457), .S0(n1755), .S1(n1754));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7622_3.INIT0 = 16'ha9aa;
    defparam add_7622_3.INIT1 = 16'ha9aa;
    defparam add_7622_3.INJECT1_0 = "NO";
    defparam add_7622_3.INJECT1_1 = "NO";
    CCU2C add_7622_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_252), .B1(n30884), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32456));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7622_1.INIT0 = 16'h0000;
    defparam add_7622_1.INIT1 = 16'heee1;
    defparam add_7622_1.INJECT1_0 = "NO";
    defparam add_7622_1.INJECT1_1 = "NO";
    CCU2C add_7621_9 (.A0(n1403), .B0(n30881), .C0(n64_adj_246), .D0(n1462), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32452), 
          .S0(n1577));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7621_9.INIT0 = 16'ha9aa;
    defparam add_7621_9.INIT1 = 16'h0000;
    defparam add_7621_9.INJECT1_0 = "NO";
    defparam add_7621_9.INJECT1_1 = "NO";
    CCU2C add_7621_7 (.A0(n1405), .B0(n30881), .C0(n64_adj_246), .D0(n2142), 
          .A1(n1404), .B1(n30881), .C1(n64_adj_246), .D1(n2141), .CIN(n32451), 
          .COUT(n32452), .S0(n1579), .S1(n1578));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7621_7.INIT0 = 16'ha9aa;
    defparam add_7621_7.INIT1 = 16'ha9aa;
    defparam add_7621_7.INJECT1_0 = "NO";
    defparam add_7621_7.INJECT1_1 = "NO";
    CCU2C add_7621_5 (.A0(n1407), .B0(n30881), .C0(n64_adj_246), .D0(n42824), 
          .A1(n1406), .B1(n30881), .C1(n64_adj_246), .D1(n42822), .CIN(n32450), 
          .COUT(n32451), .S0(n1581), .S1(n1580));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7621_5.INIT0 = 16'ha9aa;
    defparam add_7621_5.INIT1 = 16'ha9aa;
    defparam add_7621_5.INJECT1_0 = "NO";
    defparam add_7621_5.INJECT1_1 = "NO";
    CCU2C add_7621_3 (.A0(n683), .B0(n30881), .C0(n64_adj_246), .D0(n42827), 
          .A1(n1408), .B1(n30881), .C1(n64_adj_246), .D1(n42823), .CIN(n32449), 
          .COUT(n32450), .S0(n1583), .S1(n1582));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7621_3.INIT0 = 16'ha9aa;
    defparam add_7621_3.INIT1 = 16'ha9aa;
    defparam add_7621_3.INJECT1_0 = "NO";
    defparam add_7621_3.INJECT1_1 = "NO";
    CCU2C add_7621_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_246), .B1(n30881), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32449));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7621_1.INIT0 = 16'h0000;
    defparam add_7621_1.INIT1 = 16'heee1;
    defparam add_7621_1.INJECT1_0 = "NO";
    defparam add_7621_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1116 (.A(n114), .B(n117), .Z(n42815)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1116.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_57 (.A(n114), .B(n117), .C(n118_adj_225), 
         .D(n116_adj_224), .Z(n37272)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_57.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i23_2_lut_rep_783 (.A(n4666), .B(n123), 
         .Z(n42482)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i23_2_lut_rep_783.init = 16'h6666;
    LUT4 i1_2_lut_rep_1117 (.A(n115_adj_223), .B(n114), .Z(n42816)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1117.init = 16'heeee;
    LUT4 div_4016_LessThan_2513_i41_2_lut_rep_913 (.A(n3838), .B(n121_adj_227), 
         .Z(n42612)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i41_2_lut_rep_913.init = 16'h6666;
    LUT4 div_4016_i3319_4_lut (.A(n64_adj_260), .B(n22283), .C(n42786), 
         .D(n30887), .Z(n5502)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3319_4_lut.init = 16'hc0c5;
    OB x_out_pad_50 (.I(x_out_c_50), .O(x_out[50]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_51 (.I(x_out_c_51), .O(x_out[51]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_52 (.I(x_out_c_52), .O(x_out[52]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C add_7620_7 (.A0(n1227), .B0(n30878), .C0(n64_adj_241), .D0(n2142), 
          .A1(n35972), .B1(n30878), .C1(n64_adj_241), .D1(n2141), .CIN(n32444), 
          .S0(n1404), .S1(n1403));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7620_7.INIT0 = 16'ha9aa;
    defparam add_7620_7.INIT1 = 16'ha9aa;
    defparam add_7620_7.INJECT1_0 = "NO";
    defparam add_7620_7.INJECT1_1 = "NO";
    CCU2C add_7620_5 (.A0(n1229), .B0(n30878), .C0(n64_adj_241), .D0(n42824), 
          .A1(n1228), .B1(n30878), .C1(n64_adj_241), .D1(n42822), .CIN(n32443), 
          .COUT(n32444), .S0(n1406), .S1(n1405));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7620_5.INIT0 = 16'ha9aa;
    defparam add_7620_5.INIT1 = 16'ha9aa;
    defparam add_7620_5.INJECT1_0 = "NO";
    defparam add_7620_5.INJECT1_1 = "NO";
    CCU2C add_7620_3 (.A0(n682), .B0(n30878), .C0(n64_adj_241), .D0(n42827), 
          .A1(n1230), .B1(n30878), .C1(n64_adj_241), .D1(n42823), .CIN(n32442), 
          .COUT(n32443), .S0(n1408), .S1(n1407));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7620_3.INIT0 = 16'ha9aa;
    defparam add_7620_3.INIT1 = 16'ha9aa;
    defparam add_7620_3.INJECT1_0 = "NO";
    defparam add_7620_3.INJECT1_1 = "NO";
    CCU2C add_7620_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n64_adj_241), .B1(n30878), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32442));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam add_7620_1.INIT0 = 16'h0000;
    defparam add_7620_1.INIT1 = 16'heee1;
    defparam add_7620_1.INJECT1_0 = "NO";
    defparam add_7620_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_34 (.A0(i[31]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n32438), 
          .S0(n70));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_34.INIT0 = 16'h555f;
    defparam _add_1_add_4_34.INIT1 = 16'h0000;
    defparam _add_1_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_32 (.A0(i[29]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[30]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32437), 
          .COUT(n32438), .S0(n76_adj_101), .S1(n73_adj_95));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_32.INIT0 = 16'h555f;
    defparam _add_1_add_4_32.INIT1 = 16'h555f;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_30 (.A0(i[27]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[28]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32436), 
          .COUT(n32437), .S0(n82_adj_104), .S1(n79_adj_98));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_30.INIT0 = 16'h555f;
    defparam _add_1_add_4_30.INIT1 = 16'h555f;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(i[25]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[26]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32435), 
          .COUT(n32436), .S0(n88_adj_151), .S1(n85_adj_91));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_28.INIT0 = 16'h555f;
    defparam _add_1_add_4_28.INIT1 = 16'h555f;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(i[23]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[24]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32434), 
          .COUT(n32435), .S0(n94_adj_152), .S1(n91_adj_160));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_26.INIT0 = 16'h555f;
    defparam _add_1_add_4_26.INIT1 = 16'h555f;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_24 (.A0(i[21]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[22]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32433), 
          .COUT(n32434), .S0(n100_adj_161), .S1(n97_adj_153));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_24.INIT0 = 16'h555f;
    defparam _add_1_add_4_24.INIT1 = 16'h555f;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_22 (.A0(i[19]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[20]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32432), 
          .COUT(n32433), .S0(n106_adj_49), .S1(n103_adj_92));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_22.INIT0 = 16'h555f;
    defparam _add_1_add_4_22.INIT1 = 16'h555f;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_20 (.A0(i[17]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[18]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32431), 
          .COUT(n32432), .S0(n112_adj_50), .S1(n109_adj_106));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_20.INIT0 = 16'h555f;
    defparam _add_1_add_4_20.INIT1 = 16'h555f;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_18 (.A0(i[15]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32430), 
          .COUT(n32431), .S0(n118_adj_100), .S1(n115_adj_52));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_18.INIT0 = 16'h555f;
    defparam _add_1_add_4_18.INIT1 = 16'h555f;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_16 (.A0(i[13]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32429), 
          .COUT(n32430), .S0(n124_adj_154), .S1(n121_adj_150));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_14 (.A0(i[11]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32428), 
          .COUT(n32429), .S0(n130_adj_99), .S1(n127_adj_102));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_12 (.A0(i[9]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32427), 
          .COUT(n32428), .S0(n136_adj_53), .S1(n133_adj_90));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_10 (.A0(i[7]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32426), 
          .COUT(n32427), .S0(n142_adj_96), .S1(n139_adj_94));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_8 (.A0(i[5]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32425), 
          .COUT(n32426), .S0(n148_adj_113), .S1(n145_adj_103));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_8.INIT0 = 16'h555f;
    defparam _add_1_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_6 (.A0(i[3]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32424), 
          .COUT(n32425), .S0(n154_adj_158), .S1(n151_adj_159));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_6.INIT0 = 16'h555f;
    defparam _add_1_add_4_6.INIT1 = 16'h555f;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_4 (.A0(i[1]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(i[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n32423), 
          .COUT(n32424), .S0(n160_adj_156), .S1(n157_adj_157));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_4.INIT0 = 16'h555f;
    defparam _add_1_add_4_4.INIT1 = 16'h555f;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n16519), .B1(i[0]), .C1(GND_net), .D1(VCC_net), .COUT(n32423), 
          .S1(n163_adj_155));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(122[18:23])
    defparam _add_1_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_34 (.A0(n25244), .B0(\y[3] [31]), .C0(i[0]), 
          .D0(i[1]), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32422), .S0(n70_adj_87));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_34.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_34.INIT1 = 16'h0000;
    defparam _add_1_7038_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_32 (.A0(n25248), .B0(\y[3] [29]), .C0(i[0]), 
          .D0(i[1]), .A1(n25246), .B1(\y[3] [30]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32421), .COUT(n32422), .S0(n76), .S1(n73));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_32.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_32.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_30 (.A0(n25252), .B0(\y[3] [27]), .C0(i[0]), 
          .D0(i[1]), .A1(n25250), .B1(\y[3] [28]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32420), .COUT(n32421), .S0(n82), .S1(n79));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_30.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_30.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_28 (.A0(n25256), .B0(\y[3] [25]), .C0(i[0]), 
          .D0(i[1]), .A1(n25254), .B1(\y[3] [26]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32419), .COUT(n32420), .S0(n88), .S1(n85));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_28.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_28.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_26 (.A0(n25260), .B0(\y[3] [23]), .C0(i[0]), 
          .D0(i[1]), .A1(n25258), .B1(\y[3] [24]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32418), .COUT(n32419), .S0(n94), .S1(n91));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_26.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_26.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_24 (.A0(n25264), .B0(\y[3] [21]), .C0(i[0]), 
          .D0(i[1]), .A1(n25262), .B1(\y[3] [22]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32417), .COUT(n32418), .S0(n100), .S1(n97));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_24.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_24.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_22 (.A0(n25268), .B0(\y[3] [19]), .C0(i[0]), 
          .D0(i[1]), .A1(n25266), .B1(\y[3] [20]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32416), .COUT(n32417), .S0(n106), .S1(n103));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_22.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_22.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_22.INJECT1_1 = "NO";
    LUT4 i24126_3_lut_4_lut (.A(n4666), .B(n123), .C(n13_adj_674), .D(n42483), 
         .Z(n39386)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24126_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_3137_i17_2_lut (.A(n4774), .B(n125_adj_230), 
         .Z(n17_adj_711)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i17_2_lut.init = 16'h6666;
    PFUMX div_4016_LessThan_1961_i54 (.BLUT(n46_adj_351), .ALUT(n52_adj_354), 
          .C0(n37859), .Z(n54_adj_355));
    OB x_out_pad_53 (.I(x_out_c_53), .O(x_out[53]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_54 (.I(x_out_c_54), .O(x_out[54]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    CCU2C _add_1_7038_add_4_20 (.A0(n25272), .B0(\y[3] [17]), .C0(i[0]), 
          .D0(i[1]), .A1(n25270), .B1(\y[3] [18]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32415), .COUT(n32416), .S0(n112), .S1(n109));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_20.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_20.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_18 (.A0(n25276), .B0(\y[3] [15]), .C0(i[0]), 
          .D0(i[1]), .A1(n25274), .B1(\y[3] [16]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32414), .COUT(n32415), .S0(n118), .S1(n115));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_18.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_18.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_16 (.A0(n25280), .B0(\y[3] [13]), .C0(i[0]), 
          .D0(i[1]), .A1(n25278), .B1(\y[3] [14]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32413), .COUT(n32414), .S0(n124), .S1(n121));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_16.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_16.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_14 (.A0(n25284), .B0(\y[3] [11]), .C0(i[0]), 
          .D0(i[1]), .A1(n25282), .B1(\y[3] [12]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32412), .COUT(n32413), .S0(n130), .S1(n127));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_14.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_14.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_12 (.A0(n25288), .B0(\y[3] [9]), .C0(i[0]), 
          .D0(i[1]), .A1(n25286), .B1(\y[3] [10]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32411), .COUT(n32412), .S0(n136), .S1(n133));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_12.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_12.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_10 (.A0(n25292), .B0(\y[3] [7]), .C0(i[0]), 
          .D0(i[1]), .A1(n25290), .B1(\y[3] [8]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32410), .COUT(n32411), .S0(n142), .S1(n139));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_10.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_10.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_8 (.A0(n25296), .B0(\y[3] [5]), .C0(i[0]), 
          .D0(i[1]), .A1(n25294), .B1(\y[3] [6]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32409), .COUT(n32410), .S0(n148), .S1(n145));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_8.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_8.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_6 (.A0(n25300), .B0(\y[3] [3]), .C0(i[0]), 
          .D0(i[1]), .A1(n25298), .B1(\y[3] [4]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32408), .COUT(n32409), .S0(n154), .S1(n151));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_6.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_6.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_4 (.A0(n25304), .B0(\y[3] [1]), .C0(i[0]), 
          .D0(i[1]), .A1(n25302), .B1(\y[3] [2]), .C1(i[0]), .D1(i[1]), 
          .CIN(n32407), .COUT(n32408), .S0(n160), .S1(n157));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_4.INIT0 = 16'h9555;
    defparam _add_1_7038_add_4_4.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_7038_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n25306), .B1(\y[3] [0]), .C1(i[0]), .D1(i[1]), 
          .COUT(n32407), .S1(n163_adj_11));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(108[14] 112[8])
    defparam _add_1_7038_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_7038_add_4_2.INIT1 = 16'h9555;
    defparam _add_1_7038_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_7038_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_33 (.A0(n164_adj_97), .B0(n63), .C0(n5194), 
          .D0(n164_adj_28), .A1(n163_adj_107), .B1(n63), .C1(n5193), 
          .D1(n163_adj_27), .CIN(n32405), .S0(n71), .S1(n68));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_31 (.A0(n166_adj_33), .B0(n63), .C0(n5196), 
          .D0(n166_adj_144), .A1(n165_adj_105), .B1(n63), .C1(n5195), 
          .D1(n165_adj_145), .CIN(n32404), .COUT(n32405), .S0(n77), 
          .S1(n74));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_29 (.A0(n168_adj_46), .B0(n63), .C0(n5198), 
          .D0(n168_adj_25), .A1(n167_adj_32), .B1(n63), .C1(n5197), 
          .D1(n167_adj_34), .CIN(n32403), .COUT(n32404), .S0(n83), .S1(n80));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_27 (.A0(n170_adj_43), .B0(n63), .C0(n5200), 
          .D0(n170_adj_139), .A1(n169_adj_37), .B1(n63), .C1(n5199), 
          .D1(n169_adj_26), .CIN(n32402), .COUT(n32403), .S0(n89), .S1(n86));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_25 (.A0(n172_adj_45), .B0(n63), .C0(n5202), 
          .D0(n172), .A1(n171_adj_36), .B1(n63), .C1(n5201), .D1(n171_adj_138), 
          .CIN(n32401), .COUT(n32402), .S0(n95), .S1(n92));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_23 (.A0(n174_adj_29), .B0(n63), .C0(n5204), 
          .D0(n174_adj_23), .A1(n173_adj_30), .B1(n63), .C1(n5203), 
          .D1(n173_adj_22), .CIN(n32400), .COUT(n32401), .S0(n101), 
          .S1(n98));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_21 (.A0(n176_adj_41), .B0(n63), .C0(n5206), 
          .D0(n176_adj_133), .A1(n175_adj_38), .B1(n63), .C1(n5205), 
          .D1(n175_adj_24), .CIN(n32399), .COUT(n32400), .S0(n107), 
          .S1(n104));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_19 (.A0(n178_adj_39), .B0(n63), .C0(n5208), 
          .D0(n178_adj_4), .A1(n177_adj_40), .B1(n63), .C1(n5207), .D1(n177_adj_132), 
          .CIN(n32398), .COUT(n32399), .S0(n113), .S1(n110));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_17 (.A0(n180_adj_88), .B0(n63), .C0(n5210), 
          .D0(n180_adj_20), .A1(n179_adj_89), .B1(n63), .C1(n5209), 
          .D1(n179_adj_19), .CIN(n32397), .COUT(n32398), .S0(n119), 
          .S1(n116));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_15 (.A0(n182_adj_112), .B0(n63), .C0(n5212), 
          .D0(n182_adj_127), .A1(n181_adj_31), .B1(n63), .C1(n5211), 
          .D1(n181_adj_21), .CIN(n32396), .COUT(n32397), .S0(n125), 
          .S1(n122));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_13 (.A0(n184_adj_110), .B0(n63), .C0(n5214), 
          .D0(n184_adj_6), .A1(n183_adj_111), .B1(n63), .C1(n5213), 
          .D1(n183_adj_126), .CIN(n32395), .COUT(n32396), .S0(n131), 
          .S1(n128));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_11 (.A0(n186_adj_108), .B0(n63), .C0(n5216), 
          .D0(n186_adj_17), .A1(n185_adj_109), .B1(n63), .C1(n5215), 
          .D1(n185_adj_16), .CIN(n32394), .COUT(n32395), .S0(n137), 
          .S1(n134));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_9 (.A0(n188_adj_93), .B0(n63), .C0(n5218), 
          .D0(n188_adj_121), .A1(n187_adj_51), .B1(n63), .C1(n5217), 
          .D1(n187_adj_18), .CIN(n32393), .COUT(n32394), .S0(n143), 
          .S1(n140));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_7 (.A0(n190_adj_35), .B0(n63), .C0(n5220), 
          .D0(n190_adj_7), .A1(n189_adj_86), .B1(n63), .C1(n5219), .D1(n189_adj_120), 
          .CIN(n32392), .COUT(n32393), .S0(n149), .S1(n146));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_5 (.A0(n192_adj_42), .B0(n63), .C0(n5222), 
          .D0(n192_adj_14), .A1(n191_adj_47), .B1(n63), .C1(n5221), 
          .D1(n191_adj_13), .CIN(n32391), .COUT(n32392), .S0(n155), 
          .S1(n152));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_3 (.A0(n194_adj_48), .B0(n63), .C0(n5224), 
          .D0(n194_adj_115), .A1(n193_adj_44), .B1(n63), .C1(n5223), 
          .D1(n193_adj_15), .CIN(n32390), .COUT(n32391), .S0(n161), 
          .S1(n158));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_7032_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_7032_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_7032_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(i[0]), .B1(n42833), .C1(n56), .D1(n55), 
          .COUT(n32390));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(107[13:38])
    defparam _add_1_7032_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_7032_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_7032_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_7032_add_4_1.INJECT1_1 = "NO";
    LUT4 div_4016_mux_5_i10_3_lut (.A(n5482), .B(n90), .C(n5460), .Z(n123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i10_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3066_i21_2_lut_rep_784 (.A(n4667), .B(n124_adj_229), 
         .Z(n42483)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i21_2_lut_rep_784.init = 16'h6666;
    LUT4 div_4016_LessThan_3066_i12_3_lut_3_lut (.A(n4667), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n12_adj_673)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2513_i36_3_lut_3_lut (.A(n3838), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n36_adj_478)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i36_3_lut_3_lut.init = 16'hd4d4;
    OB x_out_pad_55 (.I(x_out_c_55), .O(x_out[55]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    LUT4 i9299_2_lut_4_lut_4_lut (.A(n865), .B(n131_adj_234), .C(n132), 
         .D(n42787), .Z(n60_adj_162)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(B+!((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9299_2_lut_4_lut_4_lut.init = 16'hbb2b;
    LUT4 i25837_4_lut (.A(n42495), .B(n42494), .C(n42496), .D(n39264), 
         .Z(n39289)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25837_4_lut.init = 16'hfeff;
    LUT4 div_4016_LessThan_2058_i45_2_lut_rep_985 (.A(n3161), .B(n124_adj_229), 
         .Z(n42684)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i45_2_lut_rep_985.init = 16'h6666;
    OB x_out_pad_90 (.I(x_out_c_90), .O(x_out[90]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_91 (.I(x_out_c_91), .O(x_out[91]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_92 (.I(x_out_c_92), .O(x_out[92]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_93 (.I(x_out_c_93), .O(x_out[93]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_94 (.I(x_out_c_94), .O(x_out[94]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_95 (.I(x_out_c_95), .O(x_out[95]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_96 (.I(x_out_c_96), .O(x_out[96]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_97 (.I(x_out_c_97), .O(x_out[97]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_98 (.I(x_out_c_98), .O(x_out[98]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_99 (.I(x_out_c_99), .O(x_out[99]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_100 (.I(x_out_c_100), .O(x_out[100]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_101 (.I(x_out_c_101), .O(x_out[101]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_102 (.I(x_out_c_102), .O(x_out[102]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_103 (.I(x_out_c_103), .O(x_out[103]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_104 (.I(x_out_c_104), .O(x_out[104]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_105 (.I(x_out_c_105), .O(x_out[105]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_106 (.I(x_out_c_106), .O(x_out[106]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_107 (.I(x_out_c_107), .O(x_out[107]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_108 (.I(x_out_c_108), .O(x_out[108]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_109 (.I(x_out_c_109), .O(x_out[109]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_110 (.I(x_out_c_110), .O(x_out[110]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_111 (.I(x_out_c_111), .O(x_out[111]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_112 (.I(x_out_c_112), .O(x_out[112]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_113 (.I(x_out_c_113), .O(x_out[113]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_114 (.I(x_out_c_114), .O(x_out[114]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_115 (.I(x_out_c_115), .O(x_out[115]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_116 (.I(x_out_c_116), .O(x_out[116]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_117 (.I(x_out_c_117), .O(x_out[117]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_118 (.I(x_out_c_118), .O(x_out[118]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_119 (.I(x_out_c_119), .O(x_out[119]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_120 (.I(x_out_c_120), .O(x_out[120]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_121 (.I(x_out_c_121), .O(x_out[121]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_89 (.I(x_out_c_89), .O(x_out[89]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_56 (.I(x_out_c_56), .O(x_out[56]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_57 (.I(x_out_c_57), .O(x_out[57]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_58 (.I(x_out_c_58), .O(x_out[58]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_59 (.I(x_out_c_59), .O(x_out[59]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_60 (.I(x_out_c_60), .O(x_out[60]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_61 (.I(x_out_c_61), .O(x_out[61]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_62 (.I(x_out_c_62), .O(x_out[62]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_63 (.I(x_out_c_63), .O(x_out[63]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_64 (.I(x_out_c_64), .O(x_out[64]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_65 (.I(x_out_c_65), .O(x_out[65]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_66 (.I(x_out_c_66), .O(x_out[66]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_67 (.I(x_out_c_67), .O(x_out[67]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_68 (.I(x_out_c_68), .O(x_out[68]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_69 (.I(x_out_c_69), .O(x_out[69]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_70 (.I(x_out_c_70), .O(x_out[70]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_71 (.I(x_out_c_71), .O(x_out[71]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_72 (.I(x_out_c_72), .O(x_out[72]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_73 (.I(x_out_c_73), .O(x_out[73]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_74 (.I(x_out_c_74), .O(x_out[74]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_75 (.I(x_out_c_75), .O(x_out[75]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_76 (.I(x_out_c_76), .O(x_out[76]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_77 (.I(x_out_c_77), .O(x_out[77]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_78 (.I(x_out_c_78), .O(x_out[78]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_79 (.I(x_out_c_79), .O(x_out[79]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_80 (.I(x_out_c_80), .O(x_out[80]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_81 (.I(x_out_c_81), .O(x_out[81]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_82 (.I(x_out_c_82), .O(x_out[82]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_83 (.I(x_out_c_83), .O(x_out[83]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_84 (.I(x_out_c_84), .O(x_out[84]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_85 (.I(x_out_c_85), .O(x_out[85]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_86 (.I(x_out_c_86), .O(x_out[86]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_87 (.I(x_out_c_87), .O(x_out[87]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    LUT4 div_4016_LessThan_2058_i36_3_lut_3_lut (.A(n3161), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n36_adj_364)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24004_4_lut (.A(n42497), .B(n42499), .C(n42498), .D(n39248), 
         .Z(n39264)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24004_4_lut.init = 16'h1011;
    LUT4 i22867_4_lut (.A(n42652), .B(n42653), .C(n42654), .D(n38111), 
         .Z(n38127)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22867_4_lut.init = 16'h5455;
    OB x_out_pad_124 (.I(x_out_c_124), .O(x_out[124]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_88 (.I(x_out_c_88), .O(x_out[88]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    LUT4 i23988_4_lut (.A(n42500), .B(n33_adj_654), .C(n21_adj_647), .D(n39201), 
         .Z(n39248)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23988_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_2058_i43_2_lut_rep_986 (.A(n3162), .B(n125_adj_230), 
         .Z(n42685)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i43_2_lut_rep_986.init = 16'h6666;
    LUT4 i25890_2_lut_3_lut_4_lut (.A(n3162), .B(n125_adj_230), .C(n116_adj_224), 
         .D(n3153), .Z(n37965)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25890_2_lut_3_lut_4_lut.init = 16'h6ff6;
    LUT4 div_4016_i735_3_lut_4_lut (.A(n42788), .B(n132), .C(n64), .D(n30872), 
         .Z(n1230)) /* synthesis lut_function=(A ((C+(D))+!B)+!A !((C+(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i735_3_lut_4_lut.init = 16'haaa6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.A(n115_adj_223), .B(n114), .C(n36918), 
         .D(n42817), .Z(n36994)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_58.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i15_2_lut_rep_785 (.A(n4670), .B(n127_adj_231), 
         .Z(n42484)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i15_2_lut_rep_785.init = 16'h6666;
    LUT4 div_4016_LessThan_2513_i37_2_lut_rep_914 (.A(n3840), .B(n123), 
         .Z(n42613)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i37_2_lut_rep_914.init = 16'h6666;
    LUT4 i8453_4_lut_4_lut (.A(n678), .B(n132), .C(n42784), .D(n131_adj_234), 
         .Z(n62_adj_801)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A !(B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i8453_4_lut_4_lut.init = 16'ha2fb;
    PFUMX div_4016_LessThan_1862_i62 (.BLUT(n44_adj_333), .ALUT(n60_adj_341), 
          .C0(n40086), .Z(n62_adj_342));
    LUT4 i24775_4_lut_4_lut (.A(n42439), .B(n40017), .C(n53_adj_785), 
         .D(n55_adj_787), .Z(n40035)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24775_4_lut_4_lut.init = 16'h000b;
    LUT4 div_4016_LessThan_3066_i17_2_lut_rep_786 (.A(n4669), .B(n126), 
         .Z(n42485)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i17_2_lut_rep_786.init = 16'h6666;
    LUT4 i1_2_lut_rep_1110_3_lut_4_lut (.A(n115_adj_223), .B(n114), .C(n112_adj_221), 
         .D(n113_adj_222), .Z(n42809)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1110_3_lut_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2918_i59_2_lut_rep_812 (.A(n4429), .B(n107_adj_218), 
         .Z(n42511)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i59_2_lut_rep_812.init = 16'h6666;
    LUT4 i25884_2_lut_3_lut_4_lut (.A(n3840), .B(n123), .C(n111), .D(n3828), 
         .Z(n40094)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25884_2_lut_3_lut_4_lut.init = 16'h6ff6;
    LUT4 div_4016_LessThan_2513_i39_2_lut_rep_915 (.A(n3839), .B(n122_adj_228), 
         .Z(n42614)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i39_2_lut_rep_915.init = 16'h6666;
    LUT4 div_4016_LessThan_2058_i32_4_lut (.A(n132), .B(n131_adj_234), .C(n3168), 
         .D(n880), .Z(n32_adj_361)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i32_4_lut.init = 16'h0c8e;
    LUT4 i25900_3_lut_4_lut (.A(n59_adj_791), .B(n25_adj_759), .C(n61_adj_793), 
         .D(n42437), .Z(n40074)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25900_3_lut_4_lut.init = 16'hff01;
    LUT4 div_4016_LessThan_3206_i54_3_lut_4_lut (.A(n59_adj_791), .B(n25_adj_759), 
         .C(n20_adj_754), .D(n18_adj_752), .Z(n54_adj_786)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_2918_i52_3_lut_3_lut (.A(n4429), .B(n107_adj_218), 
         .C(n50_adj_633), .Z(n52_adj_634)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25174_3_lut (.A(\U[10] [21]), .B(\U[11] [21]), .C(i[0]), .Z(n40434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25174_3_lut.init = 16'hcaca;
    LUT4 i23151_2_lut_3_lut_4_lut (.A(n3839), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3838), .Z(n38411)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23151_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i22609_4_lut (.A(n42691), .B(n42698), .C(n42699), .D(n41_adj_348), 
         .Z(n37869)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22609_4_lut.init = 16'h5554;
    LUT4 i1_2_lut_rep_1118 (.A(n117), .B(n116_adj_224), .Z(n42817)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1118.init = 16'heeee;
    LUT4 div_4016_LessThan_1961_i41_2_lut (.A(n3019), .B(n127_adj_231), 
         .Z(n41_adj_348)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i41_2_lut.init = 16'h6666;
    LUT4 div_4016_mux_3_i20_3_lut (.A(n5337), .B(n14_adj_174), .C(n5325), 
         .Z(n875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i20_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.A(n117), .B(n116_adj_224), .C(n5460), 
         .D(n68_adj_194), .Z(n37054)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_59.init = 16'hfeee;
    LUT4 div_4016_LessThan_2513_i35_2_lut_rep_916 (.A(n3841), .B(n124_adj_229), 
         .Z(n42615)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i35_2_lut_rep_916.init = 16'h6666;
    LUT4 i25173_3_lut (.A(\U[8] [21]), .B(\U[9] [21]), .C(i[0]), .Z(n40433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25173_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_3_i21_3_lut (.A(n5336), .B(n13_adj_173), .C(n5325), 
         .Z(n874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i21_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_1862_i56 (.BLUT(n48_adj_335), .ALUT(n54_adj_338), 
          .C0(n37795), .Z(n56_adj_339));
    LUT4 div_4016_LessThan_1113_i64_4_lut (.A(n60_adj_258), .B(n62_adj_259), 
         .C(n42756), .D(n37480), .Z(n64_adj_260)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i64_4_lut.init = 16'hccca;
    LUT4 div_4016_LessThan_2513_i26_3_lut_3_lut (.A(n3841), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n26_adj_472)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2993_i33_2_lut (.A(n4553), .B(n119_adj_226), 
         .Z(n33_adj_654)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i33_2_lut.init = 16'h6666;
    LUT4 div_4016_mux_3_i22_3_lut (.A(n5335), .B(n12_adj_172), .C(n5325), 
         .Z(n873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i22_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_3_i23_3_lut (.A(n5334), .B(n11_adj_171), .C(n5325), 
         .Z(n872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i23_3_lut.init = 16'hcaca;
    LUT4 i25326_3_lut (.A(\U[14] [31]), .B(\U[15] [31]), .C(i[0]), .Z(n40586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25326_3_lut.init = 16'hcaca;
    LUT4 i25172_3_lut (.A(\U[6] [21]), .B(\U[7] [21]), .C(i[0]), .Z(n40432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25172_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2918_i55_2_lut_rep_813 (.A(n4431), .B(n109_adj_219), 
         .Z(n42512)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i55_2_lut_rep_813.init = 16'h6666;
    LUT4 i22220_4_lut (.A(n42757), .B(n42758), .C(n57_adj_256), .D(n37469), 
         .Z(n37480)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22220_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_2513_i29_2_lut_rep_917 (.A(n3844), .B(n127_adj_231), 
         .Z(n42616)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i29_2_lut_rep_917.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i21_2_lut (.A(n4559), .B(n125_adj_230), 
         .Z(n21_adj_647)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i21_2_lut.init = 16'h6666;
    LUT4 i24108_2_lut_3_lut_4_lut (.A(n4669), .B(n126), .C(n127_adj_231), 
         .D(n4670), .Z(n39368)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24108_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i1_2_lut_rep_1115_3_lut_4_lut (.A(n117), .B(n116_adj_224), .C(n114), 
         .D(n115_adj_223), .Z(n42814)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1115_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1119 (.A(n116_adj_224), .B(n119_adj_226), .Z(n42818)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1119.init = 16'heeee;
    LUT4 div_4016_LessThan_2513_i31_2_lut_rep_918 (.A(n3843), .B(n126), 
         .Z(n42617)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i31_2_lut_rep_918.init = 16'h6666;
    LUT4 i23124_2_lut_3_lut_4_lut (.A(n3843), .B(n126), .C(n127_adj_231), 
         .D(n3844), .Z(n38384)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23124_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i22209_4_lut (.A(n42760), .B(n42759), .C(n1754), .D(n130_adj_233), 
         .Z(n37469)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22209_4_lut.init = 16'h1001;
    LUT4 div_4016_mux_3_i24_3_lut (.A(n5333), .B(n10_adj_170), .C(n5325), 
         .Z(n685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i24_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.A(n116_adj_224), .B(n119_adj_226), 
         .C(n117), .D(n114), .Z(n37206)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_60.init = 16'hfffe;
    LUT4 div_4016_i3324_4_lut (.A(n37154), .B(n22288), .C(n42786), .D(n64_adj_315), 
         .Z(n5507)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3324_4_lut.init = 16'hc0c5;
    PFUMX div_4016_LessThan_1761_i62 (.BLUT(n46_adj_319), .ALUT(n60_adj_326), 
          .C0(n40082), .Z(n62_adj_327));
    LUT4 div_4016_mux_3_i25_3_lut (.A(n5332), .B(n9_adj_169), .C(n5325), 
         .Z(n684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i25_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_61 (.A(n30950), .B(n37146), .C(n37148), .D(n37144), 
         .Z(n37154)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_61.init = 16'hfffe;
    LUT4 i1_4_lut_adj_62 (.A(n36956), .B(n42790), .C(n36948), .D(n36946), 
         .Z(n30887)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_62.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_63 (.A(n119_adj_226), .B(n118_adj_225), 
         .C(n116_adj_224), .D(n117), .Z(n36948)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_63.init = 16'hfffe;
    LUT4 div_4016_mux_3_i26_3_lut (.A(n5331), .B(n8_adj_168), .C(n5325), 
         .Z(n683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i26_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_1761_i58 (.BLUT(n50_adj_321), .ALUT(n56_adj_324), 
          .C0(n37738), .Z(n58_adj_325));
    LUT4 div_4016_LessThan_2513_i28_3_lut_3_lut (.A(n3843), .B(n126), .C(n127_adj_231), 
         .Z(n28_adj_473)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23113_3_lut_4_lut (.A(n3846), .B(n129), .C(n130_adj_233), .D(n3847), 
         .Z(n38373)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23113_3_lut_4_lut.init = 16'h9009;
    LUT4 i1_2_lut_rep_1120 (.A(n118_adj_225), .B(n121_adj_227), .Z(n42819)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1120.init = 16'heeee;
    LUT4 div_4016_LessThan_3066_i14_3_lut_3_lut (.A(n4669), .B(n126), .C(n127_adj_231), 
         .Z(n14_adj_675)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i14_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2513_i24_3_lut_3_lut (.A(n3846), .B(n129), .C(n130_adj_233), 
         .Z(n24_adj_471)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25325_3_lut (.A(\U[12] [31]), .B(\U[13] [31]), .C(i[0]), .Z(n40585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25325_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_64 (.A(n118_adj_225), .B(n121_adj_227), 
         .C(n119_adj_226), .D(n117), .Z(n37238)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_64.init = 16'hfffe;
    LUT4 div_4016_LessThan_2513_i27_2_lut_rep_919 (.A(n3845), .B(n128_adj_232), 
         .Z(n42618)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i27_2_lut_rep_919.init = 16'h6666;
    LUT4 i23137_2_lut_3_lut_4_lut (.A(n3845), .B(n128_adj_232), .C(n124_adj_229), 
         .D(n3841), .Z(n38397)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23137_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_1113_i57_2_lut (.A(n1751), .B(n127_adj_231), 
         .Z(n57_adj_256)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1113_i57_2_lut.init = 16'h6666;
    LUT4 i25633_4_lut_4_lut (.A(n42621), .B(n38357), .C(n54_adj_464), 
         .D(n30_adj_450), .Z(n56_adj_465)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25633_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2153_i30_4_lut (.A(n132), .B(n131_adj_234), .C(n3310), 
         .D(n881), .Z(n30_adj_379)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i30_4_lut.init = 16'h0c8e;
    LUT4 i25171_3_lut (.A(\U[4] [21]), .B(\U[5] [21]), .C(i[0]), .Z(n40431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25171_3_lut.init = 16'hcaca;
    LUT4 i25739_4_lut_4_lut (.A(n42438), .B(n39985), .C(n34_adj_768), 
         .D(n10_adj_744), .Z(n36_adj_770)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25739_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_65 (.A(n118_adj_225), .B(n120), .C(n119_adj_226), 
         .D(n116_adj_224), .Z(n37172)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_65.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_66 (.A(n118_adj_225), .B(n120), .C(n119_adj_226), 
         .D(n117), .Z(n36740)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_66.init = 16'hfffe;
    LUT4 i24727_4_lut_4_lut (.A(n42438), .B(n39794), .C(n37_adj_771), 
         .D(n39_adj_773), .Z(n39987)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24727_4_lut_4_lut.init = 16'h0004;
    LUT4 div_4016_mux_5_i11_3_lut (.A(n5481), .B(n89_adj_208), .C(n5460), 
         .Z(n122_adj_228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i11_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i63_2_lut_rep_920 (.A(n3698), .B(n111), 
         .Z(n42619)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i63_2_lut_rep_920.init = 16'h6666;
    LUT4 div_4016_LessThan_2058_i39_2_lut_rep_987 (.A(n3164), .B(n127_adj_231), 
         .Z(n42686)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i39_2_lut_rep_987.init = 16'h6666;
    LUT4 div_4016_LessThan_2426_i44_3_lut_3_lut (.A(n3698), .B(n111), .C(n36_adj_454), 
         .Z(n44_adj_458)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_5_i12_3_lut (.A(n5480), .B(n88_adj_207), .C(n5460), 
         .Z(n121_adj_227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i12_3_lut.init = 16'hcaca;
    LUT4 div_4016_i613_3_lut (.A(n42787), .B(n132), .C(n36422), .Z(n1049)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i613_3_lut.init = 16'ha6a6;
    LUT4 i25324_3_lut (.A(\U[10] [31]), .B(\U[11] [31]), .C(i[0]), .Z(n40584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25324_3_lut.init = 16'hcaca;
    LUT4 i25323_3_lut (.A(\U[8] [31]), .B(\U[9] [31]), .C(i[0]), .Z(n40583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25323_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_67 (.A(n120), .B(n121_adj_227), .C(n118_adj_225), 
         .D(n119_adj_226), .Z(n36918)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_67.init = 16'hfffe;
    LUT4 div_4016_LessThan_2426_i59_2_lut_rep_921 (.A(n3700), .B(n113_adj_222), 
         .Z(n42620)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i59_2_lut_rep_921.init = 16'h6666;
    LUT4 div_4016_LessThan_2426_i52_3_lut_3_lut (.A(n3700), .B(n113_adj_222), 
         .C(n114), .Z(n52_adj_463)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2426_i61_2_lut_rep_922 (.A(n3699), .B(n112_adj_221), 
         .Z(n42621)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i61_2_lut_rep_922.init = 16'h6666;
    LUT4 div_4016_LessThan_2918_i57_2_lut_rep_814 (.A(n4430), .B(n108), 
         .Z(n42513)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i57_2_lut_rep_814.init = 16'h6666;
    LUT4 i25170_3_lut (.A(\U[2] [21]), .B(\U[3] [21]), .C(i[0]), .Z(n40430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25170_3_lut.init = 16'hcaca;
    LUT4 i25169_3_lut (.A(\U[0] [21]), .B(\U[1] [21]), .C(i[0]), .Z(n40429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25169_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_1658_i60 (.BLUT(n52_adj_309), .ALUT(n58_adj_312), 
          .C0(n37686), .Z(n60_adj_313));
    LUT4 i1_2_lut_rep_1121 (.A(n122_adj_228), .B(n125_adj_230), .Z(n42820)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1121.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_68 (.A(n122_adj_228), .B(n125_adj_230), .C(n123), 
         .D(n121_adj_227), .Z(n36492)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_68.init = 16'hfffe;
    LUT4 div_4016_LessThan_3206_i12_3_lut (.A(n125_adj_230), .B(n116_adj_224), 
         .C(n33_adj_767), .Z(n12_adj_746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i12_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2058_i41_2_lut_rep_988 (.A(n3163), .B(n126), 
         .Z(n42687)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i41_2_lut_rep_988.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_69 (.A(n123), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n120), .Z(n36946)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_69.init = 16'hfffe;
    LUT4 div_4016_LessThan_3066_i11_2_lut_rep_787 (.A(n4672), .B(n129), 
         .Z(n42486)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i11_2_lut_rep_787.init = 16'h6666;
    LUT4 i25835_4_lut (.A(n42495), .B(n42494), .C(n42496), .D(n39273), 
         .Z(n39291)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25835_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_3137_i11_2_lut (.A(n4777), .B(n128_adj_232), 
         .Z(n11_adj_707)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i11_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_70 (.A(n124_adj_229), .B(n125_adj_230), 
         .C(n122_adj_228), .D(n123), .Z(n36916)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_70.init = 16'hfffe;
    LUT4 div_4016_mux_3_i4_3_lut (.A(n5353), .B(n30_adj_190), .C(n5325), 
         .Z(n891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 mux_4010_i4_4_lut (.A(n154), .B(n36650), .C(n15805), .D(i[1]), 
         .Z(n5353)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i4_4_lut.init = 16'hca0a;
    LUT4 i22137_2_lut_rep_1122 (.A(n124_adj_229), .B(n127_adj_231), .Z(n42821)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22137_2_lut_rep_1122.init = 16'heeee;
    LUT4 div_4016_LessThan_2426_i54_3_lut_3_lut (.A(n3699), .B(n112_adj_221), 
         .C(n52_adj_463), .Z(n54_adj_464)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i54_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_1658_i62 (.BLUT(n48_adj_307), .ALUT(n50_adj_308), 
          .C0(n40080), .Z(n62_adj_314));
    LUT4 i22145_2_lut_3_lut_4_lut (.A(n124_adj_229), .B(n127_adj_231), .C(n125_adj_230), 
         .D(n122_adj_228), .Z(n37370)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22145_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2246_i28_4_lut (.A(n132), .B(n131_adj_234), .C(n3449), 
         .D(n882), .Z(n28_adj_400)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i28_4_lut.init = 16'h0c8e;
    LUT4 i1_2_lut_adj_71 (.A(i[0]), .B(\y[3] [3]), .Z(n36650)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_71.init = 16'h8888;
    LUT4 div_4016_mux_5_i30_3_lut (.A(n5462), .B(n70_adj_195), .C(n5460), 
         .Z(n103_adj_215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i30_3_lut.init = 16'hcaca;
    LUT4 i22640_2_lut_3_lut_4_lut (.A(n3163), .B(n126), .C(n127_adj_231), 
         .D(n3164), .Z(n37900)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22640_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_3206_i23_4_lut (.A(n4771), .B(n121_adj_227), 
         .C(n22261), .D(n4783), .Z(n23_adj_757)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i23_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2918_i50_3_lut_3_lut (.A(n4430), .B(n108), .C(n109_adj_219), 
         .Z(n50_adj_633)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2058_i38_3_lut_3_lut (.A(n3163), .B(n126), .C(n127_adj_231), 
         .Z(n38_adj_365)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_5_i18_3_lut (.A(n5474), .B(n82_adj_203), .C(n5460), 
         .Z(n115_adj_223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i18_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i57_2_lut_rep_923 (.A(n3701), .B(n114), 
         .Z(n42622)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i57_2_lut_rep_923.init = 16'h6666;
    LUT4 div_4016_LessThan_2058_i35_2_lut_rep_989 (.A(n3166), .B(n129), 
         .Z(n42688)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i35_2_lut_rep_989.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i41_4_lut_rep_739 (.A(n4762), .B(n112_adj_221), 
         .C(n22252), .D(n4783), .Z(n42438)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i41_4_lut_rep_739.init = 16'h663c;
    LUT4 i23097_2_lut_3_lut_4_lut (.A(n3701), .B(n114), .C(n113_adj_222), 
         .D(n3700), .Z(n38357)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23097_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_i488_4_lut (.A(n678), .B(n42781), .C(n42775), .D(n131_adj_234), 
         .Z(n864)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i488_4_lut.init = 16'ha6a9;
    LUT4 i1_3_lut_4_lut_adj_72 (.A(n126), .B(n127_adj_231), .C(n128_adj_232), 
         .D(n129), .Z(n36802)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_72.init = 16'hfffe;
    LUT4 div_4016_LessThan_2426_i55_2_lut_rep_924 (.A(n3702), .B(n115_adj_223), 
         .Z(n42623)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i55_2_lut_rep_924.init = 16'h6666;
    LUT4 div_4016_LessThan_2058_i34_3_lut_3_lut (.A(n3166), .B(n129), .C(n130_adj_233), 
         .Z(n34_adj_363)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25597_4_lut_4_lut (.A(n42690), .B(n37876), .C(n56_adj_356), 
         .D(n34), .Z(n58_adj_357)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25597_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_3066_i10_3_lut_3_lut (.A(n4672), .B(n129), .C(n130_adj_233), 
         .Z(n10_adj_672)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_adj_73 (.A(n126), .B(n127_adj_231), .C(n125_adj_230), 
         .D(n124_adj_229), .Z(n36872)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_73.init = 16'hfffe;
    LUT4 i25915_4_lut_4_lut (.A(n42690), .B(n37869), .C(n42692), .D(n42689), 
         .Z(n37885)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25915_4_lut_4_lut.init = 16'hff04;
    LUT4 div_4016_LessThan_2426_i50_3_lut_3_lut (.A(n3702), .B(n115_adj_223), 
         .C(n32_adj_451), .Z(n50_adj_462)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25919_4_lut_4_lut (.A(n42690), .B(n37864), .C(n42692), .D(n42689), 
         .Z(n37879)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25919_4_lut_4_lut.init = 16'hfffb;
    LUT4 div_4016_i793_1_lut_rep_1123 (.A(n129), .Z(n42822)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i793_1_lut_rep_1123.init = 16'h5555;
    LUT4 i25704_4_lut_4_lut (.A(n42487), .B(n39328), .C(n28_adj_651), 
         .D(n12_adj_642), .Z(n56_adj_666)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25704_4_lut_4_lut.init = 16'hf4b0;
    LUT4 n1047_bdd_4_lut_26064_4_lut (.A(n129), .B(n42769), .C(n42825), 
         .D(n1047), .Z(n42432)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam n1047_bdd_4_lut_26064_4_lut.init = 16'hfd54;
    LUT4 div_4016_i426_1_lut_rep_1124 (.A(n131_adj_234), .Z(n42823)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i426_1_lut_rep_1124.init = 16'h5555;
    LUT4 i23086_3_lut_4_lut (.A(n3702), .B(n115_adj_223), .C(n35_adj_453), 
         .D(n42625), .Z(n38346)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23086_3_lut_4_lut.init = 16'h0009;
    LUT4 i23906_4_lut (.A(n42513), .B(n42512), .C(n42514), .D(n39150), 
         .Z(n39166)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23906_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_2426_i51_2_lut_rep_925 (.A(n3704), .B(n117), 
         .Z(n42624)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i51_2_lut_rep_925.init = 16'h6666;
    PFUMX div_4016_LessThan_1553_i62 (.BLUT(n54_adj_296), .ALUT(n60_adj_299), 
          .C0(n37637), .Z(n62_adj_300));
    LUT4 div_4016_LessThan_2426_i46_3_lut_3_lut (.A(n3704), .B(n117), .C(n34_adj_452), 
         .Z(n46_adj_459)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3137_i29_2_lut (.A(n4768), .B(n119_adj_226), 
         .Z(n29_adj_719)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i29_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i26_4_lut (.A(n132), .B(n131_adj_234), .C(n3585), 
         .D(n883), .Z(n26_adj_422)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i26_4_lut.init = 16'h0c8e;
    LUT4 i25810_3_lut_4_lut (.A(n3704), .B(n117), .C(n47_adj_460), .D(n42626), 
         .Z(n38330)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25810_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_2426_i53_2_lut_rep_926 (.A(n3703), .B(n116_adj_224), 
         .Z(n42625)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i53_2_lut_rep_926.init = 16'h6666;
    LUT4 i23908_2_lut_3_lut_4_lut (.A(n4430), .B(n108), .C(n109_adj_219), 
         .D(n4431), .Z(n39168)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23908_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2426_i32_3_lut_3_lut (.A(n3703), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n32_adj_451)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2993_i61_2_lut_rep_788 (.A(n4539), .B(n105), 
         .Z(n42487)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i61_2_lut_rep_788.init = 16'h6666;
    LUT4 div_4016_i673_1_lut_rep_1125 (.A(n130_adj_233), .Z(n42824)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i673_1_lut_rep_1125.init = 16'h5555;
    LUT4 i25631_4_lut_4_lut (.A(n42627), .B(n38301), .C(n40_adj_456), 
         .D(n26_adj_447), .Z(n42_adj_457)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25631_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i23149_4_lut (.A(n42612), .B(n42614), .C(n42613), .D(n38397), 
         .Z(n38409)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23149_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_1961_i63_2_lut_rep_990 (.A(n3008), .B(n116_adj_224), 
         .Z(n42689)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i63_2_lut_rep_990.init = 16'h6666;
    LUT4 i25887_4_lut_4_lut (.A(n42627), .B(n38294), .C(n42628), .D(n42619), 
         .Z(n40090)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25887_4_lut_4_lut.init = 16'hff04;
    LUT4 n864_bdd_4_lut_4_lut (.A(n130_adj_233), .B(n42774), .C(n23957), 
         .D(n864), .Z(n42430)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam n864_bdd_4_lut_4_lut.init = 16'hfd54;
    LUT4 div_4016_LessThan_2993_i28_3_lut_3_lut (.A(n4539), .B(n105), .C(n106_adj_217), 
         .Z(n28_adj_651)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i9576_2_lut_rep_1070_3_lut_4_lut_4_lut_4_lut (.A(n130_adj_233), .B(n42783), 
         .C(n42773), .D(n131_adj_234), .Z(n42769)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9576_2_lut_rep_1070_3_lut_4_lut_4_lut_4_lut.init = 16'h5054;
    LUT4 div_4016_LessThan_2426_i49_2_lut_rep_927 (.A(n3705), .B(n118_adj_225), 
         .Z(n42626)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i49_2_lut_rep_927.init = 16'h6666;
    LUT4 div_4016_LessThan_2426_i34_3_lut_3_lut (.A(n3705), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n34_adj_452)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25161_3_lut (.A(\U[14] [20]), .B(\U[15] [20]), .C(i[0]), .Z(n40421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25161_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i45_2_lut_rep_928 (.A(n3707), .B(n120), 
         .Z(n42627)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i45_2_lut_rep_928.init = 16'h6666;
    LUT4 i25686_4_lut_4_lut (.A(n42517), .B(n39126), .C(n42_adj_629), 
         .D(n18_adj_614), .Z(n44_adj_630)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25686_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2993_i63_2_lut_rep_789 (.A(n4538), .B(n104_adj_216), 
         .Z(n42488)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i63_2_lut_rep_789.init = 16'h6666;
    LUT4 div_4016_mux_5_i22_3_lut (.A(n5470), .B(n78), .C(n5460), .Z(n111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i22_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1961_i60_3_lut_3_lut (.A(n3008), .B(n116_adj_224), 
         .C(n42_adj_349), .Z(n60_adj_358)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23904_4_lut (.A(n42513), .B(n42512), .C(n42514), .D(n39143), 
         .Z(n39164)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23904_4_lut.init = 16'h0100;
    PFUMX div_4016_LessThan_1553_i52 (.BLUT(n42), .ALUT(n50_adj_294), .C0(n37610), 
          .Z(n52_adj_295));
    LUT4 i23883_4_lut (.A(n42515), .B(n42524), .C(n42523), .D(n39063), 
         .Z(n39143)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23883_4_lut.init = 16'h5455;
    LUT4 i15194_4_lut_4_lut_rep_1126 (.A(n130_adj_233), .B(n42773), .C(n42779), 
         .D(n1048), .Z(n42825)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i15194_4_lut_4_lut_rep_1126.init = 16'hfd00;
    LUT4 i25160_3_lut (.A(\U[12] [20]), .B(\U[13] [20]), .C(i[0]), .Z(n40420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25160_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i51_4_lut_rep_740 (.A(n4757), .B(n107_adj_218), 
         .C(n22247), .D(n4783), .Z(n42439)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i51_4_lut_rep_740.init = 16'h663c;
    LUT4 div_4016_LessThan_2993_i60_3_lut_3_lut (.A(n4538), .B(n104_adj_216), 
         .C(n58_adj_667), .Z(n60_adj_668)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1961_i61_2_lut_rep_991 (.A(n3009), .B(n117), 
         .Z(n42690)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i61_2_lut_rep_991.init = 16'h6666;
    LUT4 i9578_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n130_adj_233), .B(n42773), 
         .C(n42779), .D(n1048), .Z(n60)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9578_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hfd54;
    LUT4 i23803_4_lut (.A(n29_adj_621), .B(n42525), .C(n42526), .D(n17_adj_613), 
         .Z(n39063)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23803_4_lut.init = 16'h5554;
    LUT4 i25741_4_lut_4_lut (.A(n42439), .B(n40021), .C(n44_adj_777), 
         .D(n8_adj_742), .Z(n46_adj_779)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25741_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i23869_4_lut_4_lut (.A(n42517), .B(n39104), .C(n42519), .D(n42516), 
         .Z(n39129)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23869_4_lut_4_lut.init = 16'h0004;
    LUT4 div_4016_LessThan_2426_i40_3_lut_3_lut (.A(n3707), .B(n120), .C(n38_adj_455), 
         .Z(n40_adj_456)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i612_4_lut (.A(n865), .B(n42782), .C(n36422), .D(n131_adj_234), 
         .Z(n1048)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i612_4_lut.init = 16'ha6a9;
    LUT4 div_4016_LessThan_2426_i24_4_lut (.A(n132), .B(n131_adj_234), .C(n3718), 
         .D(n884), .Z(n24_adj_445)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i24_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2918_i29_2_lut (.A(n4444), .B(n122_adj_228), 
         .Z(n29_adj_621)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i29_2_lut.init = 16'h6666;
    LUT4 i15195_3_lut_rep_1074_4_lut (.A(n131_adj_234), .B(n132), .C(n42788), 
         .D(n1049), .Z(n42773)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i15195_3_lut_rep_1074_4_lut.init = 16'hf700;
    LUT4 div_4016_LessThan_2918_i17_2_lut (.A(n4450), .B(n128_adj_232), 
         .Z(n17_adj_613)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i17_2_lut.init = 16'h6666;
    LUT4 i25702_4_lut_4_lut (.A(n42489), .B(n39326), .C(n50_adj_663), 
         .D(n14_adj_643), .Z(n52_adj_664)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25702_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2426_i43_2_lut_rep_929 (.A(n3708), .B(n121_adj_227), 
         .Z(n42628)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i43_2_lut_rep_929.init = 16'h6666;
    LUT4 i25159_3_lut (.A(\U[10] [20]), .B(\U[11] [20]), .C(i[0]), .Z(n40419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25159_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_1446_i62 (.BLUT(n56_adj_285), .ALUT(n60_adj_287), 
          .C0(n37588), .Z(n62_adj_288));
    LUT4 div_4016_LessThan_2426_i38_3_lut_3_lut (.A(n3708), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n38_adj_455)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i53_2_lut_rep_815 (.A(n4432), .B(n110_adj_220), 
         .Z(n42514)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i53_2_lut_rep_815.init = 16'h6666;
    LUT4 i15219_3_lut_rep_1075_4_lut (.A(n131_adj_234), .B(n132), .C(n42787), 
         .D(n865), .Z(n42774)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i15219_3_lut_rep_1075_4_lut.init = 16'hf700;
    LUT4 div_4016_i427_1_lut_rep_1128 (.A(n132), .Z(n42827)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i427_1_lut_rep_1128.init = 16'h5555;
    LUT4 i25158_3_lut (.A(\U[8] [20]), .B(\U[9] [20]), .C(i[0]), .Z(n40418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25158_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i39_2_lut_rep_930 (.A(n3710), .B(n123), 
         .Z(n42629)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i39_2_lut_rep_930.init = 16'h6666;
    LUT4 i25157_3_lut (.A(\U[6] [20]), .B(\U[7] [20]), .C(i[0]), .Z(n40417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25157_3_lut.init = 16'hcaca;
    LUT4 i9569_2_lut_rep_1080_3_lut_3_lut_3_lut (.A(n132), .B(n42788), .C(n131_adj_234), 
         .Z(n42779)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9569_2_lut_rep_1080_3_lut_3_lut_3_lut.init = 16'h0d0d;
    LUT4 i25322_3_lut (.A(\U[6] [31]), .B(\U[7] [31]), .C(i[0]), .Z(n40582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25322_3_lut.init = 16'hcaca;
    LUT4 i8445_2_lut_rep_1082_4_lut_4_lut (.A(n132), .B(n5325), .C(n4_adj_164), 
         .D(n5327), .Z(n42781)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i8445_2_lut_rep_1082_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i24080_4_lut_4_lut_4_lut (.A(n42489), .B(n39328), .C(n39311), 
         .D(n42487), .Z(n39340)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24080_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i24071_4_lut_4_lut (.A(n42489), .B(n39306), .C(n42490), .D(n42491), 
         .Z(n39331)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24071_4_lut_4_lut.init = 16'h0004;
    LUT4 i25789_4_lut (.A(n42605), .B(n42604), .C(n42606), .D(n38456), 
         .Z(n38474)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25789_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2426_i36_3_lut_3_lut (.A(n3710), .B(n123), .C(n28_adj_448), 
         .Z(n36_adj_454)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25706_4_lut_4_lut (.A(n42489), .B(n39324), .C(n52_adj_664), 
         .D(n30_adj_652), .Z(n54_adj_665)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25706_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2993_i57_2_lut_rep_790 (.A(n4541), .B(n107_adj_218), 
         .Z(n42489)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i57_2_lut_rep_790.init = 16'h6666;
    LUT4 div_4016_LessThan_2426_i41_2_lut_rep_931 (.A(n3709), .B(n122_adj_228), 
         .Z(n42630)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i41_2_lut_rep_931.init = 16'h6666;
    LUT4 div_4016_i3318_4_lut (.A(n37250), .B(n22282), .C(n42786), .D(n64_adj_252), 
         .Z(n5501)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3318_4_lut.init = 16'hc0c5;
    LUT4 div_4016_i734_4_lut (.A(n1049), .B(n42783), .C(n1078), .D(n131_adj_234), 
         .Z(n1229)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i734_4_lut.init = 16'ha6a9;
    LUT4 i23041_2_lut_3_lut_4_lut (.A(n3709), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3708), .Z(n38301)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23041_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2513_i22_4_lut (.A(n132), .B(n131_adj_234), .C(n3848), 
         .D(n885), .Z(n22_adj_470)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i22_4_lut.init = 16'h0c8e;
    LUT4 i25863_4_lut (.A(n42517), .B(n42516), .C(n42519), .D(n39106), 
         .Z(n39131)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25863_4_lut.init = 16'hfeff;
    LUT4 i25156_3_lut (.A(\U[4] [20]), .B(\U[5] [20]), .C(i[0]), .Z(n40416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25156_3_lut.init = 16'hcaca;
    LUT4 i23846_4_lut (.A(n42518), .B(n42521), .C(n42520), .D(n39090), 
         .Z(n39106)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23846_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_2918_i32_3_lut_3_lut (.A(n4432), .B(n110_adj_220), 
         .C(n24_adj_618), .Z(n32_adj_623)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23830_4_lut (.A(n42522), .B(n35_adj_625), .C(n23_adj_617), .D(n39043), 
         .Z(n39090)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23830_4_lut.init = 16'h1011;
    LUT4 i1_4_lut_adj_74 (.A(n37242), .B(n35919), .C(n37244), .D(n37240), 
         .Z(n37250)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_74.init = 16'hfffe;
    LUT4 div_4016_mux_5_i23_3_lut (.A(n5469), .B(n77_adj_200), .C(n5460), 
         .Z(n110_adj_220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i23_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i37_2_lut_rep_932 (.A(n3711), .B(n124_adj_229), 
         .Z(n42631)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i37_2_lut_rep_932.init = 16'h6666;
    LUT4 i9291_2_lut_rep_1083_4_lut_4_lut (.A(n132), .B(n5325), .C(n5_adj_165), 
         .D(n5328), .Z(n42782)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9291_2_lut_rep_1083_4_lut_4_lut.init = 16'hf7d5;
    LUT4 div_4016_LessThan_2426_i28_3_lut_3_lut (.A(n3711), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n28_adj_448)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_3_i27_3_lut (.A(n5330), .B(n7_adj_167), .C(n5325), 
         .Z(n682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i27_3_lut.init = 16'hcaca;
    LUT4 i9297_2_lut_3_lut_3_lut_3_lut (.A(n132), .B(n42787), .C(n131_adj_234), 
         .Z(n23957)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9297_2_lut_3_lut_3_lut_3_lut.init = 16'h0d0d;
    LUT4 i25155_3_lut (.A(\U[2] [20]), .B(\U[3] [20]), .C(i[0]), .Z(n40415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25155_3_lut.init = 16'hcaca;
    LUT4 i9563_2_lut_rep_1084_4_lut_4_lut (.A(n132), .B(n5325), .C(n6_adj_166), 
         .D(n5329), .Z(n42783)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i9563_2_lut_rep_1084_4_lut_4_lut.init = 16'hf7d5;
    PFUMX div_4016_LessThan_1446_i54 (.BLUT(n44), .ALUT(n52_adj_283), .C0(n37568), 
          .Z(n54_adj_284));
    LUT4 i25321_3_lut (.A(\U[4] [31]), .B(\U[5] [31]), .C(i[0]), .Z(n40581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25321_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1961_i56_3_lut_3_lut (.A(n3009), .B(n117), .C(n44_adj_350), 
         .Z(n56_adj_356)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_4_lut_adj_75 (.A(n37238), .B(n37256), .C(n122_adj_228), .D(n124_adj_229), 
         .Z(n37244)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_75.init = 16'hfffe;
    LUT4 i25154_3_lut (.A(\U[0] [20]), .B(\U[1] [20]), .C(i[0]), .Z(n40414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25154_3_lut.init = 16'hcaca;
    LUT4 n1049_bdd_4_lut (.A(n1049), .B(n132), .C(n131_adj_234), .D(n42788), 
         .Z(n42835)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(B (C+!(D))+!B (C))) */ ;
    defparam n1049_bdd_4_lut.init = 16'haf2b;
    LUT4 i25146_3_lut (.A(\U[14] [19]), .B(\U[15] [19]), .C(i[0]), .Z(n40406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25146_3_lut.init = 16'hcaca;
    LUT4 mux_6984_i30_3_lut_4_lut (.A(n42829), .B(n42828), .C(n74), .D(n32356), 
         .Z(n25248)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_2918_i35_2_lut (.A(n4441), .B(n119_adj_226), 
         .Z(n35_adj_625)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i35_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2918_i23_2_lut (.A(n4447), .B(n125_adj_230), 
         .Z(n23_adj_617)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i23_2_lut.init = 16'h6666;
    LUT4 mux_6984_i32_3_lut_4_lut (.A(n42829), .B(n42828), .C(n68), .D(n32354), 
         .Z(n25244)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_76 (.A(n120), .B(n123), .Z(n37256)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_76.init = 16'heeee;
    LUT4 i25320_3_lut (.A(\U[2] [31]), .B(\U[3] [31]), .C(i[0]), .Z(n40580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25320_3_lut.init = 16'hcaca;
    LUT4 div_4016_i3175_3_lut_rep_741 (.A(n4751), .B(n22241), .C(n4783), 
         .Z(n42440)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3175_3_lut_rep_741.init = 16'hacac;
    LUT4 div_4016_LessThan_2993_i50_3_lut_3_lut (.A(n4541), .B(n107_adj_218), 
         .C(n48_adj_662), .Z(n50_adj_663)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i50_3_lut_3_lut.init = 16'hd4d4;
    PFUMX div_4016_LessThan_1337_i62 (.BLUT(n58_adj_275), .ALUT(n60_adj_276), 
          .C0(n37548), .Z(n62_adj_277));
    LUT4 div_4016_LessThan_2918_i51_2_lut_rep_816 (.A(n4433), .B(n111), 
         .Z(n42515)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i51_2_lut_rep_816.init = 16'h6666;
    LUT4 i25872_4_lut (.A(n42550), .B(n42552), .C(n42551), .D(n38866), 
         .Z(n40110)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25872_4_lut.init = 16'hfffe;
    LUT4 i25594_4_lut_4_lut (.A(n42693), .B(n37854), .C(n50_adj_353), 
         .D(n36_adj_344), .Z(n52_adj_354)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25594_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25145_3_lut (.A(\U[12] [19]), .B(\U[13] [19]), .C(i[0]), .Z(n40405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25145_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i33_2_lut_rep_933 (.A(n3713), .B(n126), 
         .Z(n42632)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i33_2_lut_rep_933.init = 16'h6666;
    LUT4 mux_6984_i31_3_lut_4_lut (.A(n42829), .B(n42828), .C(n71), .D(n32355), 
         .Z(n25246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_998_i64_4_lut (.A(n56_adj_248), .B(n62_adj_251), 
         .C(n42761), .D(n37455), .Z(n64_adj_252)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i64_4_lut.init = 16'hcacc;
    LUT4 mux_6984_i28_3_lut_4_lut (.A(n42829), .B(n42828), .C(n80), .D(n32358), 
         .Z(n25252)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22195_4_lut (.A(n42762), .B(n59), .C(n42763), .D(n37446), 
         .Z(n37455)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22195_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_2426_i30_3_lut_3_lut (.A(n3713), .B(n126), .C(n127_adj_231), 
         .Z(n30_adj_450)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_6984_i29_3_lut_4_lut (.A(n42829), .B(n42828), .C(n77), .D(n32357), 
         .Z(n25250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i26_3_lut_4_lut (.A(n42829), .B(n42828), .C(n86), .D(n32360), 
         .Z(n25256)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22604_4_lut_4_lut (.A(n42693), .B(n37843), .C(n42694), .D(n42691), 
         .Z(n37864)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22604_4_lut_4_lut.init = 16'h00fb;
    LUT4 div_4016_LessThan_2426_i31_2_lut_rep_934 (.A(n3714), .B(n127_adj_231), 
         .Z(n42633)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i31_2_lut_rep_934.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i53_2_lut_rep_791 (.A(n4543), .B(n109_adj_219), 
         .Z(n42490)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i53_2_lut_rep_791.init = 16'h6666;
    LUT4 div_4016_LessThan_1961_i57_2_lut_rep_992 (.A(n3011), .B(n119_adj_226), 
         .Z(n42691)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i57_2_lut_rep_992.init = 16'h6666;
    LUT4 i23014_2_lut_3_lut_4_lut (.A(n3714), .B(n127_adj_231), .C(n126), 
         .D(n3713), .Z(n38274)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23014_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 mux_6984_i27_3_lut_4_lut (.A(n42829), .B(n42828), .C(n83), .D(n32359), 
         .Z(n25254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i25319_3_lut (.A(\U[0] [31]), .B(\U[1] [31]), .C(i[0]), .Z(n40579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25319_3_lut.init = 16'hcaca;
    LUT4 i25144_3_lut (.A(\U[10] [19]), .B(\U[11] [19]), .C(i[0]), .Z(n40404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25144_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i27_2_lut_rep_935 (.A(n3716), .B(n129), 
         .Z(n42634)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i27_2_lut_rep_935.init = 16'h6666;
    LUT4 i25143_3_lut (.A(\U[8] [19]), .B(\U[9] [19]), .C(i[0]), .Z(n40403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25143_3_lut.init = 16'hcaca;
    LUT4 mux_6984_i24_3_lut_4_lut (.A(n42829), .B(n42828), .C(n92), .D(n32362), 
         .Z(n25260)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_2918_i24_3_lut_3_lut (.A(n4433), .B(n111), .C(n123), 
         .Z(n24_adj_618)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_6984_i25_3_lut_4_lut (.A(n42829), .B(n42828), .C(n89), .D(n32361), 
         .Z(n25258)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_3206_i63_2_lut_rep_738_4_lut (.A(n4751), .B(n22241), 
         .C(n4783), .D(n42796), .Z(n42437)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i63_2_lut_rep_738_4_lut.init = 16'h53ac;
    LUT4 div_4016_LessThan_2918_i47_2_lut_rep_817 (.A(n4435), .B(n113_adj_222), 
         .Z(n42516)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i47_2_lut_rep_817.init = 16'h6666;
    LUT4 i25730_4_lut_4_lut (.A(n42443), .B(n39698), .C(n52_adj_731), 
         .D(n8_adj_705), .Z(n54_adj_732)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25730_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25853_4_lut (.A(n42510), .B(n42524), .C(n42523), .D(n29_adj_621), 
         .Z(n39186)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25853_4_lut.init = 16'haaab;
    LUT4 mux_6984_i22_3_lut_4_lut (.A(n42829), .B(n42828), .C(n98), .D(n32364), 
         .Z(n25264)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_1961_i59_2_lut_rep_993 (.A(n3010), .B(n118_adj_225), 
         .Z(n42692)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i59_2_lut_rep_993.init = 16'h6666;
    LUT4 mux_6984_i23_3_lut_4_lut (.A(n42829), .B(n42828), .C(n95), .D(n32363), 
         .Z(n25262)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_998_i59_2_lut (.A(n1579), .B(n127_adj_231), .Z(n59)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_998_i59_2_lut.init = 16'h6666;
    LUT4 i25142_3_lut (.A(\U[6] [19]), .B(\U[7] [19]), .C(i[0]), .Z(n40402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25142_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2426_i26_3_lut_3_lut (.A(n3716), .B(n129), .C(n130_adj_233), 
         .Z(n26_adj_447)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2426_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i40_3_lut_3_lut (.A(n4435), .B(n113_adj_222), 
         .C(n114), .Z(n40_adj_628)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25311_3_lut (.A(\U[14] [30]), .B(\U[15] [30]), .C(i[0]), .Z(n40571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25311_3_lut.init = 16'hcaca;
    LUT4 i25625_4_lut_4_lut (.A(n42635), .B(n38250), .C(n56_adj_440), 
         .D(n32_adj_426), .Z(n58_adj_441)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25625_4_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6984_i20_3_lut_4_lut (.A(n42829), .B(n42828), .C(n104), .D(n32366), 
         .Z(n25268)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i21_3_lut_4_lut (.A(n42829), .B(n42828), .C(n101), .D(n32365), 
         .Z(n25266)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_2598_i20_4_lut (.A(n132), .B(n131_adj_234), .C(n3975), 
         .D(n886), .Z(n20_adj_494)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i20_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2337_i63_2_lut_rep_936 (.A(n3566), .B(n112_adj_221), 
         .Z(n42635)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i63_2_lut_rep_936.init = 16'h6666;
    LUT4 mux_6984_i18_3_lut_4_lut (.A(n42829), .B(n42828), .C(n110), .D(n32368), 
         .Z(n25272)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i25310_3_lut (.A(\U[12] [30]), .B(\U[13] [30]), .C(i[0]), .Z(n40570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25310_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_1337_i56 (.BLUT(n46), .ALUT(n54_adj_273), .C0(n37533), 
          .Z(n56_adj_274));
    LUT4 div_4016_LessThan_2337_i56_3_lut_3_lut (.A(n3566), .B(n112_adj_221), 
         .C(n54_adj_439), .Z(n56_adj_440)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_6984_i19_3_lut_4_lut (.A(n42829), .B(n42828), .C(n107), .D(n32367), 
         .Z(n25270)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i16_3_lut_4_lut (.A(n42829), .B(n42828), .C(n116), .D(n32370), 
         .Z(n25276)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i17_3_lut_4_lut (.A(n42829), .B(n42828), .C(n113), .D(n32369), 
         .Z(n25274)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_1961_i44_3_lut_3_lut (.A(n3010), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n44_adj_350)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22616_2_lut_3_lut_4_lut (.A(n3010), .B(n118_adj_225), .C(n119_adj_226), 
         .D(n3011), .Z(n37876)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22616_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i25141_3_lut (.A(\U[4] [19]), .B(\U[5] [19]), .C(i[0]), .Z(n40401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25141_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2337_i61_2_lut_rep_937 (.A(n3567), .B(n113_adj_222), 
         .Z(n42636)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i61_2_lut_rep_937.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i55_2_lut_rep_792 (.A(n4542), .B(n108), 
         .Z(n42491)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i55_2_lut_rep_792.init = 16'h6666;
    LUT4 i24066_2_lut_3_lut_4_lut (.A(n4542), .B(n108), .C(n109_adj_219), 
         .D(n4543), .Z(n39326)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24066_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 mux_6984_i14_3_lut_4_lut (.A(n42829), .B(n42828), .C(n122), .D(n32372), 
         .Z(n25280)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_77 (.A(n42791), .B(n42801), .C(n106_adj_217), .D(n108), 
         .Z(n35919)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_77.init = 16'hfffe;
    LUT4 div_4016_mux_3_i10_3_lut (.A(n5347), .B(n24_adj_184), .C(n5325), 
         .Z(n885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i10_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2337_i54_3_lut_3_lut (.A(n3567), .B(n113_adj_222), 
         .C(n114), .Z(n54_adj_439)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2337_i57_2_lut_rep_938 (.A(n3569), .B(n115_adj_223), 
         .Z(n42637)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i57_2_lut_rep_938.init = 16'h6666;
    PFUMX div_4016_LessThan_1226_i60 (.BLUT(n50_adj_261), .ALUT(n52_adj_262), 
          .C0(n37513), .Z(n60_adj_267));
    LUT4 div_4016_LessThan_2918_i49_2_lut_rep_818 (.A(n4434), .B(n112_adj_221), 
         .Z(n42517)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i49_2_lut_rep_818.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i52_3_lut_3_lut (.A(n3569), .B(n115_adj_223), 
         .C(n34_adj_427), .Z(n52_adj_438)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1961_i55_2_lut_rep_994 (.A(n3012), .B(n120), 
         .Z(n42693)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i55_2_lut_rep_994.init = 16'h6666;
    LUT4 mux_6984_i15_3_lut_4_lut (.A(n42829), .B(n42828), .C(n119), .D(n32371), 
         .Z(n25278)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_1961_i50_3_lut_3_lut (.A(n3012), .B(n120), .C(n48_adj_352), 
         .Z(n50_adj_353)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25768_4_lut_4_lut (.A(n42443), .B(n39696), .C(n42441), .D(n42442), 
         .Z(n39716)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25768_4_lut_4_lut.init = 16'hfff4;
    LUT4 mux_6984_i12_3_lut_4_lut (.A(n42829), .B(n42828), .C(n128), .D(n32374), 
         .Z(n25284)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i13_3_lut_4_lut (.A(n42829), .B(n42828), .C(n125), .D(n32373), 
         .Z(n25282)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_2993_i48_3_lut_3_lut (.A(n4542), .B(n108), .C(n109_adj_219), 
         .Z(n48_adj_662)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22979_3_lut_4_lut (.A(n3569), .B(n115_adj_223), .C(n37_adj_429), 
         .D(n42640), .Z(n38239)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22979_3_lut_4_lut.init = 16'h0009;
    LUT4 mux_6984_i10_3_lut_4_lut (.A(n42829), .B(n42828), .C(n134), .D(n32376), 
         .Z(n25288)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i25697_4_lut_4_lut (.A(n42495), .B(n39284), .C(n40_adj_658), 
         .D(n16_adj_644), .Z(n42_adj_659)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25697_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25861_4_lut (.A(n42517), .B(n42516), .C(n42519), .D(n39115), 
         .Z(n39133)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25861_4_lut.init = 16'hfffe;
    LUT4 i25140_3_lut (.A(\U[2] [19]), .B(\U[3] [19]), .C(i[0]), .Z(n40400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25140_3_lut.init = 16'hcaca;
    LUT4 i25848_2_lut (.A(done_N_1931), .B(rst_c), .Z(clk_c_enable_541)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam i25848_2_lut.init = 16'h2222;
    LUT4 i25925_4_lut (.A(n42693), .B(n42694), .C(n42695), .D(n37845), 
         .Z(n37859)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25925_4_lut.init = 16'hfffe;
    LUT4 mux_6984_i11_3_lut_4_lut (.A(n42829), .B(n42828), .C(n131), .D(n32375), 
         .Z(n25286)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_1961_i39_2_lut (.A(n3020), .B(n128_adj_232), 
         .Z(n39_adj_346)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i39_2_lut.init = 16'h6666;
    LUT4 i25309_3_lut (.A(\U[10] [30]), .B(\U[11] [30]), .C(i[0]), .Z(n40569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25309_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2337_i59_2_lut_rep_939 (.A(n3568), .B(n114), 
         .Z(n42638)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i59_2_lut_rep_939.init = 16'h6666;
    LUT4 i25139_3_lut (.A(\U[0] [19]), .B(\U[1] [19]), .C(i[0]), .Z(n40399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25139_3_lut.init = 16'hcaca;
    LUT4 i25308_3_lut (.A(\U[8] [30]), .B(\U[9] [30]), .C(i[0]), .Z(n40568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25308_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1961_i53_2_lut_rep_995 (.A(n3013), .B(n121_adj_227), 
         .Z(n42694)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i53_2_lut_rep_995.init = 16'h6666;
    LUT4 div_4016_i3323_4_lut (.A(n64_adj_301), .B(n22287), .C(n42786), 
         .D(n42789), .Z(n5506)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3323_4_lut.init = 16'hc0c5;
    LUT4 mux_6984_i8_3_lut_4_lut (.A(n42829), .B(n42828), .C(n140), .D(n32378), 
         .Z(n25292)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22990_2_lut_3_lut_4_lut (.A(n3568), .B(n114), .C(n113_adj_222), 
         .D(n3567), .Z(n38250)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22990_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2337_i53_2_lut_rep_940 (.A(n3571), .B(n117), 
         .Z(n42639)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i53_2_lut_rep_940.init = 16'h6666;
    LUT4 div_4016_LessThan_2918_i42_3_lut_3_lut (.A(n4434), .B(n112_adj_221), 
         .C(n40_adj_628), .Z(n42_adj_629)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_6984_i9_3_lut_4_lut (.A(n42829), .B(n42828), .C(n137), .D(n32377), 
         .Z(n25290)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i6_3_lut_4_lut (.A(n42829), .B(n42828), .C(n146), .D(n32380), 
         .Z(n25296)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_LessThan_3137_i61_2_lut_rep_742 (.A(n4752), .B(n103_adj_215), 
         .Z(n42441)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i61_2_lut_rep_742.init = 16'h6666;
    LUT4 div_4016_LessThan_3137_i22_3_lut_3_lut (.A(n4752), .B(n103_adj_215), 
         .C(n120), .Z(n22_adj_715)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i43_2_lut_rep_819 (.A(n4437), .B(n115_adj_223), 
         .Z(n42518)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i43_2_lut_rep_819.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i48_3_lut_3_lut (.A(n3571), .B(n117), .C(n36_adj_428), 
         .Z(n48_adj_435)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25828_3_lut_4_lut (.A(n3571), .B(n117), .C(n49_adj_436), .D(n42641), 
         .Z(n38223)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25828_3_lut_4_lut.init = 16'hfff6;
    LUT4 mux_6984_i7_3_lut_4_lut (.A(n42829), .B(n42828), .C(n143), .D(n32379), 
         .Z(n25294)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i25131_3_lut (.A(\U[14] [18]), .B(\U[15] [18]), .C(i[0]), .Z(n40391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25131_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2918_i38_3_lut_3_lut (.A(n4437), .B(n115_adj_223), 
         .C(n20_adj_615), .Z(n38_adj_627)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2681_i18_4_lut (.A(n132), .B(n131_adj_234), .C(n4099), 
         .D(n887), .Z(n18_adj_521)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i18_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2337_i55_2_lut_rep_941 (.A(n3570), .B(n116_adj_224), 
         .Z(n42640)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i55_2_lut_rep_941.init = 16'h6666;
    LUT4 mux_6984_i4_3_lut_4_lut (.A(n42829), .B(n42828), .C(n152), .D(n32382), 
         .Z(n25300)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_6984_i5_3_lut_4_lut (.A(n42829), .B(n42828), .C(n149), .D(n32381), 
         .Z(n25298)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24036_4_lut_4_lut (.A(n42495), .B(n39269), .C(n42494), .D(n42493), 
         .Z(n39296)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24036_4_lut_4_lut.init = 16'h00fb;
    LUT4 div_4016_LessThan_1961_i48_3_lut_3_lut (.A(n3013), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n48_adj_352)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_6984_i2_3_lut_4_lut (.A(n42829), .B(n42828), .C(n158), .D(n32384), 
         .Z(n25304)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i2_3_lut_4_lut.init = 16'hf1e0;
    PFUMX div_4016_LessThan_1226_i58 (.BLUT(n48), .ALUT(n56_adj_265), .C0(n37505), 
          .Z(n58_adj_266));
    LUT4 i25130_3_lut (.A(\U[12] [18]), .B(\U[13] [18]), .C(i[0]), .Z(n40390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25130_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2337_i34_3_lut_3_lut (.A(n3570), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n34_adj_427)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_6984_i3_3_lut_4_lut (.A(n42829), .B(n42828), .C(n155), .D(n32383), 
         .Z(n25302)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i25129_3_lut (.A(\U[10] [18]), .B(\U[11] [18]), .C(i[0]), .Z(n40389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25129_3_lut.init = 16'hcaca;
    LUT4 i25128_3_lut (.A(\U[8] [18]), .B(\U[9] [18]), .C(i[0]), .Z(n40388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25128_3_lut.init = 16'hcaca;
    LUT4 mux_6984_i1_3_lut_4_lut (.A(n42829), .B(n42828), .C(n161), .D(n32385), 
         .Z(n25306)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam mux_6984_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_4016_mux_3_i5_3_lut (.A(n5352), .B(n29_adj_189), .C(n5325), 
         .Z(n890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 i28_2_lut_rep_1129 (.A(n55), .B(n56), .Z(n42828)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i28_2_lut_rep_1129.init = 16'heeee;
    LUT4 i25621_4_lut_4_lut (.A(n42643), .B(n38194), .C(n42_adj_432), 
         .D(n28_adj_423), .Z(n44_adj_433)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25621_4_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_4010_i5_4_lut (.A(n151), .B(n36648), .C(n15805), .D(i[1]), 
         .Z(n5352)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i5_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_78 (.A(i[0]), .B(\y[3] [4]), .Z(n36648)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_78.init = 16'h8888;
    LUT4 div_4016_LessThan_2337_i51_2_lut_rep_942 (.A(n3572), .B(n118_adj_225), 
         .Z(n42641)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i51_2_lut_rep_942.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i36_3_lut_3_lut (.A(n3572), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n36_adj_428)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2337_i45_2_lut_rep_943 (.A(n3575), .B(n121_adj_227), 
         .Z(n42642)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i45_2_lut_rep_943.init = 16'h6666;
    LUT4 i16244_3_lut_4_lut (.A(n55), .B(n56), .C(n42833), .D(n42831), 
         .Z(n15805)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(101[15:21])
    defparam i16244_3_lut_4_lut.init = 16'hfeee;
    LUT4 i22151_3_lut (.A(done_N_1934), .B(n16519), .Z(n37411)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22151_3_lut.init = 16'heeee;
    LUT4 i12827_2_lut (.A(done_N_1929), .B(start_c), .Z(n27528)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12827_2_lut.init = 16'h2222;
    LUT4 div_4016_LessThan_1961_i51_2_lut_rep_996 (.A(n3014), .B(n122_adj_228), 
         .Z(n42695)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i51_2_lut_rep_996.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i40_3_lut_3_lut (.A(n3575), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n40_adj_431)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22594_2_lut_3_lut_4_lut (.A(n3014), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3013), .Z(n37854)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22594_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2993_i51_2_lut_rep_793 (.A(n4544), .B(n110_adj_220), 
         .Z(n42492)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i51_2_lut_rep_793.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i47_2_lut_rep_944 (.A(n3574), .B(n120), 
         .Z(n42643)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i47_2_lut_rep_944.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i30_3_lut_3_lut (.A(n4544), .B(n110_adj_220), 
         .C(n22_adj_648), .Z(n30_adj_652)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23855_3_lut_4_lut (.A(n4437), .B(n115_adj_223), .C(n23_adj_617), 
         .D(n42521), .Z(n39115)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23855_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_1961_i49_2_lut_rep_997 (.A(n3015), .B(n123), 
         .Z(n42696)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i49_2_lut_rep_997.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_79 (.A(i[0]), .B(n42833), .C(n56), .D(n55), 
         .Z(n63)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_2_lut_3_lut_4_lut_adj_79.init = 16'hfffd;
    LUT4 div_4016_LessThan_1961_i46_3_lut_3_lut (.A(n3015), .B(n123), .C(n38_adj_345), 
         .Z(n46_adj_351)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_3_lut_4_lut_adj_80 (.A(i[0]), .B(n42833), .C(n42830), .D(n37334), 
         .Z(n31021)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_3_lut_4_lut_adj_80.init = 16'h2000;
    LUT4 i25127_3_lut (.A(\U[6] [18]), .B(\U[7] [18]), .C(i[0]), .Z(n40387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25127_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2993_i49_2_lut_rep_794 (.A(n4545), .B(n111), 
         .Z(n42493)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i49_2_lut_rep_794.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i42_3_lut_3_lut (.A(n3574), .B(n120), .C(n40_adj_431), 
         .Z(n42_adj_432)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23755_4_lut (.A(n42533), .B(n42532), .C(n42535), .D(n38999), 
         .Z(n39015)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23755_4_lut.init = 16'h1011;
    LUT4 i1_3_lut_4_lut_adj_81 (.A(i[0]), .B(n42832), .C(n42830), .D(n37334), 
         .Z(n31084)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_3_lut_4_lut_adj_81.init = 16'h2000;
    LUT4 div_4016_LessThan_2337_i41_2_lut_rep_945 (.A(n3577), .B(n123), 
         .Z(n42644)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i41_2_lut_rep_945.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i38_3_lut_3_lut (.A(n3577), .B(n123), .C(n30_adj_424), 
         .Z(n38_adj_430)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25126_3_lut (.A(\U[4] [18]), .B(\U[5] [18]), .C(i[0]), .Z(n40386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25126_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_82 (.A(i[0]), .B(n42833), .C(n42830), .D(n37334), 
         .Z(n30987)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_3_lut_4_lut_adj_82.init = 16'h1000;
    LUT4 i23744_4_lut (.A(n42532), .B(n42535), .C(n42534), .D(n38924), 
         .Z(n39004)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23744_4_lut.init = 16'h0001;
    LUT4 i23664_4_lut (.A(n42544), .B(n42543), .C(n31_adj_590), .D(n38910), 
         .Z(n38924)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23664_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_2841_i31_2_lut (.A(n4329), .B(n122_adj_228), 
         .Z(n31_adj_590)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i31_2_lut.init = 16'h6666;
    LUT4 i22925_3_lut_4_lut (.A(n3577), .B(n123), .C(n31_adj_425), .D(n42646), 
         .Z(n38185)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22925_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2841_i19_2_lut (.A(n4335), .B(n128_adj_232), 
         .Z(n19_adj_582)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i19_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i43_2_lut_rep_946 (.A(n3576), .B(n122_adj_228), 
         .Z(n42645)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i43_2_lut_rep_946.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i22_3_lut_3_lut (.A(n4545), .B(n111), .C(n123), 
         .Z(n22_adj_648)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22934_2_lut_3_lut_4_lut (.A(n3576), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3575), .Z(n38194)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22934_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2337_i39_2_lut_rep_947 (.A(n3578), .B(n124_adj_229), 
         .Z(n42646)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i39_2_lut_rep_947.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i30_3_lut_3_lut (.A(n3578), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n30_adj_424)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2337_i33_2_lut_rep_948 (.A(n3581), .B(n127_adj_231), 
         .Z(n42647)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i33_2_lut_rep_948.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i45_2_lut_rep_795 (.A(n4547), .B(n113_adj_222), 
         .Z(n42494)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i45_2_lut_rep_795.init = 16'h6666;
    LUT4 div_4016_LessThan_2762_i16_4_lut (.A(n132), .B(n131_adj_234), .C(n4220), 
         .D(n888), .Z(n16_adj_550)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i16_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2337_i35_2_lut_rep_949 (.A(n3580), .B(n126), 
         .Z(n42648)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i35_2_lut_rep_949.init = 16'h6666;
    LUT4 i1_2_lut_rep_1133 (.A(i[2]), .B(i[1]), .Z(n42832)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_2_lut_rep_1133.init = 16'hbbbb;
    LUT4 i22907_2_lut_3_lut_4_lut (.A(n3580), .B(n126), .C(n127_adj_231), 
         .D(n3581), .Z(n38167)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22907_2_lut_3_lut_4_lut.init = 16'h9009;
    PFUMX div_4016_LessThan_1113_i60 (.BLUT(n50), .ALUT(n58_adj_257), .C0(n37482), 
          .Z(n60_adj_258));
    LUT4 i25889_4_lut (.A(n42701), .B(n42703), .C(n42702), .D(n37768), 
         .Z(n40086)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25889_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1132_3_lut (.A(i[2]), .B(i[1]), .C(i[0]), .Z(n42831)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_2_lut_rep_1132_3_lut.init = 16'hfbfb;
    LUT4 div_4016_LessThan_2993_i38_3_lut_3_lut (.A(n4547), .B(n113_adj_222), 
         .C(n114), .Z(n38_adj_657)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22585_3_lut_4_lut (.A(n3015), .B(n123), .C(n39_adj_346), .D(n42697), 
         .Z(n37845)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22585_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2993_i47_2_lut_rep_796 (.A(n4546), .B(n112_adj_221), 
         .Z(n42495)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i47_2_lut_rep_796.init = 16'h6666;
    LUT4 i25804_4_lut (.A(n42621), .B(n42620), .C(n42622), .D(n38337), 
         .Z(n38362)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25804_4_lut.init = 16'hfeff;
    LUT4 div_4016_LessThan_2993_i40_3_lut_3_lut (.A(n4546), .B(n112_adj_221), 
         .C(n38_adj_657), .Z(n40_adj_658)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23077_4_lut (.A(n42623), .B(n42625), .C(n42624), .D(n38321), 
         .Z(n38337)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23077_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_rep_1134 (.A(i[1]), .B(i[2]), .Z(n42833)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_2_lut_rep_1134.init = 16'heeee;
    LUT4 i25908_4_lut (.A(n42537), .B(n42536), .C(n42539), .D(n38955), 
         .Z(n38980)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25908_4_lut.init = 16'hfeff;
    LUT4 div_4016_LessThan_3137_i63_2_lut_rep_743 (.A(n4751), .B(n102), 
         .Z(n42442)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i63_2_lut_rep_743.init = 16'h6666;
    LUT4 i25307_3_lut (.A(\U[6] [30]), .B(\U[7] [30]), .C(i[0]), .Z(n40567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25307_3_lut.init = 16'hcaca;
    LUT4 i23695_4_lut (.A(n42538), .B(n42541), .C(n42540), .D(n38939), 
         .Z(n38955)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23695_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_1862_i43_2_lut (.A(n2871), .B(n127_adj_231), 
         .Z(n43_adj_332)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i43_2_lut.init = 16'h6666;
    LUT4 i25125_3_lut (.A(\U[2] [18]), .B(\U[3] [18]), .C(i[0]), .Z(n40385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25125_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i58_3_lut_3_lut (.A(n4751), .B(n102), .C(n56_adj_733), 
         .Z(n58_adj_734)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2337_i32_3_lut_3_lut (.A(n3580), .B(n126), .C(n127_adj_231), 
         .Z(n32_adj_426)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i45_2_lut_rep_820 (.A(n4436), .B(n114), 
         .Z(n42519)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i45_2_lut_rep_820.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i29_2_lut_rep_950 (.A(n3583), .B(n129), 
         .Z(n42649)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i29_2_lut_rep_950.init = 16'h6666;
    LUT4 div_4016_LessThan_1961_i47_2_lut_rep_998 (.A(n3016), .B(n124_adj_229), 
         .Z(n42697)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i47_2_lut_rep_998.init = 16'h6666;
    LUT4 i23866_2_lut_3_lut_4_lut (.A(n4436), .B(n114), .C(n113_adj_222), 
         .D(n4435), .Z(n39126)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23866_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i23061_4_lut (.A(n42626), .B(n47_adj_460), .C(n35_adj_453), .D(n38274), 
         .Z(n38321)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23061_4_lut.init = 16'h1011;
    LUT4 i23679_4_lut (.A(n42542), .B(n37_adj_594), .C(n25_adj_586), .D(n38892), 
         .Z(n38939)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23679_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_rep_1130_3_lut (.A(i[1]), .B(i[2]), .C(i[0]), .Z(n42829)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(118[13:17])
    defparam i1_2_lut_rep_1130_3_lut.init = 16'hfefe;
    LUT4 i12632_1_lut_rep_1135 (.A(rst_c), .Z(clk_c_enable_831)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i12632_1_lut_rep_1135.init = 16'h5555;
    LUT4 div_4016_LessThan_1961_i38_3_lut_3_lut (.A(n3016), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n38_adj_345)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25124_3_lut (.A(\U[0] [18]), .B(\U[1] [18]), .C(i[0]), .Z(n40384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25124_3_lut.init = 16'hcaca;
    PFUMX div_4016_LessThan_998_i62 (.BLUT(n52), .ALUT(n60_adj_250), .C0(n37462), 
          .Z(n62_adj_251));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_c), .B(i[0]), .C(n42833), 
         .D(done_N_1932), .Z(clk_c_enable_812)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 div_4016_LessThan_1961_i45_2_lut_rep_999 (.A(n3017), .B(n125_adj_230), 
         .Z(n42698)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i45_2_lut_rep_999.init = 16'h6666;
    LUT4 div_4016_LessThan_2337_i28_3_lut_3_lut (.A(n3583), .B(n129), .C(n130_adj_233), 
         .Z(n28_adj_423)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2337_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_83 (.A(rst_c), .B(i[0]), .C(n42833), 
         .D(done_N_1932), .Z(clk_c_enable_832)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_83.init = 16'h0100;
    LUT4 i1_2_lut_rep_1131_2_lut (.A(rst_c), .B(done_N_1932), .Z(n42830)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i1_2_lut_rep_1131_2_lut.init = 16'h4444;
    LUT4 i25617_4_lut_4_lut (.A(n42650), .B(n38136), .C(n56_adj_417), 
         .D(n34_adj_404), .Z(n58_adj_418)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25617_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_84 (.A(rst_c), .B(done_N_1932), 
         .C(n42832), .D(i[0]), .Z(clk_c_enable_780)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_84.init = 16'h0004;
    LUT4 div_4016_LessThan_2841_i37_2_lut (.A(n4326), .B(n119_adj_226), 
         .Z(n37_adj_594)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i37_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2246_i63_2_lut_rep_951 (.A(n3431), .B(n113_adj_222), 
         .Z(n42650)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i63_2_lut_rep_951.init = 16'h6666;
    LUT4 div_4016_LessThan_2246_i56_3_lut_3_lut (.A(n3431), .B(n113_adj_222), 
         .C(n114), .Z(n56_adj_417)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_85 (.A(rst_c), .B(i[0]), .C(n42832), 
         .D(done_N_1932), .Z(clk_c_enable_829)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_85.init = 16'h0400;
    LUT4 div_4016_LessThan_2841_i25_2_lut (.A(n4332), .B(n125_adj_230), 
         .Z(n25_adj_586)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i25_2_lut.init = 16'h6666;
    LUT4 i1_3_lut_4_lut_4_lut (.A(rst_c), .B(n42831), .C(n37334), .D(done_N_1932), 
         .Z(n31054)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 div_4016_LessThan_2246_i59_2_lut_rep_952 (.A(n3433), .B(n115_adj_223), 
         .Z(n42651)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i59_2_lut_rep_952.init = 16'h6666;
    LUT4 i12825_2_lut_2_lut (.A(rst_c), .B(done_N_1934), .Z(clk_c_enable_677)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i12825_2_lut_2_lut.init = 16'h4444;
    LUT4 i25802_4_lut (.A(n42621), .B(n42620), .C(n42622), .D(n38346), 
         .Z(n38364)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25802_4_lut.init = 16'hfffe;
    LUT4 i12977_2_lut_2_lut (.A(rst_c), .B(done_N_1931), .Z(clk_c_enable_708)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(6[24:27])
    defparam i12977_2_lut_2_lut.init = 16'h4444;
    LUT4 i22851_4_lut (.A(n51_adj_414), .B(n42659), .C(n42661), .D(n35_adj_405), 
         .Z(n38111)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22851_4_lut.init = 16'h5554;
    LUT4 i25841_4_lut (.A(n42650), .B(n38136), .C(n42651), .D(n38134), 
         .Z(n38150)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25841_4_lut.init = 16'hbfbb;
    LUT4 div_4016_mux_3_i13_3_lut (.A(n5344), .B(n21_adj_181), .C(n5325), 
         .Z(n882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i13_3_lut.init = 16'hcaca;
    LUT4 i25306_3_lut (.A(\U[4] [30]), .B(\U[5] [30]), .C(i[0]), .Z(n40566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25306_3_lut.init = 16'hcaca;
    LUT4 i25850_4_lut (.A(n42656), .B(n42655), .C(n42657), .D(n38087), 
         .Z(n38101)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25850_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2993_i43_2_lut_rep_797 (.A(n4548), .B(n114), 
         .Z(n42496)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i43_2_lut_rep_797.init = 16'h6666;
    LUT4 div_4016_LessThan_2841_i14_4_lut (.A(n132), .B(n131_adj_234), .C(n4338), 
         .D(n889), .Z(n14_adj_579)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i14_4_lut.init = 16'h0c8e;
    LUT4 i1_2_lut_adj_86 (.A(n130_adj_233), .B(n30965), .Z(n30962)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_86.init = 16'heeee;
    LUT4 div_4016_LessThan_2246_i54_3_lut_3_lut (.A(n3433), .B(n115_adj_223), 
         .C(n36_adj_406), .Z(n54_adj_416)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2246_i57_2_lut_rep_953 (.A(n3434), .B(n116_adj_224), 
         .Z(n42652)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i57_2_lut_rep_953.init = 16'h6666;
    LUT4 i1_4_lut_adj_87 (.A(n36994), .B(n30917), .C(n36916), .D(n36802), 
         .Z(n30965)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_87.init = 16'hfffe;
    LUT4 div_4016_LessThan_393_i62_4_lut (.A(n132), .B(n131_adj_234), .C(n678), 
         .D(n42784), .Z(n62_adj_798)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_393_i62_4_lut.init = 16'h0c8e;
    LUT4 i24024_2_lut_3_lut_4_lut (.A(n4548), .B(n114), .C(n113_adj_222), 
         .D(n4547), .Z(n39284)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24024_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2246_i36_3_lut_3_lut (.A(n3434), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n36_adj_406)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i39_2_lut_rep_821 (.A(n4439), .B(n117), 
         .Z(n42520)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i39_2_lut_rep_821.init = 16'h6666;
    LUT4 div_4016_LessThan_266_i64_4_lut (.A(n132), .B(n131_adj_234), .C(n35974), 
         .D(n42785), .Z(n64_adj_799)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_266_i64_4_lut.init = 16'hc0e8;
    LUT4 div_4016_LessThan_1961_i42_3_lut_3_lut (.A(n3017), .B(n125_adj_230), 
         .C(n40_adj_347), .Z(n42_adj_349)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25116_3_lut (.A(\U[14] [17]), .B(\U[15] [17]), .C(i[0]), .Z(n40376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25116_3_lut.init = 16'hcaca;
    LUT4 i25906_4_lut (.A(n42537), .B(n42536), .C(n42539), .D(n38964), 
         .Z(n38982)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25906_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_1961_i43_2_lut_rep_1000 (.A(n3018), .B(n126), 
         .Z(n42699)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i43_2_lut_rep_1000.init = 16'h6666;
    LUT4 i23034_4_lut (.A(n42630), .B(n42629), .C(n42631), .D(n29_adj_449), 
         .Z(n38294)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23034_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_1961_i40_3_lut_3_lut (.A(n3018), .B(n126), .C(n127_adj_231), 
         .Z(n40_adj_347)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2993_i41_2_lut_rep_798 (.A(n4549), .B(n115_adj_223), 
         .Z(n42497)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i41_2_lut_rep_798.init = 16'h6666;
    LUT4 div_4016_LessThan_3137_i59_2_lut_rep_744 (.A(n4753), .B(n104_adj_216), 
         .Z(n42443)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i59_2_lut_rep_744.init = 16'h6666;
    LUT4 div_4016_LessThan_1961_i37_2_lut_rep_1001 (.A(n3021), .B(n129), 
         .Z(n42700)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i37_2_lut_rep_1001.init = 16'h6666;
    LUT4 div_4016_LessThan_3137_i52_3_lut_3_lut (.A(n4753), .B(n104_adj_216), 
         .C(n24_adj_716), .Z(n52_adj_731)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_rep_1_4_lut (.A(n36636), .B(n42780), .C(n30911), .D(n37374), 
         .Z(n35974)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i1_rep_1_4_lut.init = 16'h333b;
    LUT4 i4100_2_lut (.A(start_c), .B(done_N_1929), .Z(n10098)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i4100_2_lut.init = 16'h8888;
    PFUMX div_4016_LessThan_881_i64 (.BLUT(n58_adj_243), .ALUT(n62_adj_245), 
          .C0(n37440), .Z(n64_adj_246));
    LUT4 i1_4_lut_adj_88 (.A(n36624), .B(n42819), .C(n42818), .D(n37256), 
         .Z(n36636)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i1_4_lut_adj_88.init = 16'h0002;
    LUT4 div_4016_LessThan_2246_i55_2_lut_rep_954 (.A(n3435), .B(n117), 
         .Z(n42653)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i55_2_lut_rep_954.init = 16'h6666;
    LUT4 i25115_3_lut (.A(\U[12] [17]), .B(\U[13] [17]), .C(i[0]), .Z(n40375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25115_3_lut.init = 16'hcaca;
    LUT4 i22149_4_lut (.A(n37370), .B(n37364), .C(n128_adj_232), .D(n131_adj_234), 
         .Z(n37374)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22149_4_lut.init = 16'hfffe;
    LUT4 i12832_3_lut (.A(done_N_1932), .B(done_N_1931), .C(n16519), .Z(n27533)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i12832_3_lut.init = 16'hcece;
    LUT4 i1_3_lut (.A(n130_adj_233), .B(n117), .C(n132), .Z(n36624)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i1_3_lut.init = 16'h1010;
    LUT4 div_4016_LessThan_2246_i50_3_lut_3_lut (.A(n3435), .B(n117), .C(n38_adj_407), 
         .Z(n50_adj_413)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i34_3_lut_3_lut (.A(n4439), .B(n117), .C(n22_adj_616), 
         .Z(n34_adj_624)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25933_4_lut (.A(n42704), .B(n42705), .C(n42706), .D(n37781), 
         .Z(n37795)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25933_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_1862_i41_2_lut (.A(n2872), .B(n128_adj_232), 
         .Z(n41)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i41_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_1961_i36_3_lut_3_lut (.A(n3021), .B(n129), .C(n130_adj_233), 
         .Z(n36_adj_344)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1961_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25591_4_lut_4_lut (.A(n42701), .B(n37812), .C(n58_adj_340), 
         .D(n36), .Z(n60_adj_341)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25591_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_1761_i61_2_lut (.A(n2712), .B(n119_adj_226), 
         .Z(n37742)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i61_2_lut.init = 16'h9999;
    LUT4 div_4016_LessThan_1862_i63_2_lut_rep_1002 (.A(n2861), .B(n117), 
         .Z(n42701)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i63_2_lut_rep_1002.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i25_4_lut (.A(n4770), .B(n120), .C(n22260), 
         .D(n4783), .Z(n25_adj_759)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i25_4_lut.init = 16'h663c;
    LUT4 div_4016_mux_5_i3_3_lut (.A(n5489), .B(n97_adj_213), .C(n5460), 
         .Z(n130_adj_233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i3_3_lut.init = 16'hcaca;
    LUT4 i25892_4_lut (.A(n42711), .B(n37742), .C(n42717), .D(n37706), 
         .Z(n40082)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25892_4_lut.init = 16'hbfbb;
    LUT4 i25114_3_lut (.A(\U[10] [17]), .B(\U[11] [17]), .C(i[0]), .Z(n40374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25114_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1862_i58_3_lut_3_lut (.A(n2861), .B(n117), .C(n46_adj_334), 
         .Z(n58_adj_340)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25305_3_lut (.A(\U[2] [30]), .B(\U[3] [30]), .C(i[0]), .Z(n40565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25305_3_lut.init = 16'hcaca;
    LUT4 i25113_3_lut (.A(\U[8] [17]), .B(\U[9] [17]), .C(i[0]), .Z(n40373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25113_3_lut.init = 16'hcaca;
    LUT4 i25304_3_lut (.A(\U[0] [30]), .B(\U[1] [30]), .C(i[0]), .Z(n40564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25304_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i57_2_lut_rep_745 (.A(n4754), .B(n105), 
         .Z(n42444)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i57_2_lut_rep_745.init = 16'h6666;
    LUT4 i25870_3_lut_4_lut (.A(n4439), .B(n117), .C(n35_adj_625), .D(n42522), 
         .Z(n39099)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25870_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_mux_5_i4_3_lut (.A(n5488), .B(n96), .C(n5460), .Z(n129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i4_3_lut.init = 16'hcaca;
    LUT4 i25112_3_lut (.A(\U[6] [17]), .B(\U[7] [17]), .C(i[0]), .Z(n40372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25112_3_lut.init = 16'hcaca;
    LUT4 i25588_4_lut_4_lut (.A(n42704), .B(n37790), .C(n52_adj_337), 
         .D(n38_adj_329), .Z(n54_adj_338)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25588_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2918_i41_2_lut_rep_822 (.A(n4438), .B(n116_adj_224), 
         .Z(n42521)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i41_2_lut_rep_822.init = 16'h6666;
    LUT4 i25111_3_lut (.A(\U[4] [17]), .B(\U[5] [17]), .C(i[0]), .Z(n40371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25111_3_lut.init = 16'hcaca;
    LUT4 i22533_4_lut_4_lut (.A(n42704), .B(n37774), .C(n42706), .D(n42705), 
         .Z(n37793)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22533_4_lut_4_lut.init = 16'h0004;
    LUT4 div_4016_LessThan_1862_i59_2_lut_rep_1003 (.A(n2863), .B(n119_adj_226), 
         .Z(n42702)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i59_2_lut_rep_1003.init = 16'h6666;
    LUT4 i22139_2_lut (.A(n126), .B(n129), .Z(n37364)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22139_2_lut.init = 16'heeee;
    LUT4 div_4016_LessThan_3137_i24_3_lut_3_lut (.A(n4754), .B(n105), .C(n106_adj_217), 
         .Z(n24_adj_716)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25949_4_lut (.A(n42712), .B(n42713), .C(n42714), .D(n37724), 
         .Z(n37738)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25949_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2918_i20_3_lut_3_lut (.A(n4438), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n20_adj_615)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_mux_3_i6_3_lut (.A(n5351), .B(n28_adj_188), .C(n5325), 
         .Z(n889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i6_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1862_i61_2_lut_rep_1004 (.A(n2862), .B(n118_adj_225), 
         .Z(n42703)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i61_2_lut_rep_1004.init = 16'h6666;
    LUT4 i25846_3_lut_4_lut (.A(n3435), .B(n117), .C(n51_adj_414), .D(n42654), 
         .Z(n38125)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25846_3_lut_4_lut.init = 16'hfff6;
    PFUMX div_4016_LessThan_762_i64 (.BLUT(n60_adj_239), .ALUT(n62_adj_240), 
          .C0(n37427), .Z(n64_adj_241));
    LUT4 mux_4010_i6_4_lut (.A(n148), .B(n36652), .C(n15805), .D(i[1]), 
         .Z(n5351)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i6_4_lut.init = 16'hca0a;
    LUT4 i22552_2_lut_3_lut_4_lut (.A(n2862), .B(n118_adj_225), .C(n119_adj_226), 
         .D(n2863), .Z(n37812)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22552_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_mux_3_i11_3_lut (.A(n5346), .B(n23_adj_183), .C(n5325), 
         .Z(n884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 i25613_4_lut_4_lut (.A(n42656), .B(n38096), .C(n44_adj_410), 
         .D(n30_adj_401), .Z(n46_adj_411)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25613_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_adj_89 (.A(i[0]), .B(\y[3] [5]), .Z(n36652)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_89.init = 16'h8888;
    LUT4 i25110_3_lut (.A(\U[2] [17]), .B(\U[3] [17]), .C(i[0]), .Z(n40370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25110_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_90 (.A(n36760), .B(n36752), .C(n42799), .D(n36734), 
         .Z(n35916)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_90.init = 16'hfffe;
    PFUMX div_4016_LessThan_641_i64 (.BLUT(n58), .ALUT(n62), .C0(n37417), 
          .Z(n64));
    LUT4 i25109_3_lut (.A(\U[0] [17]), .B(\U[1] [17]), .C(i[0]), .Z(n40369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25109_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i43_2_lut (.A(n2721), .B(n128_adj_232), 
         .Z(n43)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i43_2_lut.init = 16'h6666;
    LUT4 i25101_3_lut (.A(\U[14] [16]), .B(\U[15] [16]), .C(i[0]), .Z(n40361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25101_3_lut.init = 16'hcaca;
    LUT4 i25726_4_lut_4_lut (.A(n42445), .B(n39671), .C(n46_adj_728), 
         .D(n10_adj_706), .Z(n48_adj_729)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25726_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2918_i37_2_lut_rep_823 (.A(n4440), .B(n118_adj_225), 
         .Z(n42522)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i37_2_lut_rep_823.init = 16'h6666;
    LUT4 i1_4_lut_adj_91 (.A(n36756), .B(n36744), .C(n36720), .D(n42796), 
         .Z(n36760)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_91.init = 16'hfffe;
    LUT4 div_4016_LessThan_1862_i46_3_lut_3_lut (.A(n2862), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n46_adj_334)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_4_lut_adj_92 (.A(n36740), .B(n121_adj_227), .C(n103_adj_215), 
         .D(n122_adj_228), .Z(n36752)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_92.init = 16'hfffe;
    LUT4 div_4016_LessThan_1862_i57_2_lut_rep_1005 (.A(n2864), .B(n120), 
         .Z(n42704)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i57_2_lut_rep_1005.init = 16'h6666;
    LUT4 div_4016_LessThan_2918_i22_3_lut_3_lut (.A(n4440), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n22_adj_616)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25100_3_lut (.A(\U[12] [16]), .B(\U[13] [16]), .C(i[0]), .Z(n40360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25100_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2993_i36_3_lut_3_lut (.A(n4549), .B(n115_adj_223), 
         .C(n18_adj_645), .Z(n36_adj_656)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2246_i53_2_lut_rep_955 (.A(n3436), .B(n118_adj_225), 
         .Z(n42654)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i53_2_lut_rep_955.init = 16'h6666;
    LUT4 i1_3_lut_adj_93 (.A(n104_adj_216), .B(n123), .C(n125_adj_230), 
         .Z(n36734)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_93.init = 16'hfefe;
    PFUMX div_4016_LessThan_518_i64 (.BLUT(n60_adj_795), .ALUT(n62_adj_796), 
          .C0(n40078), .Z(n64_adj_797));
    LUT4 div_4016_LessThan_1862_i52_3_lut_3_lut (.A(n2864), .B(n120), .C(n50_adj_336), 
         .Z(n52_adj_337)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3137_i53_2_lut_rep_746 (.A(n4756), .B(n107_adj_218), 
         .Z(n42445)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i53_2_lut_rep_746.init = 16'h6666;
    LUT4 div_4016_LessThan_2246_i38_3_lut_3_lut (.A(n3436), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n38_adj_407)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25753_4_lut (.A(n42722), .B(n42723), .C(n42724), .D(n37672), 
         .Z(n37686)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25753_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_94 (.A(n42803), .B(n36746), .C(n37252), .D(n109_adj_219), 
         .Z(n36756)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_94.init = 16'hfffe;
    LUT4 i1_4_lut_adj_95 (.A(n113_adj_222), .B(n42812), .C(n128_adj_232), 
         .D(n130_adj_233), .Z(n36744)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_95.init = 16'hfffe;
    LUT4 div_4016_LessThan_1658_i45_2_lut (.A(n2567), .B(n128_adj_232), 
         .Z(n45_adj_304)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i45_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_96 (.A(n108), .B(n42810), .C(n127_adj_231), .D(n129), 
         .Z(n36746)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_96.init = 16'hfffe;
    LUT4 div_4016_LessThan_2246_i47_2_lut_rep_956 (.A(n3439), .B(n121_adj_227), 
         .Z(n42655)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i47_2_lut_rep_956.init = 16'h6666;
    LUT4 div_4016_LessThan_2918_i31_2_lut_rep_824 (.A(n4443), .B(n121_adj_227), 
         .Z(n42523)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i31_2_lut_rep_824.init = 16'h6666;
    LUT4 i25099_3_lut (.A(\U[10] [16]), .B(\U[11] [16]), .C(i[0]), .Z(n40359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25099_3_lut.init = 16'hcaca;
    FD1P3IX x_3___i126 (.D(n5496), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i126.GSR = "ENABLED";
    LUT4 div_4016_LessThan_1862_i55_2_lut_rep_1006 (.A(n2865), .B(n121_adj_227), 
         .Z(n42705)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i55_2_lut_rep_1006.init = 16'h6666;
    LUT4 i25098_3_lut (.A(\U[8] [16]), .B(\U[9] [16]), .C(i[0]), .Z(n40358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25098_3_lut.init = 16'hcaca;
    LUT4 i25296_3_lut (.A(\U[14] [29]), .B(\U[15] [29]), .C(i[0]), .Z(n40556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25296_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1658_i40_4_lut (.A(n132), .B(n131_adj_234), .C(n2570), 
         .D(n876), .Z(n40)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i40_4_lut.init = 16'h0c8e;
    L6MUX21 i24868 (.D0(n40126), .D1(n40127), .SD(n9901), .Z(n5491));
    LUT4 i24013_3_lut_4_lut (.A(n4549), .B(n115_adj_223), .C(n21_adj_647), 
         .D(n42499), .Z(n39273)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24013_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_1862_i50_3_lut_3_lut (.A(n2865), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n50_adj_336)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i50_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i24883 (.D0(n40141), .D1(n40142), .SD(n9901), .Z(n5490));
    LUT4 div_4016_LessThan_2918_i26_3_lut_3_lut (.A(n4443), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n26_adj_619)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i26_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i24898 (.D0(n40156), .D1(n40157), .SD(n9901), .Z(n5489));
    LUT4 i1_2_lut_adj_97 (.A(n124_adj_229), .B(n126), .Z(n37252)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_97.init = 16'heeee;
    LUT4 i1_4_lut_adj_98 (.A(done_N_1934), .B(done_c), .C(done_N_1932), 
         .D(done_N_1931), .Z(done_N_1928)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i1_4_lut_adj_98.init = 16'heeea;
    LUT4 i25097_3_lut (.A(\U[6] [16]), .B(\U[7] [16]), .C(i[0]), .Z(n40357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25097_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2918_i33_2_lut_rep_825 (.A(n4442), .B(n120), 
         .Z(n42524)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i33_2_lut_rep_825.init = 16'h6666;
    L6MUX21 i24913 (.D0(n40171), .D1(n40172), .SD(n9901), .Z(n5488));
    LUT4 div_4016_i362_4_lut (.A(n35974), .B(n62_adj_800), .C(n42777), 
         .D(n131_adj_234), .Z(n35964)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i362_4_lut.init = 16'ha6a9;
    LUT4 i25893_4_lut (.A(n42721), .B(n42726), .C(n42728), .D(n47_adj_306), 
         .Z(n40080)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25893_4_lut.init = 16'haaab;
    LUT4 div_4016_LessThan_1862_i53_2_lut_rep_1007 (.A(n2866), .B(n122_adj_228), 
         .Z(n42706)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i53_2_lut_rep_1007.init = 16'h6666;
    LUT4 div_4016_LessThan_1658_i47_2_lut (.A(n2566), .B(n127_adj_231), 
         .Z(n47_adj_306)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i47_2_lut.init = 16'h6666;
    FD1P3IX x_3___i127 (.D(n5495), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i127.GSR = "ENABLED";
    LUT4 i25096_3_lut (.A(\U[4] [16]), .B(\U[5] [16]), .C(i[0]), .Z(n40356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25096_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2993_i37_2_lut_rep_799 (.A(n4551), .B(n117), 
         .Z(n42498)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i37_2_lut_rep_799.init = 16'h6666;
    LUT4 i1_4_lut_adj_99 (.A(n36882), .B(n30923), .C(n36946), .D(n36872), 
         .Z(n30872)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_99.init = 16'hfffe;
    L6MUX21 i24928 (.D0(n40186), .D1(n40187), .SD(n9901), .Z(n5487));
    LUT4 i25295_3_lut (.A(\U[12] [29]), .B(\U[13] [29]), .C(i[0]), .Z(n40555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25295_3_lut.init = 16'hcaca;
    L6MUX21 i24943 (.D0(n40201), .D1(n40202), .SD(n9901), .Z(n5486));
    LUT4 div_4016_LessThan_3137_i46_3_lut_3_lut (.A(n4756), .B(n107_adj_218), 
         .C(n44_adj_727), .Z(n46_adj_728)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i46_3_lut_3_lut.init = 16'hd4d4;
    FD1P3IX x_3___i128 (.D(n5494), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [31]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i128.GSR = "ENABLED";
    LUT4 i25929_4_lut (.A(n42556), .B(n42555), .C(n42557), .D(n38815), 
         .Z(n38840)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25929_4_lut.init = 16'hfeff;
    L6MUX21 i24958 (.D0(n40216), .D1(n40217), .SD(n9901), .Z(n5485));
    LUT4 div_4016_LessThan_3206_i7_4_lut (.A(n4779), .B(n129), .C(n22269), 
         .D(n4783), .Z(n7_adj_741)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i7_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2246_i42_3_lut_3_lut (.A(n3439), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n42_adj_409)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i42_3_lut_3_lut.init = 16'hd4d4;
    FD1P3IX x_3___i1 (.D(n5525), .SP(clk_c_enable_829), .CD(n31084), .CK(clk_c), 
            .Q(\x[3] [0]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i1.GSR = "ENABLED";
    LUT4 i25095_3_lut (.A(\U[2] [16]), .B(\U[3] [16]), .C(i[0]), .Z(n40355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25095_3_lut.init = 16'hcaca;
    LUT4 i22530_2_lut_3_lut_4_lut (.A(n2866), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n2865), .Z(n37790)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22530_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i23555_4_lut (.A(n42558), .B(n42560), .C(n42559), .D(n38799), 
         .Z(n38815)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23555_4_lut.init = 16'h1011;
    LUT4 i25094_3_lut (.A(\U[0] [16]), .B(\U[1] [16]), .C(i[0]), .Z(n40354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25094_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2918_i28_3_lut_3_lut (.A(n4442), .B(n120), .C(n26_adj_619), 
         .Z(n28_adj_620)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23539_4_lut (.A(n42561), .B(n39_adj_565), .C(n27_adj_556), .D(n38752), 
         .Z(n38799)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23539_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_2918_i27_2_lut_rep_826 (.A(n4445), .B(n123), 
         .Z(n42525)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i27_2_lut_rep_826.init = 16'h6666;
    LUT4 i1_2_lut_adj_100 (.A(n128_adj_232), .B(n30872), .Z(n30968)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_100.init = 16'heeee;
    LUT4 div_4016_LessThan_2246_i49_2_lut_rep_957 (.A(n3438), .B(n120), 
         .Z(n42656)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i49_2_lut_rep_957.init = 16'h6666;
    L6MUX21 i24973 (.D0(n40231), .D1(n40232), .SD(n9901), .Z(n5484));
    LUT4 i1_2_lut_adj_101 (.A(n126), .B(n30881), .Z(n30878)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_101.init = 16'heeee;
    LUT4 i1_2_lut_adj_102 (.A(n124_adj_229), .B(n30887), .Z(n30884)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_102.init = 16'heeee;
    LUT4 div_4016_LessThan_3137_i55_2_lut_rep_747 (.A(n4755), .B(n106_adj_217), 
         .Z(n42446)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i55_2_lut_rep_747.init = 16'h6666;
    LUT4 i25294_3_lut (.A(\U[10] [29]), .B(\U[11] [29]), .C(i[0]), .Z(n40554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25294_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1862_i51_2_lut_rep_1008 (.A(n2867), .B(n123), 
         .Z(n42707)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i51_2_lut_rep_1008.init = 16'h6666;
    L6MUX21 i24988 (.D0(n40246), .D1(n40247), .SD(n9901), .Z(n5483));
    L6MUX21 i25003 (.D0(n40261), .D1(n40262), .SD(n9901), .Z(n5482));
    LUT4 div_4016_LessThan_1862_i48_3_lut_3_lut (.A(n2867), .B(n123), .C(n40_adj_330), 
         .Z(n48_adj_335)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 select_5271_Select_31_i5_4_lut (.A(n70), .B(i[31]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[31])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_31_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_i3317_4_lut (.A(n64_adj_246), .B(n22281), .C(n42786), 
         .D(n30881), .Z(n5500)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3317_4_lut.init = 16'hc0c5;
    LUT4 i23890_2_lut_3_lut_4_lut (.A(n4445), .B(n123), .C(n111), .D(n4433), 
         .Z(n39150)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23890_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i24438_2_lut_3_lut_4_lut (.A(n4755), .B(n106_adj_217), .C(n105), 
         .D(n4754), .Z(n39698)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24438_2_lut_3_lut_4_lut.init = 16'h9009;
    FD1P3AX U_15___i511 (.D(\U[0] [30]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [30]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i511.GSR = "ENABLED";
    FD1P3AX U_15___i510 (.D(\U[0] [29]), .SP(clk_c_enable_831), .CK(clk_c), 
            .Q(\U[0] [29]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam U_15___i510.GSR = "ENABLED";
    LUT4 select_5271_Select_30_i5_4_lut (.A(n73_adj_95), .B(i[30]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[30])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_30_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_2246_i44_3_lut_3_lut (.A(n3438), .B(n120), .C(n42_adj_409), 
         .Z(n44_adj_410)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25814_4_lut (.A(n42730), .B(n42731), .C(n42732), .D(n37623), 
         .Z(n37637)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25814_4_lut.init = 16'hfffe;
    L6MUX21 i25018 (.D0(n40276), .D1(n40277), .SD(n9901), .Z(n5481));
    LUT4 i1_2_lut_adj_103 (.A(n122_adj_228), .B(n30893), .Z(n30890)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_103.init = 16'heeee;
    LUT4 select_5271_Select_29_i5_4_lut (.A(n76_adj_101), .B(i[29]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[29])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_29_i5_4_lut.init = 16'heca0;
    OB x_out_pad_125 (.I(x_out_c_125), .O(x_out[125]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_126 (.I(x_out_c_126), .O(x_out[126]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB x_out_pad_127 (.I(x_out_c_127), .O(x_out[127]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(14[24:29])
    OB done_pad (.I(done_c), .O(done));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(12[24:28])
    LUT4 i22521_3_lut_4_lut (.A(n2867), .B(n123), .C(n41), .D(n42708), 
         .Z(n37781)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22521_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_1553_i47_2_lut (.A(n2410), .B(n128_adj_232), 
         .Z(n47)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i47_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_1862_i49_2_lut_rep_1009 (.A(n2868), .B(n124_adj_229), 
         .Z(n42708)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i49_2_lut_rep_1009.init = 16'h6666;
    LUT4 i25086_3_lut (.A(\U[14] [15]), .B(\U[15] [15]), .C(i[0]), .Z(n40346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25086_3_lut.init = 16'hcaca;
    L6MUX21 i25033 (.D0(n40291), .D1(n40292), .SD(n9901), .Z(n5480));
    L6MUX21 i25048 (.D0(n40306), .D1(n40307), .SD(n9901), .Z(n5479));
    L6MUX21 i25063 (.D0(n40321), .D1(n40322), .SD(n9901), .Z(n5478));
    LUT4 i1_2_lut_adj_104 (.A(n118_adj_225), .B(n30905), .Z(n30902)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_104.init = 16'heeee;
    LUT4 select_5271_Select_28_i5_4_lut (.A(n79_adj_98), .B(i[28]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_28_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_1862_i40_3_lut_3_lut (.A(n2868), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n40_adj_330)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25085_3_lut (.A(\U[12] [15]), .B(\U[13] [15]), .C(i[0]), .Z(n40345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25085_3_lut.init = 16'hcaca;
    L6MUX21 i25078 (.D0(n40336), .D1(n40337), .SD(n9901), .Z(n5477));
    LUT4 i1_4_lut_adj_105 (.A(n36926), .B(n30929), .C(n36918), .D(n36916), 
         .Z(n30881)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_105.init = 16'hfffe;
    LUT4 div_4016_LessThan_2918_i25_2_lut_rep_827 (.A(n4446), .B(n124_adj_229), 
         .Z(n42526)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i25_2_lut_rep_827.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i22_3_lut (.A(n106_adj_217), .B(n105), .C(n55_adj_787), 
         .Z(n22_adj_756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i22_3_lut.init = 16'hcaca;
    L6MUX21 i25093 (.D0(n40351), .D1(n40352), .SD(n9901), .Z(n5476));
    L6MUX21 i25108 (.D0(n40366), .D1(n40367), .SD(n9901), .Z(n5475));
    LUT4 i1_2_lut_adj_106 (.A(n116_adj_224), .B(n30911), .Z(n30908)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_106.init = 16'heeee;
    LUT4 i1_2_lut_adj_107 (.A(n114), .B(n30917), .Z(n30914)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_107.init = 16'heeee;
    L6MUX21 i25123 (.D0(n40381), .D1(n40382), .SD(n9901), .Z(n5474));
    L6MUX21 i25138 (.D0(n40396), .D1(n40397), .SD(n9901), .Z(n5473));
    LUT4 div_4016_LessThan_2918_i16_3_lut_3_lut (.A(n4446), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n16_adj_612)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i16_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i25153 (.D0(n40411), .D1(n40412), .SD(n9901), .Z(n5472));
    IB U_in_pad_41 (.I(U_in[41]), .O(U_in_c_41));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_40 (.I(U_in[40]), .O(U_in_c_40));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_39 (.I(U_in[39]), .O(U_in_c_39));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_38 (.I(U_in[38]), .O(U_in_c_38));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_37 (.I(U_in[37]), .O(U_in_c_37));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_36 (.I(U_in[36]), .O(U_in_c_36));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_35 (.I(U_in[35]), .O(U_in_c_35));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_34 (.I(U_in[34]), .O(U_in_c_34));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_33 (.I(U_in[33]), .O(U_in_c_33));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_32 (.I(U_in[32]), .O(U_in_c_32));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_31 (.I(U_in[31]), .O(U_in_c_31));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_30 (.I(U_in[30]), .O(U_in_c_30));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_29 (.I(U_in[29]), .O(U_in_c_29));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_28 (.I(U_in[28]), .O(U_in_c_28));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_27 (.I(U_in[27]), .O(U_in_c_27));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_26 (.I(U_in[26]), .O(U_in_c_26));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_25 (.I(U_in[25]), .O(U_in_c_25));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_24 (.I(U_in[24]), .O(U_in_c_24));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_23 (.I(U_in[23]), .O(U_in_c_23));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_22 (.I(U_in[22]), .O(U_in_c_22));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_21 (.I(U_in[21]), .O(U_in_c_21));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_20 (.I(U_in[20]), .O(U_in_c_20));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_19 (.I(U_in[19]), .O(U_in_c_19));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_18 (.I(U_in[18]), .O(U_in_c_18));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_17 (.I(U_in[17]), .O(U_in_c_17));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_16 (.I(U_in[16]), .O(U_in_c_16));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_15 (.I(U_in[15]), .O(U_in_c_15));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_14 (.I(U_in[14]), .O(U_in_c_14));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_13 (.I(U_in[13]), .O(U_in_c_13));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_12 (.I(U_in[12]), .O(U_in_c_12));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_11 (.I(U_in[11]), .O(U_in_c_11));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_10 (.I(U_in[10]), .O(U_in_c_10));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_9 (.I(U_in[9]), .O(U_in_c_9));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_8 (.I(U_in[8]), .O(U_in_c_8));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_7 (.I(U_in[7]), .O(U_in_c_7));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_6 (.I(U_in[6]), .O(U_in_c_6));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_5 (.I(U_in[5]), .O(U_in_c_5));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_4 (.I(U_in[4]), .O(U_in_c_4));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_3 (.I(U_in[3]), .O(U_in_c_3));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_2 (.I(U_in[2]), .O(U_in_c_2));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_1 (.I(U_in[1]), .O(U_in_c_1));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB U_in_pad_0 (.I(U_in[0]), .O(U_in_c_0));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(9[24:28])
    IB y_in_pad_127 (.I(y_in[127]), .O(y_in_c_127));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_126 (.I(y_in[126]), .O(y_in_c_126));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_125 (.I(y_in[125]), .O(y_in_c_125));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_124 (.I(y_in[124]), .O(y_in_c_124));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_123 (.I(y_in[123]), .O(y_in_c_123));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_122 (.I(y_in[122]), .O(y_in_c_122));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_121 (.I(y_in[121]), .O(y_in_c_121));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_120 (.I(y_in[120]), .O(y_in_c_120));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_119 (.I(y_in[119]), .O(y_in_c_119));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_118 (.I(y_in[118]), .O(y_in_c_118));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_117 (.I(y_in[117]), .O(y_in_c_117));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_116 (.I(y_in[116]), .O(y_in_c_116));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_115 (.I(y_in[115]), .O(y_in_c_115));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_114 (.I(y_in[114]), .O(y_in_c_114));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_113 (.I(y_in[113]), .O(y_in_c_113));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_112 (.I(y_in[112]), .O(y_in_c_112));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_111 (.I(y_in[111]), .O(y_in_c_111));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_110 (.I(y_in[110]), .O(y_in_c_110));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_109 (.I(y_in[109]), .O(y_in_c_109));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_108 (.I(y_in[108]), .O(y_in_c_108));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_107 (.I(y_in[107]), .O(y_in_c_107));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_106 (.I(y_in[106]), .O(y_in_c_106));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_105 (.I(y_in[105]), .O(y_in_c_105));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_104 (.I(y_in[104]), .O(y_in_c_104));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_103 (.I(y_in[103]), .O(y_in_c_103));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_102 (.I(y_in[102]), .O(y_in_c_102));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_101 (.I(y_in[101]), .O(y_in_c_101));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_100 (.I(y_in[100]), .O(y_in_c_100));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_99 (.I(y_in[99]), .O(y_in_c_99));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_98 (.I(y_in[98]), .O(y_in_c_98));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_97 (.I(y_in[97]), .O(y_in_c_97));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_96 (.I(y_in[96]), .O(y_in_c_96));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_95 (.I(y_in[95]), .O(y_in_c_95));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_94 (.I(y_in[94]), .O(y_in_c_94));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_93 (.I(y_in[93]), .O(y_in_c_93));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_92 (.I(y_in[92]), .O(y_in_c_92));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_91 (.I(y_in[91]), .O(y_in_c_91));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_90 (.I(y_in[90]), .O(y_in_c_90));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_89 (.I(y_in[89]), .O(y_in_c_89));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_88 (.I(y_in[88]), .O(y_in_c_88));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_87 (.I(y_in[87]), .O(y_in_c_87));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_86 (.I(y_in[86]), .O(y_in_c_86));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_85 (.I(y_in[85]), .O(y_in_c_85));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_84 (.I(y_in[84]), .O(y_in_c_84));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_83 (.I(y_in[83]), .O(y_in_c_83));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_82 (.I(y_in[82]), .O(y_in_c_82));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_81 (.I(y_in[81]), .O(y_in_c_81));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_80 (.I(y_in[80]), .O(y_in_c_80));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_79 (.I(y_in[79]), .O(y_in_c_79));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_78 (.I(y_in[78]), .O(y_in_c_78));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_77 (.I(y_in[77]), .O(y_in_c_77));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_76 (.I(y_in[76]), .O(y_in_c_76));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_75 (.I(y_in[75]), .O(y_in_c_75));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_74 (.I(y_in[74]), .O(y_in_c_74));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_73 (.I(y_in[73]), .O(y_in_c_73));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_72 (.I(y_in[72]), .O(y_in_c_72));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_71 (.I(y_in[71]), .O(y_in_c_71));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_70 (.I(y_in[70]), .O(y_in_c_70));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_69 (.I(y_in[69]), .O(y_in_c_69));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_68 (.I(y_in[68]), .O(y_in_c_68));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_67 (.I(y_in[67]), .O(y_in_c_67));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_66 (.I(y_in[66]), .O(y_in_c_66));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_65 (.I(y_in[65]), .O(y_in_c_65));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_64 (.I(y_in[64]), .O(y_in_c_64));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_63 (.I(y_in[63]), .O(y_in_c_63));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_62 (.I(y_in[62]), .O(y_in_c_62));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_61 (.I(y_in[61]), .O(y_in_c_61));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_60 (.I(y_in[60]), .O(y_in_c_60));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_59 (.I(y_in[59]), .O(y_in_c_59));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_58 (.I(y_in[58]), .O(y_in_c_58));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_57 (.I(y_in[57]), .O(y_in_c_57));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_56 (.I(y_in[56]), .O(y_in_c_56));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_55 (.I(y_in[55]), .O(y_in_c_55));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_54 (.I(y_in[54]), .O(y_in_c_54));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_53 (.I(y_in[53]), .O(y_in_c_53));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_52 (.I(y_in[52]), .O(y_in_c_52));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_51 (.I(y_in[51]), .O(y_in_c_51));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_50 (.I(y_in[50]), .O(y_in_c_50));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_49 (.I(y_in[49]), .O(y_in_c_49));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_48 (.I(y_in[48]), .O(y_in_c_48));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_47 (.I(y_in[47]), .O(y_in_c_47));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_46 (.I(y_in[46]), .O(y_in_c_46));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_45 (.I(y_in[45]), .O(y_in_c_45));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_44 (.I(y_in[44]), .O(y_in_c_44));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_43 (.I(y_in[43]), .O(y_in_c_43));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_42 (.I(y_in[42]), .O(y_in_c_42));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_41 (.I(y_in[41]), .O(y_in_c_41));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_40 (.I(y_in[40]), .O(y_in_c_40));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_39 (.I(y_in[39]), .O(y_in_c_39));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_38 (.I(y_in[38]), .O(y_in_c_38));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_37 (.I(y_in[37]), .O(y_in_c_37));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_36 (.I(y_in[36]), .O(y_in_c_36));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_35 (.I(y_in[35]), .O(y_in_c_35));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_34 (.I(y_in[34]), .O(y_in_c_34));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_33 (.I(y_in[33]), .O(y_in_c_33));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_32 (.I(y_in[32]), .O(y_in_c_32));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_31 (.I(y_in[31]), .O(y_in_c_31));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_30 (.I(y_in[30]), .O(y_in_c_30));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_29 (.I(y_in[29]), .O(y_in_c_29));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_28 (.I(y_in[28]), .O(y_in_c_28));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_27 (.I(y_in[27]), .O(y_in_c_27));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_26 (.I(y_in[26]), .O(y_in_c_26));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_25 (.I(y_in[25]), .O(y_in_c_25));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_24 (.I(y_in[24]), .O(y_in_c_24));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_23 (.I(y_in[23]), .O(y_in_c_23));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_22 (.I(y_in[22]), .O(y_in_c_22));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_21 (.I(y_in[21]), .O(y_in_c_21));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_20 (.I(y_in[20]), .O(y_in_c_20));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_19 (.I(y_in[19]), .O(y_in_c_19));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_18 (.I(y_in[18]), .O(y_in_c_18));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_17 (.I(y_in[17]), .O(y_in_c_17));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_16 (.I(y_in[16]), .O(y_in_c_16));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_15 (.I(y_in[15]), .O(y_in_c_15));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_14 (.I(y_in[14]), .O(y_in_c_14));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_13 (.I(y_in[13]), .O(y_in_c_13));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_12 (.I(y_in[12]), .O(y_in_c_12));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_11 (.I(y_in[11]), .O(y_in_c_11));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_10 (.I(y_in[10]), .O(y_in_c_10));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_9 (.I(y_in[9]), .O(y_in_c_9));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_8 (.I(y_in[8]), .O(y_in_c_8));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_7 (.I(y_in[7]), .O(y_in_c_7));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_6 (.I(y_in[6]), .O(y_in_c_6));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_5 (.I(y_in[5]), .O(y_in_c_5));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_4 (.I(y_in[4]), .O(y_in_c_4));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_3 (.I(y_in[3]), .O(y_in_c_3));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_2 (.I(y_in[2]), .O(y_in_c_2));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_1 (.I(y_in[1]), .O(y_in_c_1));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    IB y_in_pad_0 (.I(y_in[0]), .O(y_in_c_0));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(11[24:28])
    LUT4 div_4016_LessThan_2918_i19_2_lut_rep_828 (.A(n4449), .B(n127_adj_231), 
         .Z(n42527)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i19_2_lut_rep_828.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i32_3_lut_3_lut (.A(n4551), .B(n117), .C(n20_adj_646), 
         .Z(n32_adj_653)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i32_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i25168 (.D0(n40426), .D1(n40427), .SD(n9901), .Z(n5471));
    LUT4 div_4016_LessThan_2918_i12_4_lut (.A(n132), .B(n131_adj_234), .C(n4453), 
         .D(n890), .Z(n12_adj_609)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i12_4_lut.init = 16'h0c8e;
    LUT4 div_4016_mux_5_i29_3_lut (.A(n5463), .B(n71_adj_196), .C(n5460), 
         .Z(n104_adj_216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i29_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_108 (.A(n112_adj_221), .B(n30923), .Z(n30920)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_108.init = 16'heeee;
    LUT4 div_4016_LessThan_1862_i47_2_lut_rep_1010 (.A(n2869), .B(n125_adj_230), 
         .Z(n42709)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i47_2_lut_rep_1010.init = 16'h6666;
    L6MUX21 i25183 (.D0(n40441), .D1(n40442), .SD(n9901), .Z(n5470));
    LUT4 div_4016_LessThan_2513_i64_4_lut (.A(n58_adj_490), .B(n62_adj_492), 
         .C(n42603), .D(n38479), .Z(n64_adj_493)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2513_i64_4_lut.init = 16'hcacc;
    LUT4 div_4016_LessThan_1862_i44_3_lut_3_lut (.A(n2869), .B(n125_adj_230), 
         .C(n42_adj_331), .Z(n44_adj_333)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22508_3_lut_4_lut (.A(n2869), .B(n125_adj_230), .C(n43_adj_332), 
         .D(n42710), .Z(n37768)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22508_3_lut_4_lut.init = 16'h0009;
    L6MUX21 i25198 (.D0(n40456), .D1(n40457), .SD(n9901), .Z(n5469));
    LUT4 select_5271_Select_27_i5_4_lut (.A(n82_adj_104), .B(i[27]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[27])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_27_i5_4_lut.init = 16'heca0;
    LUT4 select_5271_Select_26_i5_4_lut (.A(n85_adj_91), .B(i[26]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[26])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_26_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_1553_i49_2_lut (.A(n2409), .B(n127_adj_231), 
         .Z(n49_adj_293)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i49_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i57_4_lut (.A(n4754), .B(n104_adj_216), 
         .C(n22244), .D(n4783), .Z(n57_adj_789)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i57_4_lut.init = 16'h663c;
    LUT4 i23192_4_lut (.A(n42606), .B(n42607), .C(n42609), .D(n38429), 
         .Z(n38452)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23192_4_lut.init = 16'h0100;
    L6MUX21 i25213 (.D0(n40471), .D1(n40472), .SD(n9901), .Z(n5468));
    LUT4 i23169_4_lut (.A(n42608), .B(n42610), .C(n45_adj_483), .D(n38414), 
         .Z(n38429)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23169_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_1446_i61_2_lut (.A(n2244), .B(n122_adj_228), 
         .Z(n37578)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i61_2_lut.init = 16'h9999;
    LUT4 div_4016_LessThan_3137_i49_2_lut_rep_748 (.A(n4758), .B(n109_adj_219), 
         .Z(n42447)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i49_2_lut_rep_748.init = 16'h6666;
    LUT4 select_5271_Select_25_i5_4_lut (.A(n88_adj_151), .B(i[25]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[25])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_25_i5_4_lut.init = 16'heca0;
    LUT4 i23135_4_lut (.A(n42613), .B(n42615), .C(n33_adj_476), .D(n38382), 
         .Z(n38395)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23135_4_lut.init = 16'h1011;
    L6MUX21 i25228 (.D0(n40486), .D1(n40487), .SD(n9901), .Z(n5467));
    LUT4 i23122_4_lut (.A(n42617), .B(n42616), .C(n42618), .D(n38373), 
         .Z(n38382)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23122_4_lut.init = 16'h1011;
    LUT4 div_4016_mux_5_i27_3_lut (.A(n5465), .B(n73_adj_197), .C(n5460), 
         .Z(n106_adj_217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i27_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1862_i45_2_lut_rep_1011 (.A(n2870), .B(n126), 
         .Z(n42710)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i45_2_lut_rep_1011.init = 16'h6666;
    L6MUX21 i25243 (.D0(n40501), .D1(n40502), .SD(n9901), .Z(n5466));
    L6MUX21 i25258 (.D0(n40516), .D1(n40517), .SD(n9901), .Z(n5465));
    LUT4 i25939_4_lut (.A(n42737), .B(n37578), .C(n42738), .D(n37576), 
         .Z(n37588)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25939_4_lut.init = 16'hbfbb;
    LUT4 div_4016_LessThan_2246_i45_2_lut_rep_958 (.A(n3440), .B(n122_adj_228), 
         .Z(n42657)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i45_2_lut_rep_958.init = 16'h6666;
    LUT4 select_5271_Select_24_i5_4_lut (.A(n91_adj_160), .B(i[24]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[24])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_24_i5_4_lut.init = 16'heca0;
    L6MUX21 i25273 (.D0(n40531), .D1(n40532), .SD(n9901), .Z(n5464));
    L6MUX21 i25288 (.D0(n40546), .D1(n40547), .SD(n9901), .Z(n5463));
    LUT4 div_4016_LessThan_1862_i42_3_lut_3_lut (.A(n2870), .B(n126), .C(n127_adj_231), 
         .Z(n42_adj_331)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25293_3_lut (.A(\U[8] [29]), .B(\U[9] [29]), .C(i[0]), .Z(n40553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25293_3_lut.init = 16'hcaca;
    L6MUX21 i25303 (.D0(n40561), .D1(n40562), .SD(n9901), .Z(n5462));
    LUT4 i25084_3_lut (.A(\U[10] [15]), .B(\U[11] [15]), .C(i[0]), .Z(n40344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25084_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2993_i16_3_lut_3_lut (.A(n4560), .B(n126), .C(n127_adj_231), 
         .Z(n16_adj_644)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i16_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i25318 (.D0(n40576), .D1(n40577), .SD(n9901), .Z(n5461));
    LUT4 i1_2_lut_adj_109 (.A(n110_adj_220), .B(n30929), .Z(n30926)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_109.init = 16'heeee;
    LUT4 i25292_3_lut (.A(\U[6] [29]), .B(\U[7] [29]), .C(i[0]), .Z(n40552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25292_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2918_i21_2_lut_rep_829 (.A(n4448), .B(n126), 
         .Z(n42528)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i21_2_lut_rep_829.init = 16'h6666;
    LUT4 i23783_2_lut_3_lut_4_lut (.A(n4448), .B(n126), .C(n127_adj_231), 
         .D(n4449), .Z(n39043)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23783_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 select_5271_Select_23_i5_4_lut (.A(n94_adj_152), .B(i[23]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[23])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_23_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_1446_i51_2_lut (.A(n2249), .B(n127_adj_231), 
         .Z(n51_adj_282)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i51_2_lut.init = 16'h6666;
    L6MUX21 i24866 (.D0(n40122), .D1(n40123), .SD(n9902), .Z(n40126));
    LUT4 i1_4_lut_adj_110 (.A(n42808), .B(n42797), .C(n42798), .D(n42796), 
         .Z(n30929)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_110.init = 16'hfffe;
    LUT4 mux_4010_i26_4_lut (.A(n88), .B(n36694), .C(n15805), .D(i[1]), 
         .Z(n5331)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i26_4_lut.init = 16'hca0a;
    LUT4 i25291_3_lut (.A(\U[4] [29]), .B(\U[5] [29]), .C(i[0]), .Z(n40551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25291_3_lut.init = 16'hcaca;
    LUT4 i25083_3_lut (.A(\U[8] [15]), .B(\U[9] [15]), .C(i[0]), .Z(n40343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25083_3_lut.init = 16'hcaca;
    LUT4 i22492_3_lut_4_lut (.A(n2873), .B(n129), .C(n130_adj_233), .D(n2874), 
         .Z(n37752)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22492_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_mux_5_i28_3_lut (.A(n5464), .B(n72), .C(n5460), .Z(n105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i28_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1862_i38_3_lut_3_lut (.A(n2873), .B(n129), .C(n130_adj_233), 
         .Z(n38_adj_329)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1862_i38_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i24867 (.D0(n40124), .D1(n40125), .SD(n9902), .Z(n40127));
    L6MUX21 i24881 (.D0(n40137), .D1(n40138), .SD(n9902), .Z(n40141));
    LUT4 div_4016_LessThan_2918_i18_3_lut_3_lut (.A(n4448), .B(n126), .C(n127_adj_231), 
         .Z(n18_adj_614)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i15_2_lut_rep_830 (.A(n4451), .B(n129), 
         .Z(n42529)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i15_2_lut_rep_830.init = 16'h6666;
    LUT4 i23464_4_lut (.A(n38723), .B(n42569), .C(n42570), .D(n38707), 
         .Z(n38724)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23464_4_lut.init = 16'h0002;
    L6MUX21 i24882 (.D0(n40139), .D1(n40140), .SD(n9902), .Z(n40142));
    LUT4 div_4016_LessThan_2918_i14_3_lut_3_lut (.A(n4451), .B(n129), .C(n130_adj_233), 
         .Z(n14_adj_611)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i14_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25290_3_lut (.A(\U[2] [29]), .B(\U[3] [29]), .C(i[0]), .Z(n40550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25290_3_lut.init = 16'hcaca;
    LUT4 i25585_4_lut_4_lut (.A(n42711), .B(n37742), .C(n48_adj_320), 
         .D(n38), .Z(n60_adj_326)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25585_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25951_4_lut (.A(n42744), .B(n42745), .C(n42747), .D(n51), 
         .Z(n37548)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25951_4_lut.init = 16'haaab;
    LUT4 i25583_4_lut_4_lut (.A(n42712), .B(n37733), .C(n54_adj_323), 
         .D(n40_adj_316), .Z(n56_adj_324)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25583_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25289_3_lut (.A(\U[0] [29]), .B(\U[1] [29]), .C(i[0]), .Z(n40549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25289_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1337_i51_2_lut (.A(n2087), .B(n128_adj_232), 
         .Z(n51)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i51_2_lut.init = 16'h6666;
    LUT4 i25944_4_lut_4_lut (.A(n42712), .B(n37729), .C(n37742), .D(n42711), 
         .Z(n37746)) /* synthesis lut_function=(A ((D)+!C)+!A (B+((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25944_4_lut_4_lut.init = 16'hff4f;
    LUT4 i25680_4_lut_4_lut (.A(n42531), .B(n39017), .C(n54_adj_603), 
         .D(n18_adj_581), .Z(n56_adj_604)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25680_4_lut_4_lut.init = 16'hf4b0;
    LUT4 select_5271_Select_22_i5_4_lut (.A(n97_adj_153), .B(i[22]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[22])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_22_i5_4_lut.init = 16'heca0;
    LUT4 i25895_4_lut_4_lut (.A(n42531), .B(n39004), .C(n42533), .D(n42530), 
         .Z(n39028)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25895_4_lut_4_lut.init = 16'hff04;
    LUT4 i25082_3_lut (.A(\U[6] [15]), .B(\U[7] [15]), .C(i[0]), .Z(n40342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25082_3_lut.init = 16'hcaca;
    LUT4 i25081_3_lut (.A(\U[4] [15]), .B(\U[5] [15]), .C(i[0]), .Z(n40341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25081_3_lut.init = 16'hcaca;
    L6MUX21 i24896 (.D0(n40152), .D1(n40153), .SD(n9902), .Z(n40156));
    L6MUX21 i24897 (.D0(n40154), .D1(n40155), .SD(n9902), .Z(n40157));
    L6MUX21 i24911 (.D0(n40167), .D1(n40168), .SD(n9902), .Z(n40171));
    LUT4 i23422_4_lut (.A(n42574), .B(n42576), .C(n42575), .D(n38661), 
         .Z(n38682)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23422_4_lut.init = 16'h0100;
    L6MUX21 i24912 (.D0(n40169), .D1(n40170), .SD(n9902), .Z(n40172));
    L6MUX21 i24926 (.D0(n40182), .D1(n40183), .SD(n9902), .Z(n40186));
    LUT4 div_4016_LessThan_1337_i53_2_lut (.A(n2086), .B(n127_adj_231), 
         .Z(n53)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1337_i53_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_1761_i63_2_lut_rep_1012 (.A(n2711), .B(n118_adj_225), 
         .Z(n42711)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i63_2_lut_rep_1012.init = 16'h6666;
    L6MUX21 i24927 (.D0(n40184), .D1(n40185), .SD(n9902), .Z(n40187));
    LUT4 i23751_4_lut_4_lut (.A(n42531), .B(n38990), .C(n42532), .D(n42533), 
         .Z(n39011)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23751_4_lut_4_lut.init = 16'h0004;
    LUT4 select_5271_Select_21_i5_4_lut (.A(n100_adj_161), .B(i[21]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[21])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_21_i5_4_lut.init = 16'heca0;
    L6MUX21 i24941 (.D0(n40197), .D1(n40198), .SD(n9902), .Z(n40201));
    LUT4 i25839_3_lut_4_lut (.A(n4551), .B(n117), .C(n33_adj_654), .D(n42500), 
         .Z(n39257)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25839_3_lut_4_lut.init = 16'hfff6;
    L6MUX21 i24942 (.D0(n40199), .D1(n40200), .SD(n9902), .Z(n40202));
    LUT4 i25080_3_lut (.A(\U[2] [15]), .B(\U[3] [15]), .C(i[0]), .Z(n40340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25080_3_lut.init = 16'hcaca;
    LUT4 i25281_3_lut (.A(\U[14] [28]), .B(\U[15] [28]), .C(i[0]), .Z(n40541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25281_3_lut.init = 16'hcaca;
    LUT4 i23401_4_lut (.A(n42577), .B(n41_adj_537), .C(n42579), .D(n38644), 
         .Z(n38661)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23401_4_lut.init = 16'h1011;
    L6MUX21 i24956 (.D0(n40212), .D1(n40213), .SD(n9902), .Z(n40216));
    L6MUX21 i24957 (.D0(n40214), .D1(n40215), .SD(n9902), .Z(n40217));
    LUT4 div_4016_LessThan_881_i61_2_lut (.A(n1404), .B(n127_adj_231), .Z(n61)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_881_i61_2_lut.init = 16'h9999;
    L6MUX21 i24971 (.D0(n40227), .D1(n40228), .SD(n9902), .Z(n40231));
    LUT4 select_5271_Select_20_i5_4_lut (.A(n103_adj_92), .B(i[20]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[20])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_20_i5_4_lut.init = 16'heca0;
    LUT4 select_5271_Select_19_i5_4_lut (.A(n106_adj_49), .B(i[19]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[19])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_19_i5_4_lut.init = 16'heca0;
    L6MUX21 i24972 (.D0(n40229), .D1(n40230), .SD(n9902), .Z(n40232));
    LUT4 i25079_3_lut (.A(\U[0] [15]), .B(\U[1] [15]), .C(i[0]), .Z(n40339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25079_3_lut.init = 16'hcaca;
    L6MUX21 i24986 (.D0(n40242), .D1(n40243), .SD(n9902), .Z(n40246));
    LUT4 i23384_4_lut (.A(n42578), .B(n35_adj_533), .C(n42580), .D(n38629), 
         .Z(n38644)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23384_4_lut.init = 16'h0100;
    LUT4 i25280_3_lut (.A(\U[12] [28]), .B(\U[13] [28]), .C(i[0]), .Z(n40540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25280_3_lut.init = 16'hcaca;
    LUT4 i25852_4_lut (.A(n42764), .B(n61), .C(n42765), .D(n37431), 
         .Z(n37440)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25852_4_lut.init = 16'hbfbb;
    LUT4 div_4016_LessThan_2762_i39_2_lut (.A(n4208), .B(n119_adj_226), 
         .Z(n39_adj_565)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i39_2_lut.init = 16'h6666;
    L6MUX21 i24987 (.D0(n40244), .D1(n40245), .SD(n9902), .Z(n40247));
    L6MUX21 i25001 (.D0(n40257), .D1(n40258), .SD(n9902), .Z(n40261));
    LUT4 i25071_3_lut (.A(\U[14] [14]), .B(\U[15] [14]), .C(i[0]), .Z(n40331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25071_3_lut.init = 16'hcaca;
    LUT4 select_5271_Select_18_i5_4_lut (.A(n109_adj_106), .B(i[18]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[18])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_18_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_762_i56_4_lut (.A(n132), .B(n131_adj_234), .C(n1230), 
         .D(n682), .Z(n56_adj_237)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i56_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_1761_i48_3_lut_3_lut (.A(n2711), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n48_adj_320)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i48_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i25002 (.D0(n40259), .D1(n40260), .SD(n9902), .Z(n40262));
    L6MUX21 i25016 (.D0(n40272), .D1(n40273), .SD(n9902), .Z(n40276));
    LUT4 i25070_3_lut (.A(\U[12] [14]), .B(\U[13] [14]), .C(i[0]), .Z(n40330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25070_3_lut.init = 16'hcaca;
    L6MUX21 i25017 (.D0(n40274), .D1(n40275), .SD(n9902), .Z(n40277));
    LUT4 i23369_4_lut (.A(n42581), .B(n29_adj_529), .C(n42583), .D(n38616), 
         .Z(n38629)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23369_4_lut.init = 16'h5455;
    LUT4 i25682_4_lut_4_lut (.A(n42531), .B(n39015), .C(n56_adj_604), 
         .D(n34_adj_592), .Z(n58_adj_605)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25682_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i25279_3_lut (.A(\U[10] [28]), .B(\U[11] [28]), .C(i[0]), .Z(n40539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25279_3_lut.init = 16'hcaca;
    LUT4 i25864_4_lut (.A(n42766), .B(n42768), .C(n42767), .D(n57), 
         .Z(n37427)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25864_4_lut.init = 16'haaab;
    L6MUX21 i25031 (.D0(n40287), .D1(n40288), .SD(n9902), .Z(n40291));
    L6MUX21 i25032 (.D0(n40289), .D1(n40290), .SD(n9902), .Z(n40292));
    LUT4 div_4016_LessThan_762_i57_2_lut (.A(n1229), .B(n130_adj_233), .Z(n57)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_762_i57_2_lut.init = 16'h6666;
    L6MUX21 i25046 (.D0(n40302), .D1(n40303), .SD(n9902), .Z(n40306));
    LUT4 div_4016_LessThan_2762_i27_2_lut (.A(n4214), .B(n125_adj_230), 
         .Z(n27_adj_556)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i27_2_lut.init = 16'h6666;
    LUT4 i25069_3_lut (.A(\U[10] [14]), .B(\U[11] [14]), .C(i[0]), .Z(n40329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25069_3_lut.init = 16'hcaca;
    L6MUX21 i25047 (.D0(n40304), .D1(n40305), .SD(n9902), .Z(n40307));
    LUT4 i6999_2_lut (.A(i[0]), .B(i[2]), .Z(n9902)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[29:36])
    defparam i6999_2_lut.init = 16'h6666;
    LUT4 i23356_4_lut (.A(n42582), .B(n23_adj_525), .C(n42584), .D(n19_adj_522), 
         .Z(n38616)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23356_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_2681_i19_2_lut (.A(n4098), .B(n130_adj_233), 
         .Z(n19_adj_522)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i19_2_lut.init = 16'h6666;
    L6MUX21 i25061 (.D0(n40317), .D1(n40318), .SD(n9902), .Z(n40321));
    LUT4 div_4016_LessThan_1761_i59_2_lut_rep_1013 (.A(n2713), .B(n120), 
         .Z(n42712)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i59_2_lut_rep_1013.init = 16'h6666;
    LUT4 i22663_4_lut (.A(n42681), .B(n42682), .C(n42683), .D(n37908), 
         .Z(n37923)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22663_4_lut.init = 16'h0100;
    L6MUX21 i25062 (.D0(n40319), .D1(n40320), .SD(n9902), .Z(n40322));
    LUT4 div_4016_LessThan_2841_i63_2_lut_rep_831 (.A(n4313), .B(n106_adj_217), 
         .Z(n42530)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i63_2_lut_rep_831.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i39_2_lut_rep_800 (.A(n4550), .B(n116_adj_224), 
         .Z(n42499)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i39_2_lut_rep_800.init = 16'h6666;
    LUT4 i25068_3_lut (.A(\U[8] [14]), .B(\U[9] [14]), .C(i[0]), .Z(n40328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25068_3_lut.init = 16'hcaca;
    LUT4 i22648_4_lut (.A(n42684), .B(n42685), .C(n42687), .D(n37895), 
         .Z(n37908)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22648_4_lut.init = 16'h5455;
    LUT4 i22635_4_lut (.A(n42686), .B(n37), .C(n42688), .D(n33_adj_362), 
         .Z(n37895)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22635_4_lut.init = 16'h5554;
    L6MUX21 i25076 (.D0(n40332), .D1(n40333), .SD(n9902), .Z(n40336));
    L6MUX21 i25077 (.D0(n40334), .D1(n40335), .SD(n9902), .Z(n40337));
    LUT4 div_4016_LessThan_1761_i54_3_lut_3_lut (.A(n2713), .B(n120), .C(n52_adj_322), 
         .Z(n54_adj_323)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2058_i33_2_lut (.A(n3167), .B(n130_adj_233), 
         .Z(n33_adj_362)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i33_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2598_i64_4_lut (.A(n56_adj_516), .B(n62_adj_519), 
         .C(n42585), .D(n38597), .Z(n64_adj_520)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2598_i64_4_lut.init = 16'hcacc;
    L6MUX21 i25091 (.D0(n40347), .D1(n40348), .SD(n9902), .Z(n40351));
    LUT4 div_4016_LessThan_3137_i51_2_lut_rep_749 (.A(n4757), .B(n108), 
         .Z(n42448)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i51_2_lut_rep_749.init = 16'h6666;
    LUT4 i25770_4_lut (.A(n42442), .B(n42441), .C(n42443), .D(n39687), 
         .Z(n39714)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25770_4_lut.init = 16'hfeff;
    L6MUX21 i25092 (.D0(n40349), .D1(n40350), .SD(n9902), .Z(n40352));
    L6MUX21 i25106 (.D0(n40362), .D1(n40363), .SD(n9902), .Z(n40366));
    LUT4 select_5271_Select_17_i5_4_lut (.A(n112_adj_50), .B(i[17]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[17])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_17_i5_4_lut.init = 16'heca0;
    L6MUX21 i25107 (.D0(n40364), .D1(n40365), .SD(n9902), .Z(n40367));
    L6MUX21 i25121 (.D0(n40377), .D1(n40378), .SD(n9902), .Z(n40381));
    LUT4 i22583_4_lut (.A(n42695), .B(n42696), .C(n42697), .D(n37830), 
         .Z(n37843)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22583_4_lut.init = 16'h0001;
    LUT4 select_5271_Select_16_i5_4_lut (.A(n115_adj_52), .B(i[16]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[16])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_16_i5_4_lut.init = 16'heca0;
    LUT4 i22570_4_lut (.A(n42698), .B(n42699), .C(n41_adj_348), .D(n37819), 
         .Z(n37830)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22570_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_2841_i60_3_lut_3_lut (.A(n4313), .B(n106_adj_217), 
         .C(n32_adj_591), .Z(n60_adj_606)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i60_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 i25122 (.D0(n40379), .D1(n40380), .SD(n9902), .Z(n40382));
    LUT4 i24427_4_lut (.A(n42444), .B(n42446), .C(n42445), .D(n39667), 
         .Z(n39687)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24427_4_lut.init = 16'h1011;
    LUT4 i22559_4_lut (.A(n39_adj_346), .B(n42700), .C(n3022), .D(n130_adj_233), 
         .Z(n37819)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22559_4_lut.init = 16'h1001;
    L6MUX21 i25136 (.D0(n40392), .D1(n40393), .SD(n9902), .Z(n40396));
    LUT4 div_4016_LessThan_2841_i61_2_lut_rep_832 (.A(n4314), .B(n107_adj_218), 
         .Z(n42531)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i61_2_lut_rep_832.init = 16'h6666;
    L6MUX21 i25137 (.D0(n40394), .D1(n40395), .SD(n9902), .Z(n40397));
    LUT4 div_4016_LessThan_1761_i57_2_lut_rep_1014 (.A(n2714), .B(n121_adj_227), 
         .Z(n42713)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i57_2_lut_rep_1014.init = 16'h6666;
    L6MUX21 i25151 (.D0(n40407), .D1(n40408), .SD(n9902), .Z(n40411));
    LUT4 div_4016_LessThan_3206_i55_4_lut (.A(n4755), .B(n105), .C(n22245), 
         .D(n4783), .Z(n55_adj_787)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i55_4_lut.init = 16'h663c;
    L6MUX21 i25152 (.D0(n40409), .D1(n40410), .SD(n9902), .Z(n40412));
    LUT4 i25931_4_lut (.A(n42701), .B(n42703), .C(n42702), .D(n37793), 
         .Z(n37808)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25931_4_lut.init = 16'hfffe;
    LUT4 i22514_4_lut (.A(n42707), .B(n42708), .C(n42709), .D(n37761), 
         .Z(n37774)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22514_4_lut.init = 16'h1011;
    LUT4 i22501_4_lut (.A(n42710), .B(n43_adj_332), .C(n41), .D(n37752), 
         .Z(n37761)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22501_4_lut.init = 16'h1011;
    LUT4 i25067_3_lut (.A(\U[6] [14]), .B(\U[7] [14]), .C(i[0]), .Z(n40327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25067_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i52_3_lut_3_lut (.A(n2714), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n52_adj_322)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i22469_4_lut (.A(n42713), .B(n42714), .C(n42715), .D(n37714), 
         .Z(n37729)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22469_4_lut.init = 16'h0100;
    L6MUX21 i25166 (.D0(n40422), .D1(n40423), .SD(n9902), .Z(n40426));
    LUT4 i25066_3_lut (.A(\U[4] [14]), .B(\U[5] [14]), .C(i[0]), .Z(n40326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25066_3_lut.init = 16'hcaca;
    LUT4 i25278_3_lut (.A(\U[8] [28]), .B(\U[9] [28]), .C(i[0]), .Z(n40538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25278_3_lut.init = 16'hcaca;
    L6MUX21 i25167 (.D0(n40424), .D1(n40425), .SD(n9902), .Z(n40427));
    LUT4 i22454_4_lut (.A(n42716), .B(n42717), .C(n42719), .D(n37701), 
         .Z(n37714)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22454_4_lut.init = 16'h5455;
    LUT4 i22441_4_lut (.A(n42718), .B(n43), .C(n42720), .D(n39), .Z(n37701)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22441_4_lut.init = 16'h5554;
    LUT4 i22836_2_lut_3_lut_4_lut (.A(n3440), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3439), .Z(n38096)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22836_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i25065_3_lut (.A(\U[2] [14]), .B(\U[3] [14]), .C(i[0]), .Z(n40325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25065_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i39_2_lut (.A(n2723), .B(n130_adj_233), 
         .Z(n39)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i39_2_lut.init = 16'h6666;
    FD1P3IX x_3___i125 (.D(n5497), .SP(clk_c_enable_832), .CD(n30987), 
            .CK(clk_c), .Q(\x[0] [28]));   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(35[10] 137[6])
    defparam x_3___i125.GSR = "ENABLED";
    LUT4 i22410_4_lut (.A(n42724), .B(n42725), .C(n42727), .D(n37657), 
         .Z(n37670)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22410_4_lut.init = 16'h0001;
    LUT4 i22397_4_lut (.A(n42726), .B(n42728), .C(n47_adj_306), .D(n37646), 
         .Z(n37657)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22397_4_lut.init = 16'h0001;
    L6MUX21 i25181 (.D0(n40437), .D1(n40438), .SD(n9902), .Z(n40441));
    L6MUX21 i25182 (.D0(n40439), .D1(n40440), .SD(n9902), .Z(n40442));
    L6MUX21 i25196 (.D0(n40452), .D1(n40453), .SD(n9902), .Z(n40456));
    LUT4 i22386_4_lut (.A(n45_adj_304), .B(n42729), .C(n2569), .D(n130_adj_233), 
         .Z(n37646)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22386_4_lut.init = 16'h1001;
    LUT4 i25064_3_lut (.A(\U[0] [14]), .B(\U[1] [14]), .C(i[0]), .Z(n40324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25064_3_lut.init = 16'hcaca;
    L6MUX21 i25197 (.D0(n40454), .D1(n40455), .SD(n9902), .Z(n40457));
    LUT4 div_4016_LessThan_1761_i55_2_lut_rep_1015 (.A(n2715), .B(n122_adj_228), 
         .Z(n42714)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i55_2_lut_rep_1015.init = 16'h6666;
    L6MUX21 i25211 (.D0(n40467), .D1(n40468), .SD(n9902), .Z(n40471));
    L6MUX21 i25212 (.D0(n40469), .D1(n40470), .SD(n9902), .Z(n40472));
    LUT4 i25277_3_lut (.A(\U[6] [28]), .B(\U[7] [28]), .C(i[0]), .Z(n40537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25277_3_lut.init = 16'hcaca;
    LUT4 i25816_4_lut (.A(n42730), .B(n42731), .C(n42732), .D(n37616), 
         .Z(n37635)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25816_4_lut.init = 16'hfeff;
    LUT4 i22356_4_lut (.A(n42733), .B(n42735), .C(n42734), .D(n37603), 
         .Z(n37616)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22356_4_lut.init = 16'h1011;
    L6MUX21 i25226 (.D0(n40482), .D1(n40483), .SD(n9902), .Z(n40486));
    LUT4 i22343_4_lut (.A(n42736), .B(n49_adj_293), .C(n47), .D(n37594), 
         .Z(n37603)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22343_4_lut.init = 16'h1011;
    LUT4 i25941_4_lut (.A(n42737), .B(n37578), .C(n42738), .D(n37571), 
         .Z(n37586)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25941_4_lut.init = 16'hfbff;
    L6MUX21 i25227 (.D0(n40484), .D1(n40485), .SD(n9902), .Z(n40487));
    LUT4 i23316_4_lut (.A(n42588), .B(n42590), .C(n42591), .D(n38551), 
         .Z(n38576)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23316_4_lut.init = 16'h0100;
    LUT4 i22311_4_lut (.A(n42740), .B(n42739), .C(n42741), .D(n37558), 
         .Z(n37571)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22311_4_lut.init = 16'h5455;
    L6MUX21 i25241 (.D0(n40497), .D1(n40498), .SD(n9902), .Z(n40501));
    L6MUX21 i25242 (.D0(n40499), .D1(n40500), .SD(n9902), .Z(n40502));
    L6MUX21 i25256 (.D0(n40512), .D1(n40513), .SD(n9902), .Z(n40516));
    LUT4 i22473_2_lut_3_lut_4_lut (.A(n2715), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n2714), .Z(n37733)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22473_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i22298_4_lut (.A(n51_adj_282), .B(n42743), .C(n42742), .D(n45), 
         .Z(n37558)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22298_4_lut.init = 16'h5554;
    LUT4 i25056_3_lut (.A(\U[14] [13]), .B(\U[15] [13]), .C(i[0]), .Z(n40316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25056_3_lut.init = 16'hcaca;
    LUT4 i23291_4_lut (.A(n42593), .B(n42592), .C(n42594), .D(n38536), 
         .Z(n38551)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23291_4_lut.init = 16'h0100;
    LUT4 i23276_4_lut (.A(n43_adj_509), .B(n42596), .C(n42595), .D(n38515), 
         .Z(n38536)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23276_4_lut.init = 16'h5455;
    LUT4 i23255_4_lut (.A(n37_adj_505), .B(n42597), .C(n42598), .D(n38502), 
         .Z(n38515)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23255_4_lut.init = 16'h0001;
    LUT4 i24407_4_lut (.A(n42448), .B(n42447), .C(n42449), .D(n39646), 
         .Z(n39667)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24407_4_lut.init = 16'h0100;
    LUT4 i25055_3_lut (.A(\U[12] [13]), .B(\U[13] [13]), .C(i[0]), .Z(n40315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25055_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i53_2_lut_rep_1016 (.A(n2716), .B(n123), 
         .Z(n42715)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i53_2_lut_rep_1016.init = 16'h6666;
    L6MUX21 i25257 (.D0(n40514), .D1(n40515), .SD(n9902), .Z(n40517));
    LUT4 select_5271_Select_15_i5_4_lut (.A(n118_adj_100), .B(i[15]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[15])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_15_i5_4_lut.init = 16'heca0;
    LUT4 select_5271_Select_14_i5_4_lut (.A(n121_adj_150), .B(i[14]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[14])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_14_i5_4_lut.init = 16'heca0;
    LUT4 i23242_4_lut (.A(n31_adj_501), .B(n42600), .C(n42599), .D(n38491), 
         .Z(n38502)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23242_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_1446_i45_2_lut (.A(n2252), .B(n130_adj_233), 
         .Z(n45)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1446_i45_2_lut.init = 16'h6666;
    LUT4 i23231_4_lut (.A(n25_adj_497), .B(n42601), .C(n3974), .D(n130_adj_233), 
         .Z(n38491)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23231_4_lut.init = 16'h1001;
    L6MUX21 i25271 (.D0(n40527), .D1(n40528), .SD(n9902), .Z(n40531));
    LUT4 i25953_4_lut (.A(n42744), .B(n42745), .C(n42747), .D(n37531), 
         .Z(n37544)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25953_4_lut.init = 16'hfffe;
    LUT4 i24386_4_lut (.A(n42450), .B(n42459), .C(n42458), .D(n39566), 
         .Z(n39646)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24386_4_lut.init = 16'h5455;
    L6MUX21 i25272 (.D0(n40529), .D1(n40530), .SD(n9902), .Z(n40532));
    L6MUX21 i25286 (.D0(n40542), .D1(n40543), .SD(n9902), .Z(n40546));
    LUT4 div_4016_LessThan_2841_i64_4_lut (.A(n50_adj_601), .B(n62_adj_607), 
         .C(n42530), .D(n39011), .Z(n64_adj_608)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i64_4_lut.init = 16'hcacc;
    L6MUX21 i25287 (.D0(n40544), .D1(n40545), .SD(n9902), .Z(n40547));
    LUT4 i22271_4_lut (.A(n42746), .B(n42748), .C(n53), .D(n37520), 
         .Z(n37531)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22271_4_lut.init = 16'h0001;
    LUT4 select_5271_Select_13_i5_4_lut (.A(n124_adj_154), .B(i[13]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[13])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_13_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_2246_i43_2_lut_rep_959 (.A(n3441), .B(n123), 
         .Z(n42658)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i43_2_lut_rep_959.init = 16'h6666;
    LUT4 i22260_4_lut (.A(n51), .B(n42749), .C(n2089), .D(n130_adj_233), 
         .Z(n37520)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22260_4_lut.init = 16'h1001;
    LUT4 select_5271_Select_12_i5_4_lut (.A(n127_adj_102), .B(i[12]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[12])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_12_i5_4_lut.init = 16'heca0;
    LUT4 i25054_3_lut (.A(\U[10] [13]), .B(\U[11] [13]), .C(i[0]), .Z(n40314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25054_3_lut.init = 16'hcaca;
    LUT4 i25053_3_lut (.A(\U[8] [13]), .B(\U[9] [13]), .C(i[0]), .Z(n40313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25053_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i50_3_lut_3_lut (.A(n2716), .B(n123), .C(n42_adj_317), 
         .Z(n50_adj_321)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25052_3_lut (.A(\U[6] [13]), .B(\U[7] [13]), .C(i[0]), .Z(n40312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25052_3_lut.init = 16'hcaca;
    L6MUX21 i25301 (.D0(n40557), .D1(n40558), .SD(n9902), .Z(n40561));
    LUT4 i23709_4_lut (.A(n42536), .B(n42539), .C(n42538), .D(n38944), 
         .Z(n38969)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23709_4_lut.init = 16'h0100;
    LUT4 i25276_3_lut (.A(\U[4] [28]), .B(\U[5] [28]), .C(i[0]), .Z(n40536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25276_3_lut.init = 16'hcaca;
    L6MUX21 i25302 (.D0(n40559), .D1(n40560), .SD(n9902), .Z(n40562));
    LUT4 i22464_3_lut_4_lut (.A(n2716), .B(n123), .C(n43), .D(n42716), 
         .Z(n37724)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22464_3_lut_4_lut.init = 16'h0009;
    LUT4 i25051_3_lut (.A(\U[4] [13]), .B(\U[5] [13]), .C(i[0]), .Z(n40311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25051_3_lut.init = 16'hcaca;
    LUT4 i24411_2_lut_3_lut_4_lut (.A(n4757), .B(n108), .C(n109_adj_219), 
         .D(n4758), .Z(n39671)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24411_2_lut_3_lut_4_lut.init = 16'h9009;
    L6MUX21 i25316 (.D0(n40572), .D1(n40573), .SD(n9902), .Z(n40576));
    LUT4 div_4016_LessThan_2841_i54_3_lut_3_lut (.A(n4314), .B(n107_adj_218), 
         .C(n52_adj_602), .Z(n54_adj_603)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2841_i57_2_lut_rep_833 (.A(n4316), .B(n109_adj_219), 
         .Z(n42532)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i57_2_lut_rep_833.init = 16'h6666;
    LUT4 div_4016_LessThan_3137_i44_3_lut_3_lut (.A(n4757), .B(n108), .C(n109_adj_219), 
         .Z(n44_adj_727)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2841_i59_2_lut_rep_834 (.A(n4315), .B(n108), 
         .Z(n42533)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i59_2_lut_rep_834.init = 16'h6666;
    LUT4 i25275_3_lut (.A(\U[2] [28]), .B(\U[3] [28]), .C(i[0]), .Z(n40535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25275_3_lut.init = 16'hcaca;
    LUT4 i23684_4_lut (.A(n42541), .B(n42540), .C(n42542), .D(n38929), 
         .Z(n38944)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23684_4_lut.init = 16'h0100;
    L6MUX21 i25317 (.D0(n40574), .D1(n40575), .SD(n9902), .Z(n40577));
    L6MUX21 i25331 (.D0(n40587), .D1(n40588), .SD(n9902), .Z(n40591));
    L6MUX21 i25332 (.D0(n40589), .D1(n40590), .SD(n9902), .Z(n40592));
    LUT4 i23669_4_lut (.A(n37_adj_594), .B(n42544), .C(n42543), .D(n38908), 
         .Z(n38929)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23669_4_lut.init = 16'h5455;
    LUT4 i25050_3_lut (.A(\U[2] [13]), .B(\U[3] [13]), .C(i[0]), .Z(n40310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25050_3_lut.init = 16'hcaca;
    PFUMX i24862 (.BLUT(n40114), .ALUT(n40115), .C0(i[1]), .Z(n40122));
    LUT4 div_4016_LessThan_2841_i52_3_lut_3_lut (.A(n4315), .B(n108), .C(n109_adj_219), 
         .Z(n52_adj_602)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i52_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25180 (.BLUT(n40435), .ALUT(n40436), .C0(i[1]), .Z(n40440));
    LUT4 i23757_2_lut_3_lut_4_lut (.A(n4315), .B(n108), .C(n109_adj_219), 
         .D(n4316), .Z(n39017)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23757_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i25049_3_lut (.A(\U[0] [13]), .B(\U[1] [13]), .C(i[0]), .Z(n40309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25049_3_lut.init = 16'hcaca;
    PFUMX i24863 (.BLUT(n40116), .ALUT(n40117), .C0(i[1]), .Z(n40123));
    LUT4 div_4016_LessThan_1761_i51_2_lut_rep_1017 (.A(n2717), .B(n124_adj_229), 
         .Z(n42716)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i51_2_lut_rep_1017.init = 16'h6666;
    LUT4 i25274_3_lut (.A(\U[0] [28]), .B(\U[1] [28]), .C(i[0]), .Z(n40534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25274_3_lut.init = 16'hcaca;
    LUT4 i23648_4_lut (.A(n31_adj_590), .B(n42545), .C(n42546), .D(n38895), 
         .Z(n38908)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23648_4_lut.init = 16'h0001;
    PFUMX i24864 (.BLUT(n40118), .ALUT(n40119), .C0(i[1]), .Z(n40124));
    LUT4 div_4016_LessThan_3137_i47_2_lut_rep_750 (.A(n4759), .B(n110_adj_220), 
         .Z(n42449)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i47_2_lut_rep_750.init = 16'h6666;
    LUT4 i25266_3_lut (.A(\U[14] [27]), .B(\U[15] [27]), .C(i[0]), .Z(n40526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25266_3_lut.init = 16'hcaca;
    LUT4 i25676_4_lut_4_lut (.A(n42537), .B(n38975), .C(n44_adj_598), 
         .D(n20_adj_583), .Z(n46_adj_599)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25676_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i23635_4_lut (.A(n25_adj_586), .B(n42548), .C(n42547), .D(n38884), 
         .Z(n38895)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23635_4_lut.init = 16'h0001;
    PFUMX i24865 (.BLUT(n40120), .ALUT(n40121), .C0(i[1]), .Z(n40125));
    LUT4 i25041_3_lut (.A(\U[14] [12]), .B(\U[15] [12]), .C(i[0]), .Z(n40301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25041_3_lut.init = 16'hcaca;
    LUT4 i23730_4_lut_4_lut (.A(n42537), .B(n38969), .C(n42534), .D(n42535), 
         .Z(n38990)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23730_4_lut_4_lut.init = 16'h000b;
    LUT4 div_4016_LessThan_3137_i26_3_lut_3_lut (.A(n4759), .B(n110_adj_220), 
         .C(n18_adj_712), .Z(n26_adj_717)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i26_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i24877 (.BLUT(n40129), .ALUT(n40130), .C0(i[1]), .Z(n40137));
    LUT4 i25040_3_lut (.A(\U[12] [12]), .B(\U[13] [12]), .C(i[0]), .Z(n40300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25040_3_lut.init = 16'hcaca;
    PFUMX i25192 (.BLUT(n40444), .ALUT(n40445), .C0(i[1]), .Z(n40452));
    PFUMX i24878 (.BLUT(n40131), .ALUT(n40132), .C0(i[1]), .Z(n40138));
    LUT4 div_4016_LessThan_2841_i53_2_lut_rep_835 (.A(n4318), .B(n111), 
         .Z(n42534)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i53_2_lut_rep_835.init = 16'h6666;
    LUT4 i23624_4_lut (.A(n19_adj_582), .B(n42549), .C(n4337), .D(n130_adj_233), 
         .Z(n38884)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23624_4_lut.init = 16'h1001;
    LUT4 div_4016_LessThan_1761_i42_3_lut_3_lut (.A(n2717), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n42_adj_317)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25039_3_lut (.A(\U[10] [12]), .B(\U[11] [12]), .C(i[0]), .Z(n40299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25039_3_lut.init = 16'hcaca;
    PFUMX i24879 (.BLUT(n40133), .ALUT(n40134), .C0(i[1]), .Z(n40139));
    LUT4 select_5271_Select_11_i5_4_lut (.A(n130_adj_99), .B(i[11]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[11])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_11_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_1761_i49_2_lut_rep_1018 (.A(n2718), .B(n125_adj_230), 
         .Z(n42717)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i49_2_lut_rep_1018.init = 16'h6666;
    LUT4 div_4016_LessThan_1761_i46_3_lut_3_lut (.A(n2718), .B(n125_adj_230), 
         .C(n44_adj_318), .Z(n46_adj_319)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2246_i40_3_lut_3_lut (.A(n3441), .B(n123), .C(n32_adj_402), 
         .Z(n40_adj_408)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25038_3_lut (.A(\U[8] [12]), .B(\U[9] [12]), .C(i[0]), .Z(n40298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25038_3_lut.init = 16'hcaca;
    LUT4 i23602_4_lut (.A(n42552), .B(n42551), .C(n42554), .D(n38847), 
         .Z(n38862)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23602_4_lut.init = 16'h0100;
    LUT4 select_5271_Select_10_i5_4_lut (.A(n133_adj_90), .B(i[10]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[10])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_10_i5_4_lut.init = 16'heca0;
    LUT4 i23560_4_lut (.A(n42557), .B(n42558), .C(n42560), .D(n38797), 
         .Z(n38820)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23560_4_lut.init = 16'h0100;
    LUT4 i25902_3_lut (.A(n57_adj_789), .B(n55_adj_787), .C(n53_adj_785), 
         .Z(n40053)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25902_3_lut.init = 16'hfefe;
    PFUMX i24880 (.BLUT(n40135), .ALUT(n40136), .C0(i[1]), .Z(n40140));
    LUT4 i25265_3_lut (.A(\U[12] [27]), .B(\U[13] [27]), .C(i[0]), .Z(n40525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25265_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i45_2_lut_rep_1019 (.A(n2720), .B(n127_adj_231), 
         .Z(n42718)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i45_2_lut_rep_1019.init = 16'h6666;
    LUT4 div_4016_LessThan_1761_i47_2_lut_rep_1020 (.A(n2719), .B(n126), 
         .Z(n42719)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i47_2_lut_rep_1020.init = 16'h6666;
    LUT4 select_5271_Select_9_i5_4_lut (.A(n136_adj_53), .B(i[9]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[9])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_9_i5_4_lut.init = 16'heca0;
    LUT4 i22446_2_lut_3_lut_4_lut (.A(n2719), .B(n126), .C(n127_adj_231), 
         .D(n2720), .Z(n37706)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22446_2_lut_3_lut_4_lut.init = 16'h9009;
    PFUMX i24892 (.BLUT(n40144), .ALUT(n40145), .C0(i[1]), .Z(n40152));
    LUT4 i22827_3_lut_4_lut (.A(n3441), .B(n123), .C(n33_adj_403), .D(n42660), 
         .Z(n38087)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22827_3_lut_4_lut.init = 16'h0009;
    PFUMX i25193 (.BLUT(n40446), .ALUT(n40447), .C0(i[1]), .Z(n40453));
    LUT4 i23537_4_lut (.A(n42559), .B(n42561), .C(n39_adj_565), .D(n38782), 
         .Z(n38797)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23537_4_lut.init = 16'h0001;
    LUT4 i23522_4_lut (.A(n42563), .B(n42562), .C(n33_adj_561), .D(n38763), 
         .Z(n38782)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23522_4_lut.init = 16'h0100;
    LUT4 i25037_3_lut (.A(\U[6] [12]), .B(\U[7] [12]), .C(i[0]), .Z(n40297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25037_3_lut.init = 16'hcaca;
    LUT4 i23503_4_lut (.A(n31_adj_559), .B(n42564), .C(n27_adj_556), .D(n38750), 
         .Z(n38763)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23503_4_lut.init = 16'h1011;
    PFUMX i24893 (.BLUT(n40146), .ALUT(n40147), .C0(i[1]), .Z(n40153));
    LUT4 i25264_3_lut (.A(\U[10] [27]), .B(\U[11] [27]), .C(i[0]), .Z(n40524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25264_3_lut.init = 16'hcaca;
    PFUMX i24894 (.BLUT(n40148), .ALUT(n40149), .C0(i[1]), .Z(n40154));
    PFUMX i24895 (.BLUT(n40150), .ALUT(n40151), .C0(i[1]), .Z(n40155));
    LUT4 div_4016_LessThan_1761_i44_3_lut_3_lut (.A(n2719), .B(n126), .C(n127_adj_231), 
         .Z(n44_adj_318)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1761_i41_2_lut_rep_1021 (.A(n2722), .B(n129), 
         .Z(n42720)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i41_2_lut_rep_1021.init = 16'h6666;
    LUT4 i25036_3_lut (.A(\U[4] [12]), .B(\U[5] [12]), .C(i[0]), .Z(n40296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25036_3_lut.init = 16'hcaca;
    LUT4 i25263_3_lut (.A(\U[8] [27]), .B(\U[9] [27]), .C(i[0]), .Z(n40523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25263_3_lut.init = 16'hcaca;
    LUT4 select_5271_Select_8_i5_4_lut (.A(n139_adj_94), .B(i[8]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[8])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_8_i5_4_lut.init = 16'heca0;
    LUT4 i25035_3_lut (.A(\U[2] [12]), .B(\U[3] [12]), .C(i[0]), .Z(n40295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25035_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1761_i40_3_lut_3_lut (.A(n2722), .B(n129), .C(n130_adj_233), 
         .Z(n40_adj_316)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1761_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25034_3_lut (.A(\U[0] [12]), .B(\U[1] [12]), .C(i[0]), .Z(n40294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25034_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i53_4_lut (.A(n4756), .B(n106_adj_217), 
         .C(n22246), .D(n4783), .Z(n53_adj_785)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i53_4_lut.init = 16'h663c;
    PFUMX i24907 (.BLUT(n40159), .ALUT(n40160), .C0(i[1]), .Z(n40167));
    LUT4 div_4016_LessThan_2246_i39_2_lut_rep_960 (.A(n3443), .B(n125_adj_230), 
         .Z(n42659)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i39_2_lut_rep_960.init = 16'h6666;
    PFUMX i25194 (.BLUT(n40448), .ALUT(n40449), .C0(i[1]), .Z(n40454));
    LUT4 i25262_3_lut (.A(\U[6] [27]), .B(\U[7] [27]), .C(i[0]), .Z(n40522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25262_3_lut.init = 16'hcaca;
    LUT4 i23490_4_lut (.A(n42566), .B(n42565), .C(n42567), .D(n38741), 
         .Z(n38750)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23490_4_lut.init = 16'h1011;
    PFUMX i24908 (.BLUT(n40161), .ALUT(n40162), .C0(i[1]), .Z(n40168));
    LUT4 i24306_4_lut (.A(n42460), .B(n21_adj_714), .C(n42461), .D(n11_adj_707), 
         .Z(n39566)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24306_4_lut.init = 16'h5554;
    LUT4 i25261_3_lut (.A(\U[4] [27]), .B(\U[5] [27]), .C(i[0]), .Z(n40521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25261_3_lut.init = 16'hcaca;
    LUT4 i25927_4_lut (.A(n42556), .B(n42555), .C(n42557), .D(n38824), 
         .Z(n38842)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25927_4_lut.init = 16'hfffe;
    PFUMX i24909 (.BLUT(n40163), .ALUT(n40164), .C0(i[1]), .Z(n40169));
    LUT4 i25260_3_lut (.A(\U[2] [27]), .B(\U[3] [27]), .C(i[0]), .Z(n40520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25260_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i26_3_lut_3_lut (.A(n4318), .B(n111), .C(n123), 
         .Z(n26_adj_587)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1658_i63_2_lut_rep_1022 (.A(n2558), .B(n119_adj_226), 
         .Z(n42721)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i63_2_lut_rep_1022.init = 16'h6666;
    LUT4 i25026_3_lut (.A(\U[14] [11]), .B(\U[15] [11]), .C(i[0]), .Z(n40286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25026_3_lut.init = 16'hcaca;
    PFUMX i24910 (.BLUT(n40165), .ALUT(n40166), .C0(i[1]), .Z(n40170));
    PFUMX i24922 (.BLUT(n40174), .ALUT(n40175), .C0(i[1]), .Z(n40182));
    PFUMX i25195 (.BLUT(n40450), .ALUT(n40451), .C0(i[1]), .Z(n40455));
    LUT4 div_4016_LessThan_1658_i50_3_lut_3_lut (.A(n2558), .B(n119_adj_226), 
         .C(n40), .Z(n50_adj_308)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25025_3_lut (.A(\U[12] [11]), .B(\U[13] [11]), .C(i[0]), .Z(n40285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25025_3_lut.init = 16'hcaca;
    PFUMX i24923 (.BLUT(n40176), .ALUT(n40177), .C0(i[1]), .Z(n40183));
    LUT4 div_4016_LessThan_2841_i55_2_lut_rep_836 (.A(n4317), .B(n110_adj_220), 
         .Z(n42535)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i55_2_lut_rep_836.init = 16'h6666;
    LUT4 select_5271_Select_7_i5_4_lut (.A(n142_adj_96), .B(i[7]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[7])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_7_i5_4_lut.init = 16'heca0;
    LUT4 select_5271_Select_6_i5_4_lut (.A(n145_adj_103), .B(i[6]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[6])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_6_i5_4_lut.init = 16'heca0;
    PFUMX i24924 (.BLUT(n40178), .ALUT(n40179), .C0(i[1]), .Z(n40184));
    LUT4 i25024_3_lut (.A(\U[10] [11]), .B(\U[11] [11]), .C(i[0]), .Z(n40284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25024_3_lut.init = 16'hcaca;
    LUT4 i25579_4_lut_4_lut (.A(n42722), .B(n37681), .C(n56_adj_311), 
         .D(n42_adj_302), .Z(n58_adj_312)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25579_4_lut_4_lut.init = 16'hf4b0;
    PFUMX i24925 (.BLUT(n40180), .ALUT(n40181), .C0(i[1]), .Z(n40185));
    PFUMX i25207 (.BLUT(n40459), .ALUT(n40460), .C0(i[1]), .Z(n40467));
    LUT4 div_4016_LessThan_2841_i34_3_lut_3_lut (.A(n4317), .B(n110_adj_220), 
         .C(n26_adj_587), .Z(n34_adj_592)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25259_3_lut (.A(\U[0] [27]), .B(\U[1] [27]), .C(i[0]), .Z(n40519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25259_3_lut.init = 16'hcaca;
    LUT4 i25958_4_lut_4_lut (.A(n42722), .B(n37670), .C(n42723), .D(n42721), 
         .Z(n37691)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25958_4_lut_4_lut.init = 16'hff04;
    LUT4 div_4016_LessThan_2993_i64_4_lut (.A(n46_adj_661), .B(n62_adj_669), 
         .C(n42488), .D(n39340), .Z(n64_adj_670)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i64_4_lut.init = 16'hcacc;
    LUT4 i22874_2_lut_3_lut_4_lut (.A(n3443), .B(n125_adj_230), .C(n116_adj_224), 
         .D(n3434), .Z(n38134)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22874_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i25023_3_lut (.A(\U[8] [11]), .B(\U[9] [11]), .C(i[0]), .Z(n40283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25023_3_lut.init = 16'hcaca;
    PFUMX i24937 (.BLUT(n40189), .ALUT(n40190), .C0(i[1]), .Z(n40197));
    LUT4 div_4016_LessThan_2841_i49_2_lut_rep_837 (.A(n4320), .B(n113_adj_222), 
         .Z(n42536)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i49_2_lut_rep_837.init = 16'h6666;
    PFUMX i24938 (.BLUT(n40191), .ALUT(n40192), .C0(i[1]), .Z(n40198));
    LUT4 i24051_4_lut (.A(n42491), .B(n42490), .C(n42492), .D(n39296), 
         .Z(n39311)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24051_4_lut.init = 16'h0100;
    LUT4 i25251_3_lut (.A(\U[14] [26]), .B(\U[15] [26]), .C(i[0]), .Z(n40511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25251_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1658_i61_2_lut_rep_1023 (.A(n2559), .B(n120), 
         .Z(n42722)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i61_2_lut_rep_1023.init = 16'h6666;
    PFUMX i24939 (.BLUT(n40193), .ALUT(n40194), .C0(i[1]), .Z(n40199));
    LUT4 i25022_3_lut (.A(\U[6] [11]), .B(\U[7] [11]), .C(i[0]), .Z(n40282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25022_3_lut.init = 16'hcaca;
    LUT4 i25021_3_lut (.A(\U[4] [11]), .B(\U[5] [11]), .C(i[0]), .Z(n40281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25021_3_lut.init = 16'hcaca;
    PFUMX i25208 (.BLUT(n40461), .ALUT(n40462), .C0(i[1]), .Z(n40468));
    PFUMX i24940 (.BLUT(n40195), .ALUT(n40196), .C0(i[1]), .Z(n40200));
    LUT4 i24009_4_lut (.A(n42496), .B(n42497), .C(n42499), .D(n39246), 
         .Z(n39269)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24009_4_lut.init = 16'h0100;
    LUT4 i25250_3_lut (.A(\U[12] [26]), .B(\U[13] [26]), .C(i[0]), .Z(n40510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25250_3_lut.init = 16'hcaca;
    LUT4 i23986_4_lut (.A(n42498), .B(n42500), .C(n33_adj_654), .D(n39231), 
         .Z(n39246)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23986_4_lut.init = 16'h0001;
    L6MUX21 div_4016_LessThan_2058_i64 (.D0(n52_adj_372), .D1(n62_adj_377), 
            .SD(n37961), .Z(n64_adj_378));
    LUT4 i25249_3_lut (.A(\U[10] [26]), .B(\U[11] [26]), .C(i[0]), .Z(n40509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25249_3_lut.init = 16'hcaca;
    LUT4 i25248_3_lut (.A(\U[8] [26]), .B(\U[9] [26]), .C(i[0]), .Z(n40508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25248_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_3_i7_3_lut (.A(n5350), .B(n27_adj_187), .C(n5325), 
         .Z(n888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i7_3_lut.init = 16'hcaca;
    LUT4 i23971_4_lut (.A(n42502), .B(n42501), .C(n42503), .D(n39212), 
         .Z(n39231)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23971_4_lut.init = 16'h0100;
    LUT4 i23952_4_lut (.A(n42504), .B(n42505), .C(n21_adj_647), .D(n39199), 
         .Z(n39212)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23952_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_1658_i56_3_lut_3_lut (.A(n2559), .B(n120), .C(n54_adj_310), 
         .Z(n56_adj_311)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i56_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i24952 (.BLUT(n40204), .ALUT(n40205), .C0(i[1]), .Z(n40212));
    LUT4 i25020_3_lut (.A(\U[2] [11]), .B(\U[3] [11]), .C(i[0]), .Z(n40280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25020_3_lut.init = 16'hcaca;
    LUT4 select_5271_Select_5_i5_4_lut (.A(n148_adj_113), .B(i[5]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_5_i5_4_lut.init = 16'heca0;
    PFUMX i24953 (.BLUT(n40206), .ALUT(n40207), .C0(i[1]), .Z(n40213));
    PFUMX i25209 (.BLUT(n40463), .ALUT(n40464), .C0(i[1]), .Z(n40469));
    LUT4 i25019_3_lut (.A(\U[0] [11]), .B(\U[1] [11]), .C(i[0]), .Z(n40279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25019_3_lut.init = 16'hcaca;
    PFUMX i24954 (.BLUT(n40208), .ALUT(n40209), .C0(i[1]), .Z(n40214));
    LUT4 div_4016_LessThan_1658_i59_2_lut_rep_1024 (.A(n2560), .B(n121_adj_227), 
         .Z(n42723)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i59_2_lut_rep_1024.init = 16'h6666;
    LUT4 i25247_3_lut (.A(\U[6] [26]), .B(\U[7] [26]), .C(i[0]), .Z(n40507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25247_3_lut.init = 16'hcaca;
    PFUMX i24955 (.BLUT(n40210), .ALUT(n40211), .C0(i[1]), .Z(n40215));
    LUT4 i25011_3_lut (.A(\U[14] [10]), .B(\U[15] [10]), .C(i[0]), .Z(n40271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25011_3_lut.init = 16'hcaca;
    LUT4 i25246_3_lut (.A(\U[4] [26]), .B(\U[5] [26]), .C(i[0]), .Z(n40506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25246_3_lut.init = 16'hcaca;
    PFUMX i24967 (.BLUT(n40219), .ALUT(n40220), .C0(i[1]), .Z(n40227));
    LUT4 i23939_4_lut (.A(n42507), .B(n42506), .C(n42508), .D(n39190), 
         .Z(n39199)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23939_4_lut.init = 16'h1011;
    L6MUX21 div_4016_LessThan_1961_i64 (.D0(n54_adj_355), .D1(n62_adj_359), 
            .SD(n37879), .Z(n64_adj_360));
    LUT4 i25010_3_lut (.A(\U[12] [10]), .B(\U[13] [10]), .C(i[0]), .Z(n40270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25010_3_lut.init = 16'hcaca;
    LUT4 i25009_3_lut (.A(\U[10] [10]), .B(\U[11] [10]), .C(i[0]), .Z(n40269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25009_3_lut.init = 16'hcaca;
    LUT4 select_5271_Select_4_i5_4_lut (.A(n151_adj_159), .B(i[4]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[4])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_4_i5_4_lut.init = 16'heca0;
    LUT4 div_4016_LessThan_2246_i41_2_lut_rep_961 (.A(n3442), .B(n124_adj_229), 
         .Z(n42660)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i41_2_lut_rep_961.init = 16'h6666;
    LUT4 i25008_3_lut (.A(\U[8] [10]), .B(\U[9] [10]), .C(i[0]), .Z(n40268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25008_3_lut.init = 16'hcaca;
    LUT4 i25007_3_lut (.A(\U[6] [10]), .B(\U[7] [10]), .C(i[0]), .Z(n40267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25007_3_lut.init = 16'hcaca;
    PFUMX i24968 (.BLUT(n40221), .ALUT(n40222), .C0(i[1]), .Z(n40228));
    LUT4 div_4016_LessThan_2841_i42_3_lut_3_lut (.A(n4320), .B(n113_adj_222), 
         .C(n114), .Z(n42_adj_597)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i42_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 div_4016_LessThan_1862_i64 (.D0(n56_adj_339), .D1(n62_adj_342), 
            .SD(n37808), .Z(n64_adj_343));
    LUT4 div_4016_LessThan_2918_i64_4_lut (.A(n48_adj_632), .B(n62_adj_639), 
         .C(n42509), .D(n39171), .Z(n64_adj_640)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i64_4_lut.init = 16'hcacc;
    PFUMX i25210 (.BLUT(n40465), .ALUT(n40466), .C0(i[1]), .Z(n40470));
    LUT4 i25245_3_lut (.A(\U[2] [26]), .B(\U[3] [26]), .C(i[0]), .Z(n40505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25245_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2993_i10_4_lut (.A(n132), .B(n131_adj_234), .C(n4565), 
         .D(n891), .Z(n10_adj_641)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i10_4_lut.init = 16'h0c8e;
    LUT4 i23886_4_lut (.A(n42512), .B(n42514), .C(n42515), .D(n39129), 
         .Z(n39146)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23886_4_lut.init = 16'h0001;
    LUT4 i24400_3_lut_4_lut (.A(n4759), .B(n110_adj_220), .C(n21_adj_714), 
         .D(n42450), .Z(n39660)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24400_3_lut_4_lut.init = 16'h0009;
    PFUMX i24969 (.BLUT(n40223), .ALUT(n40224), .C0(i[1]), .Z(n40229));
    LUT4 div_4016_LessThan_2841_i51_2_lut_rep_838 (.A(n4319), .B(n112_adj_221), 
         .Z(n42537)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i51_2_lut_rep_838.init = 16'h6666;
    PFUMX i24970 (.BLUT(n40225), .ALUT(n40226), .C0(i[1]), .Z(n40230));
    LUT4 i25244_3_lut (.A(\U[0] [26]), .B(\U[1] [26]), .C(i[0]), .Z(n40504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25244_3_lut.init = 16'hcaca;
    PFUMX i24982 (.BLUT(n40234), .ALUT(n40235), .C0(i[1]), .Z(n40242));
    LUT4 i25006_3_lut (.A(\U[4] [10]), .B(\U[5] [10]), .C(i[0]), .Z(n40266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25006_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i45_2_lut_rep_751 (.A(n4760), .B(n111), 
         .Z(n42450)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i45_2_lut_rep_751.init = 16'h6666;
    LUT4 select_5271_Select_3_i5_4_lut (.A(n154_adj_158), .B(i[3]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_3_i5_4_lut.init = 16'heca0;
    PFUMX i24983 (.BLUT(n40236), .ALUT(n40237), .C0(i[1]), .Z(n40243));
    LUT4 i25236_3_lut (.A(\U[14] [25]), .B(\U[15] [25]), .C(i[0]), .Z(n40496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25236_3_lut.init = 16'hcaca;
    PFUMX i24984 (.BLUT(n40238), .ALUT(n40239), .C0(i[1]), .Z(n40244));
    LUT4 div_4016_LessThan_2841_i44_3_lut_3_lut (.A(n4319), .B(n112_adj_221), 
         .C(n42_adj_597), .Z(n44_adj_598)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25005_3_lut (.A(\U[2] [10]), .B(\U[3] [10]), .C(i[0]), .Z(n40265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25005_3_lut.init = 16'hcaca;
    PFUMX i25222 (.BLUT(n40474), .ALUT(n40475), .C0(i[1]), .Z(n40482));
    PFUMX i24985 (.BLUT(n40240), .ALUT(n40241), .C0(i[1]), .Z(n40245));
    LUT4 i25004_3_lut (.A(\U[0] [10]), .B(\U[1] [10]), .C(i[0]), .Z(n40264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25004_3_lut.init = 16'hcaca;
    LUT4 i25235_3_lut (.A(\U[12] [25]), .B(\U[13] [25]), .C(i[0]), .Z(n40495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25235_3_lut.init = 16'hcaca;
    PFUMX i25223 (.BLUT(n40476), .ALUT(n40477), .C0(i[1]), .Z(n40483));
    PFUMX i24997 (.BLUT(n40249), .ALUT(n40250), .C0(i[1]), .Z(n40257));
    PFUMX i25224 (.BLUT(n40478), .ALUT(n40479), .C0(i[1]), .Z(n40484));
    LUT4 div_4016_LessThan_2841_i45_2_lut_rep_839 (.A(n4322), .B(n115_adj_223), 
         .Z(n42538)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i45_2_lut_rep_839.init = 16'h6666;
    PFUMX i24998 (.BLUT(n40251), .ALUT(n40252), .C0(i[1]), .Z(n40258));
    PFUMX i25225 (.BLUT(n40480), .ALUT(n40481), .C0(i[1]), .Z(n40485));
    PFUMX i24999 (.BLUT(n40253), .ALUT(n40254), .C0(i[1]), .Z(n40259));
    LUT4 i24996_3_lut (.A(\U[14] [9]), .B(\U[15] [9]), .C(i[0]), .Z(n40256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24996_3_lut.init = 16'hcaca;
    PFUMX i25237 (.BLUT(n40489), .ALUT(n40490), .C0(i[1]), .Z(n40497));
    PFUMX i25238 (.BLUT(n40491), .ALUT(n40492), .C0(i[1]), .Z(n40498));
    LUT4 i23844_4_lut (.A(n42518), .B(n42521), .C(n42520), .D(n39083), 
         .Z(n39104)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23844_4_lut.init = 16'h0100;
    PFUMX i25239 (.BLUT(n40493), .ALUT(n40494), .C0(i[1]), .Z(n40499));
    LUT4 select_5271_Select_2_i5_4_lut (.A(n157_adj_157), .B(i[2]), .C(done_N_1932), 
         .D(n13381), .Z(i_31__N_1607[2])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam select_5271_Select_2_i5_4_lut.init = 16'heca0;
    PFUMX i25000 (.BLUT(n40255), .ALUT(n40256), .C0(i[1]), .Z(n40260));
    LUT4 div_4016_LessThan_3137_i18_3_lut_3_lut (.A(n4760), .B(n111), .C(n123), 
         .Z(n18_adj_712)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23823_4_lut (.A(n42522), .B(n35_adj_625), .C(n42524), .D(n39066), 
         .Z(n39083)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23823_4_lut.init = 16'h1011;
    PFUMX i25240 (.BLUT(n40495), .ALUT(n40496), .C0(i[1]), .Z(n40500));
    PFUMX i25012 (.BLUT(n40264), .ALUT(n40265), .C0(i[1]), .Z(n40272));
    LUT4 i23806_4_lut (.A(n42523), .B(n29_adj_621), .C(n42525), .D(n39051), 
         .Z(n39066)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23806_4_lut.init = 16'h0100;
    LUT4 i23791_4_lut (.A(n42526), .B(n23_adj_617), .C(n42528), .D(n39038), 
         .Z(n39051)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23791_4_lut.init = 16'h5455;
    LUT4 div_4016_LessThan_2246_i32_3_lut_3_lut (.A(n3442), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n32_adj_402)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i32_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25252 (.BLUT(n40504), .ALUT(n40505), .C0(i[1]), .Z(n40512));
    PFUMX i25013 (.BLUT(n40266), .ALUT(n40267), .C0(i[1]), .Z(n40273));
    LUT4 i24995_3_lut (.A(\U[12] [9]), .B(\U[13] [9]), .C(i[0]), .Z(n40255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24995_3_lut.init = 16'hcaca;
    PFUMX i25014 (.BLUT(n40268), .ALUT(n40269), .C0(i[1]), .Z(n40274));
    PFUMX i25253 (.BLUT(n40506), .ALUT(n40507), .C0(i[1]), .Z(n40513));
    LUT4 i25234_3_lut (.A(\U[10] [25]), .B(\U[11] [25]), .C(i[0]), .Z(n40494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25234_3_lut.init = 16'hcaca;
    PFUMX i25015 (.BLUT(n40270), .ALUT(n40271), .C0(i[1]), .Z(n40275));
    LUT4 i25233_3_lut (.A(\U[8] [25]), .B(\U[9] [25]), .C(i[0]), .Z(n40493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25233_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i40_3_lut_3_lut (.A(n4322), .B(n115_adj_223), 
         .C(n22_adj_584), .Z(n40_adj_596)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23704_3_lut_4_lut (.A(n4322), .B(n115_adj_223), .C(n25_adj_586), 
         .D(n42541), .Z(n38964)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23704_3_lut_4_lut.init = 16'h0009;
    PFUMX i25027 (.BLUT(n40279), .ALUT(n40280), .C0(i[1]), .Z(n40287));
    LUT4 i25232_3_lut (.A(\U[6] [25]), .B(\U[7] [25]), .C(i[0]), .Z(n40492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25232_3_lut.init = 16'hcaca;
    LUT4 i23778_4_lut (.A(n42527), .B(n17_adj_613), .C(n42529), .D(n13_adj_610), 
         .Z(n39038)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23778_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_2918_i13_2_lut (.A(n4452), .B(n130_adj_233), 
         .Z(n13_adj_610)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i13_2_lut.init = 16'h6666;
    PFUMX i25254 (.BLUT(n40508), .ALUT(n40509), .C0(i[1]), .Z(n40514));
    LUT4 div_4016_LessThan_2246_i37_2_lut_rep_962 (.A(n3444), .B(n126), 
         .Z(n42661)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i37_2_lut_rep_962.init = 16'h6666;
    LUT4 div_4016_LessThan_2841_i47_2_lut_rep_840 (.A(n4321), .B(n114), 
         .Z(n42539)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i47_2_lut_rep_840.init = 16'h6666;
    PFUMX i25028 (.BLUT(n40281), .ALUT(n40282), .C0(i[1]), .Z(n40288));
    PFUMX i25255 (.BLUT(n40510), .ALUT(n40511), .C0(i[1]), .Z(n40515));
    LUT4 i25231_3_lut (.A(\U[4] [25]), .B(\U[5] [25]), .C(i[0]), .Z(n40491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25231_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2246_i34_3_lut_3_lut (.A(n3444), .B(n126), .C(n127_adj_231), 
         .Z(n34_adj_404)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i34_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25267 (.BLUT(n40519), .ALUT(n40520), .C0(i[1]), .Z(n40527));
    PFUMX i25029 (.BLUT(n40283), .ALUT(n40284), .C0(i[1]), .Z(n40289));
    LUT4 i23715_2_lut_3_lut_4_lut (.A(n4321), .B(n114), .C(n113_adj_222), 
         .D(n4320), .Z(n38975)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23715_2_lut_3_lut_4_lut.init = 16'h9009;
    L6MUX21 div_4016_LessThan_1761_i64 (.D0(n58_adj_325), .D1(n62_adj_327), 
            .SD(n37746), .Z(n64_adj_328));
    LUT4 i25230_3_lut (.A(\U[2] [25]), .B(\U[3] [25]), .C(i[0]), .Z(n40490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25230_3_lut.init = 16'hcaca;
    LUT4 i25229_3_lut (.A(\U[0] [25]), .B(\U[1] [25]), .C(i[0]), .Z(n40489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25229_3_lut.init = 16'hcaca;
    PFUMX i25030 (.BLUT(n40285), .ALUT(n40286), .C0(i[1]), .Z(n40290));
    LUT4 i24994_3_lut (.A(\U[10] [9]), .B(\U[11] [9]), .C(i[0]), .Z(n40254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24994_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1658_i54_3_lut_3_lut (.A(n2560), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n54_adj_310)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2993_i18_3_lut_3_lut (.A(n4550), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n18_adj_645)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3066_i64_4_lut (.A(n44_adj_693), .B(n62_adj_702), 
         .C(n42464), .D(n39514), .Z(n64_adj_703)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i64_4_lut.init = 16'hcacc;
    PFUMX i25042 (.BLUT(n40294), .ALUT(n40295), .C0(i[1]), .Z(n40302));
    PFUMX i25268 (.BLUT(n40521), .ALUT(n40522), .C0(i[1]), .Z(n40528));
    LUT4 i22798_3_lut_4_lut (.A(n3447), .B(n129), .C(n130_adj_233), .D(n3448), 
         .Z(n38058)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22798_3_lut_4_lut.init = 16'h9009;
    PFUMX i25269 (.BLUT(n40523), .ALUT(n40524), .C0(i[1]), .Z(n40529));
    LUT4 i24993_3_lut (.A(\U[8] [9]), .B(\U[9] [9]), .C(i[0]), .Z(n40253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24993_3_lut.init = 16'hcaca;
    LUT4 i25221_3_lut (.A(\U[14] [24]), .B(\U[15] [24]), .C(i[0]), .Z(n40481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25221_3_lut.init = 16'hcaca;
    PFUMX i25043 (.BLUT(n40296), .ALUT(n40297), .C0(i[1]), .Z(n40303));
    LUT4 div_4016_LessThan_1658_i57_2_lut_rep_1025 (.A(n2561), .B(n122_adj_228), 
         .Z(n42724)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i57_2_lut_rep_1025.init = 16'h6666;
    LUT4 i24185_4_lut (.A(n42473), .B(n42475), .C(n42476), .D(n39420), 
         .Z(n39445)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24185_4_lut.init = 16'h0100;
    LUT4 i24773_4_lut_4_lut (.A(n42439), .B(n40007), .C(n53_adj_785), 
         .D(n55_adj_787), .Z(n40033)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24773_4_lut_4_lut.init = 16'h0004;
    LUT4 i24992_3_lut (.A(\U[6] [9]), .B(\U[7] [9]), .C(i[0]), .Z(n40252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24992_3_lut.init = 16'hcaca;
    PFUMX i25044 (.BLUT(n40298), .ALUT(n40299), .C0(i[1]), .Z(n40304));
    LUT4 i24160_4_lut (.A(n42478), .B(n42477), .C(n42479), .D(n39405), 
         .Z(n39420)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24160_4_lut.init = 16'h0100;
    PFUMX i25270 (.BLUT(n40525), .ALUT(n40526), .C0(i[1]), .Z(n40530));
    LUT4 i25220_3_lut (.A(\U[12] [24]), .B(\U[13] [24]), .C(i[0]), .Z(n40480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25220_3_lut.init = 16'hcaca;
    LUT4 i24991_3_lut (.A(\U[4] [9]), .B(\U[5] [9]), .C(i[0]), .Z(n40251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24991_3_lut.init = 16'hcaca;
    LUT4 i25219_3_lut (.A(\U[10] [24]), .B(\U[11] [24]), .C(i[0]), .Z(n40479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25219_3_lut.init = 16'hcaca;
    LUT4 i25921_4_lut (.A(n42438), .B(n39_adj_773), .C(n37_adj_771), .D(n39975), 
         .Z(n39991)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25921_4_lut.init = 16'hfffe;
    PFUMX i25045 (.BLUT(n40300), .ALUT(n40301), .C0(i[1]), .Z(n40305));
    PFUMX i25057 (.BLUT(n40309), .ALUT(n40310), .C0(i[1]), .Z(n40317));
    LUT4 i24715_3_lut (.A(n35_adj_769), .B(n33_adj_767), .C(n15_adj_749), 
         .Z(n39975)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24715_3_lut.init = 16'h0101;
    PFUMX i25282 (.BLUT(n40534), .ALUT(n40535), .C0(i[1]), .Z(n40542));
    LUT4 i22421_2_lut_3_lut_4_lut (.A(n2561), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n2560), .Z(n37681)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22421_2_lut_3_lut_4_lut.init = 16'h9009;
    PFUMX i25058 (.BLUT(n40311), .ALUT(n40312), .C0(i[1]), .Z(n40318));
    LUT4 i25218_3_lut (.A(\U[8] [24]), .B(\U[9] [24]), .C(i[0]), .Z(n40478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25218_3_lut.init = 16'hcaca;
    L6MUX21 div_4016_LessThan_1658_i64 (.D0(n60_adj_313), .D1(n62_adj_314), 
            .SD(n37691), .Z(n64_adj_315));
    LUT4 i24145_4_lut (.A(n31_adj_686), .B(n42481), .C(n42480), .D(n39384), 
         .Z(n39405)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24145_4_lut.init = 16'h5455;
    PFUMX i25283 (.BLUT(n40536), .ALUT(n40537), .C0(i[1]), .Z(n40543));
    LUT4 div_4016_LessThan_2993_i35_2_lut_rep_801 (.A(n4552), .B(n118_adj_225), 
         .Z(n42500)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i35_2_lut_rep_801.init = 16'h6666;
    LUT4 div_4016_LessThan_1658_i55_2_lut_rep_1026 (.A(n2562), .B(n123), 
         .Z(n42725)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i55_2_lut_rep_1026.init = 16'h6666;
    PFUMX i25059 (.BLUT(n40313), .ALUT(n40314), .C0(i[1]), .Z(n40319));
    LUT4 div_4016_LessThan_1658_i52_3_lut_3_lut (.A(n2562), .B(n123), .C(n44_adj_303), 
         .Z(n52_adj_309)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i52_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25060 (.BLUT(n40315), .ALUT(n40316), .C0(i[1]), .Z(n40320));
    LUT4 i24990_3_lut (.A(\U[2] [9]), .B(\U[3] [9]), .C(i[0]), .Z(n40250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24990_3_lut.init = 16'hcaca;
    PFUMX i25072 (.BLUT(n40324), .ALUT(n40325), .C0(i[1]), .Z(n40332));
    LUT4 i25722_4_lut_4_lut (.A(n42452), .B(n39629), .C(n36_adj_723), 
         .D(n12_adj_708), .Z(n38_adj_724)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25722_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_4016_LessThan_2993_i20_3_lut_3_lut (.A(n4552), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n20_adj_646)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24989_3_lut (.A(\U[0] [9]), .B(\U[1] [9]), .C(i[0]), .Z(n40249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24989_3_lut.init = 16'hcaca;
    LUT4 i25217_3_lut (.A(\U[6] [24]), .B(\U[7] [24]), .C(i[0]), .Z(n40477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25217_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i41_2_lut_rep_841 (.A(n4324), .B(n117), 
         .Z(n42540)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i41_2_lut_rep_841.init = 16'h6666;
    LUT4 i24124_4_lut (.A(n25_adj_682), .B(n42482), .C(n42483), .D(n39371), 
         .Z(n39384)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24124_4_lut.init = 16'h0001;
    PFUMX i25284 (.BLUT(n40538), .ALUT(n40539), .C0(i[1]), .Z(n40544));
    LUT4 i24111_4_lut (.A(n19_adj_678), .B(n42485), .C(n42484), .D(n39360), 
         .Z(n39371)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24111_4_lut.init = 16'h0001;
    PFUMX i25073 (.BLUT(n40326), .ALUT(n40327), .C0(i[1]), .Z(n40333));
    LUT4 i24100_4_lut (.A(n13_adj_674), .B(n42486), .C(n4673), .D(n130_adj_233), 
         .Z(n39360)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24100_4_lut.init = 16'h1001;
    LUT4 div_4016_LessThan_2246_i30_3_lut_3_lut (.A(n3447), .B(n129), .C(n130_adj_233), 
         .Z(n30_adj_401)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2246_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25216_3_lut (.A(\U[4] [24]), .B(\U[5] [24]), .C(i[0]), .Z(n40476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25216_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2153_i63_2_lut_rep_963 (.A(n3293), .B(n114), 
         .Z(n42662)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i63_2_lut_rep_963.init = 16'h6666;
    LUT4 div_4016_LessThan_2153_i58_3_lut_3_lut (.A(n3293), .B(n114), .C(n36_adj_383), 
         .Z(n58_adj_396)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2993_i29_2_lut_rep_802 (.A(n4555), .B(n121_adj_227), 
         .Z(n42501)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i29_2_lut_rep_802.init = 16'h6666;
    LUT4 i22412_3_lut_4_lut (.A(n2562), .B(n123), .C(n45_adj_304), .D(n42727), 
         .Z(n37672)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22412_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2153_i61_2_lut_rep_964 (.A(n3294), .B(n115_adj_223), 
         .Z(n42663)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i61_2_lut_rep_964.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i24_3_lut_3_lut (.A(n4555), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n24_adj_649)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i24_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25074 (.BLUT(n40328), .ALUT(n40329), .C0(i[1]), .Z(n40334));
    LUT4 div_4016_LessThan_2153_i56_3_lut_3_lut (.A(n3294), .B(n115_adj_223), 
         .C(n38_adj_385), .Z(n56_adj_395)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2153_i57_2_lut_rep_965 (.A(n3296), .B(n117), 
         .Z(n42664)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i57_2_lut_rep_965.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i31_2_lut_rep_803 (.A(n4554), .B(n120), 
         .Z(n42502)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i31_2_lut_rep_803.init = 16'h6666;
    LUT4 div_4016_LessThan_2153_i52_3_lut_3_lut (.A(n3296), .B(n117), .C(n40_adj_386), 
         .Z(n52_adj_392)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i52_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3206_i62_4_lut (.A(n40_adj_774), .B(n60_adj_792), 
         .C(n61_adj_793), .D(n39888), .Z(n62_adj_794)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i62_4_lut.init = 16'hcacc;
    LUT4 i25874_4_lut (.A(n42550), .B(n42552), .C(n42551), .D(n38857), 
         .Z(n40108)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25874_4_lut.init = 16'hfeff;
    LUT4 div_4016_LessThan_3206_i60_3_lut (.A(n48_adj_781), .B(n58_adj_790), 
         .C(n40059), .Z(n60_adj_792)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i60_3_lut.init = 16'hacac;
    LUT4 i24628_4_lut (.A(n59_adj_791), .B(n57_adj_789), .C(n55_adj_787), 
         .D(n39861), .Z(n39888)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24628_4_lut.init = 16'h0100;
    LUT4 i23597_4_lut (.A(n42554), .B(n42553), .C(n42563), .D(n38777), 
         .Z(n38857)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23597_4_lut.init = 16'h1011;
    PFUMX i25285 (.BLUT(n40540), .ALUT(n40541), .C0(i[1]), .Z(n40545));
    PFUMX i25075 (.BLUT(n40330), .ALUT(n40331), .C0(i[1]), .Z(n40335));
    LUT4 i24981_3_lut (.A(\U[14] [8]), .B(\U[15] [8]), .C(i[0]), .Z(n40241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24981_3_lut.init = 16'hcaca;
    LUT4 i23517_4_lut (.A(n42562), .B(n33_adj_561), .C(n31_adj_559), .D(n38765), 
         .Z(n38777)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23517_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_3206_i58_3_lut (.A(n52_adj_784), .B(n56_adj_788), 
         .C(n40061), .Z(n58_adj_790)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i58_3_lut.init = 16'hacac;
    LUT4 i25820_4_lut (.A(n42635), .B(n42636), .C(n42638), .D(n38230), 
         .Z(n38255)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25820_4_lut.init = 16'hfeff;
    LUT4 div_4016_LessThan_3206_i56_3_lut (.A(n54_adj_786), .B(n102), .C(n61_adj_793), 
         .Z(n56_adj_788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i56_3_lut.init = 16'hcaca;
    LUT4 i24576_4_lut (.A(n47_adj_780), .B(n45_adj_778), .C(n43_adj_776), 
         .D(n39987), .Z(n39836)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24576_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_2993_i26_3_lut_3_lut (.A(n4554), .B(n120), .C(n24_adj_649), 
         .Z(n26_adj_650)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i26_3_lut_3_lut.init = 16'hd4d4;
    L6MUX21 div_4016_LessThan_1553_i64 (.D0(n52_adj_295), .D1(n62_adj_300), 
            .SD(n37635), .Z(n64_adj_301));
    LUT4 i25866_3_lut_4_lut (.A(n3296), .B(n117), .C(n53_adj_393), .D(n42666), 
         .Z(n38036)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25866_3_lut_4_lut.init = 16'hfff6;
    PFUMX i25087 (.BLUT(n40339), .ALUT(n40340), .C0(i[1]), .Z(n40347));
    LUT4 div_4016_LessThan_3206_i59_4_lut (.A(n4753), .B(n103_adj_215), 
         .C(n22243), .D(n4783), .Z(n59_adj_791)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i59_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2153_i59_2_lut_rep_966 (.A(n3295), .B(n116_adj_224), 
         .Z(n42665)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i59_2_lut_rep_966.init = 16'h6666;
    LUT4 i24436_4_lut (.A(n42444), .B(n42446), .C(n42459), .D(n39573), 
         .Z(n39696)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24436_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_3137_i41_2_lut_rep_752 (.A(n4762), .B(n113_adj_222), 
         .Z(n42451)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i41_2_lut_rep_752.init = 16'h6666;
    LUT4 i24534_4_lut (.A(n35_adj_769), .B(n33_adj_767), .C(n31_adj_765), 
         .D(n39773), .Z(n39794)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24534_4_lut.init = 16'h0100;
    LUT4 i22970_4_lut (.A(n42637), .B(n42640), .C(n42639), .D(n38214), 
         .Z(n38230)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22970_4_lut.init = 16'h1011;
    LUT4 i25215_3_lut (.A(\U[2] [24]), .B(\U[3] [24]), .C(i[0]), .Z(n40475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25215_3_lut.init = 16'hcaca;
    LUT4 i24513_4_lut (.A(n29_adj_763), .B(n27_adj_761), .C(n25_adj_759), 
         .D(n39756), .Z(n39773)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24513_4_lut.init = 16'h1011;
    PFUMX i25088 (.BLUT(n40341), .ALUT(n40342), .C0(i[1]), .Z(n40348));
    LUT4 i24496_4_lut (.A(n23_adj_757), .B(n21_adj_755), .C(n19_adj_753), 
         .D(n39741), .Z(n39756)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24496_4_lut.init = 16'h0100;
    LUT4 div_4016_LessThan_2153_i38_3_lut_3_lut (.A(n3295), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n38_adj_385)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i38_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24481_4_lut (.A(n17_adj_751), .B(n15_adj_749), .C(n13_adj_747), 
         .D(n39728), .Z(n39741)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24481_4_lut.init = 16'h5455;
    LUT4 i25607_4_lut_4_lut (.A(n42667), .B(n38007), .C(n46_adj_389), 
         .D(n32_adj_381), .Z(n48_adj_390)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25607_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i24468_4_lut (.A(n11_adj_745), .B(n9_adj_743), .C(n7_adj_741), 
         .D(n5_adj_739), .Z(n39728)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24468_4_lut.init = 16'h5554;
    LUT4 div_4016_LessThan_3206_i5_4_lut (.A(n4780), .B(n130_adj_233), .C(n22270), 
         .D(n4783), .Z(n5_adj_739)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i5_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2993_i27_2_lut_rep_804 (.A(n4556), .B(n122_adj_228), 
         .Z(n42503)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i27_2_lut_rep_804.init = 16'h6666;
    LUT4 i25214_3_lut (.A(\U[0] [24]), .B(\U[1] [24]), .C(i[0]), .Z(n40474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25214_3_lut.init = 16'hcaca;
    LUT4 i24980_3_lut (.A(\U[12] [8]), .B(\U[13] [8]), .C(i[0]), .Z(n40240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24980_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1658_i51_2_lut_rep_1027 (.A(n2564), .B(n125_adj_230), 
         .Z(n42726)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i51_2_lut_rep_1027.init = 16'h6666;
    LUT4 div_4016_LessThan_2153_i55_2_lut_rep_967 (.A(n3297), .B(n118_adj_225), 
         .Z(n42666)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i55_2_lut_rep_967.init = 16'h6666;
    PFUMX i25297 (.BLUT(n40549), .ALUT(n40550), .C0(i[1]), .Z(n40557));
    LUT4 i24979_3_lut (.A(\U[10] [8]), .B(\U[11] [8]), .C(i[0]), .Z(n40239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24979_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2153_i40_3_lut_3_lut (.A(n3297), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n40_adj_386)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23968_2_lut_3_lut_4_lut (.A(n4556), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n4555), .Z(n39228)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23968_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_3206_i9_4_lut (.A(n4778), .B(n128_adj_232), .C(n22268), 
         .D(n4783), .Z(n9_adj_743)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i9_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2762_i33_2_lut (.A(n4211), .B(n122_adj_228), 
         .Z(n33_adj_561)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i33_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i25_2_lut_rep_805 (.A(n4557), .B(n123), 
         .Z(n42504)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i25_2_lut_rep_805.init = 16'h6666;
    PFUMX i25089 (.BLUT(n40343), .ALUT(n40344), .C0(i[1]), .Z(n40349));
    LUT4 i22954_4_lut (.A(n42641), .B(n49_adj_436), .C(n37_adj_429), .D(n38167), 
         .Z(n38214)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22954_4_lut.init = 16'h1011;
    LUT4 i24048_2_lut_3_lut_4_lut (.A(n4557), .B(n123), .C(n111), .D(n4545), 
         .Z(n39308)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24048_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2762_i31_2_lut (.A(n4212), .B(n123), .Z(n31_adj_559)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2762_i31_2_lut.init = 16'h6666;
    LUT4 div_4016_LessThan_2993_i23_2_lut_rep_806 (.A(n4558), .B(n124_adj_229), 
         .Z(n42505)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i23_2_lut_rep_806.init = 16'h6666;
    LUT4 div_4016_LessThan_1658_i48_3_lut_3_lut (.A(n2564), .B(n125_adj_230), 
         .C(n46_adj_305), .Z(n48_adj_307)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i48_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25298 (.BLUT(n40551), .ALUT(n40552), .C0(i[1]), .Z(n40558));
    LUT4 div_4016_LessThan_2993_i14_3_lut_3_lut (.A(n4558), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n14_adj_643)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i14_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2153_i51_2_lut_rep_968 (.A(n3299), .B(n120), 
         .Z(n42667)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i51_2_lut_rep_968.init = 16'h6666;
    LUT4 i24801_4_lut (.A(n61_adj_793), .B(n59_adj_791), .C(n57_adj_789), 
         .D(n40043), .Z(n40061)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24801_4_lut.init = 16'h1011;
    LUT4 i24783_4_lut (.A(n55_adj_787), .B(n53_adj_785), .C(n25_adj_759), 
         .D(n39760), .Z(n40043)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24783_4_lut.init = 16'h1011;
    LUT4 i24500_2_lut (.A(n23_adj_757), .B(n21_adj_755), .Z(n39760)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24500_2_lut.init = 16'h1111;
    PFUMX i25299 (.BLUT(n40553), .ALUT(n40554), .C0(i[1]), .Z(n40559));
    LUT4 div_4016_LessThan_2841_i36_3_lut_3_lut (.A(n4324), .B(n117), .C(n24_adj_585), 
         .Z(n36_adj_593)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3206_i21_4_lut (.A(n4772), .B(n122_adj_228), 
         .C(n22262), .D(n4783), .Z(n21_adj_755)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i21_4_lut.init = 16'h663c;
    LUT4 i25206_3_lut (.A(\U[14] [23]), .B(\U[15] [23]), .C(i[0]), .Z(n40466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25206_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2153_i46_3_lut_3_lut (.A(n3299), .B(n120), .C(n44_adj_388), 
         .Z(n46_adj_389)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3066_i8_4_lut (.A(n132), .B(n131_adj_234), .C(n4674), 
         .D(n892), .Z(n8_adj_671)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3066_i8_4_lut.init = 16'h0c8e;
    LUT4 div_4016_LessThan_2153_i49_2_lut_rep_969 (.A(n3300), .B(n121_adj_227), 
         .Z(n42668)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i49_2_lut_rep_969.init = 16'h6666;
    LUT4 mux_4010_i30_4_lut (.A(n76), .B(n36704), .C(n15805), .D(i[1]), 
         .Z(n5327)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i30_4_lut.init = 16'hca0a;
    LUT4 i24978_3_lut (.A(\U[8] [8]), .B(\U[9] [8]), .C(i[0]), .Z(n40238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24978_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_111 (.A(i[0]), .B(\y[3] [29]), .Z(n36704)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_111.init = 16'h8888;
    LUT4 mux_4010_i31_4_lut (.A(n73), .B(n36702), .C(n15805), .D(i[1]), 
         .Z(n5326)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i31_4_lut.init = 16'hca0a;
    PFUMX i25090 (.BLUT(n40345), .ALUT(n40346), .C0(i[1]), .Z(n40350));
    LUT4 div_4016_LessThan_2993_i17_2_lut_rep_807 (.A(n4561), .B(n127_adj_231), 
         .Z(n42506)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i17_2_lut_rep_807.init = 16'h6666;
    LUT4 i25205_3_lut (.A(\U[12] [23]), .B(\U[13] [23]), .C(i[0]), .Z(n40465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25205_3_lut.init = 16'hcaca;
    LUT4 i24601_4_lut_4_lut (.A(n42439), .B(n39836), .C(n49_adj_782), 
         .D(n53_adj_785), .Z(n39861)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24601_4_lut_4_lut.init = 16'h0004;
    LUT4 i24799_4_lut (.A(n61_adj_793), .B(n59_adj_791), .C(n57_adj_789), 
         .D(n40035), .Z(n40059)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24799_4_lut.init = 16'h0100;
    LUT4 div_4016_LessThan_2153_i44_3_lut_3_lut (.A(n3300), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n44_adj_388)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_112 (.A(i[0]), .B(\y[3] [30]), .Z(n36702)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_112.init = 16'h8888;
    LUT4 i24757_4_lut (.A(n49_adj_782), .B(n47_adj_780), .C(n45_adj_778), 
         .D(n39999), .Z(n40017)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24757_4_lut.init = 16'h0100;
    LUT4 i24739_4_lut (.A(n43_adj_776), .B(n25_adj_759), .C(n23_adj_757), 
         .D(n39753), .Z(n39999)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24739_4_lut.init = 16'h5455;
    LUT4 div_4016_LessThan_2153_i45_2_lut_rep_970 (.A(n3302), .B(n123), 
         .Z(n42669)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i45_2_lut_rep_970.init = 16'h6666;
    LUT4 mux_4010_i28_4_lut (.A(n82), .B(n36696), .C(n15805), .D(i[1]), 
         .Z(n5329)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i28_4_lut.init = 16'hca0a;
    LUT4 i24977_3_lut (.A(\U[6] [8]), .B(\U[7] [8]), .C(i[0]), .Z(n40237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24977_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_113 (.A(i[0]), .B(\y[3] [27]), .Z(n36696)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_113.init = 16'h8888;
    LUT4 i24493_4_lut (.A(n21_adj_755), .B(n19_adj_753), .C(n17_adj_751), 
         .D(n9_adj_743), .Z(n39753)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24493_4_lut.init = 16'h5554;
    LUT4 mux_4010_i29_4_lut (.A(n79), .B(n36698), .C(n15805), .D(i[1]), 
         .Z(n5328)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i29_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_114 (.A(i[0]), .B(\y[3] [28]), .Z(n36698)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_114.init = 16'h8888;
    LUT4 i22738_3_lut_4_lut (.A(n3302), .B(n123), .C(n35), .D(n42672), 
         .Z(n37998)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22738_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2153_i47_2_lut_rep_971 (.A(n3301), .B(n122_adj_228), 
         .Z(n42670)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i47_2_lut_rep_971.init = 16'h6666;
    LUT4 i22747_2_lut_3_lut_4_lut (.A(n3301), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3300), .Z(n38007)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22747_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i1_2_lut_adj_115 (.A(i[0]), .B(\y[3] [25]), .Z(n36694)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_115.init = 16'h8888;
    LUT4 i24976_3_lut (.A(\U[4] [8]), .B(\U[5] [8]), .C(i[0]), .Z(n40236)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24976_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2153_i42_3_lut_3_lut (.A(n3302), .B(n123), .C(n34_adj_382), 
         .Z(n42_adj_387)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i42_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25102 (.BLUT(n40354), .ALUT(n40355), .C0(i[1]), .Z(n40362));
    LUT4 div_4016_LessThan_2993_i19_2_lut_rep_808 (.A(n4560), .B(n126), 
         .Z(n42507)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i19_2_lut_rep_808.init = 16'h6666;
    LUT4 i25857_4_lut (.A(n42662), .B(n42663), .C(n42665), .D(n42671), 
         .Z(n38054)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25857_4_lut.init = 16'haaab;
    LUT4 div_4016_LessThan_2153_i41_2_lut_rep_972 (.A(n3304), .B(n125_adj_230), 
         .Z(n42671)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i41_2_lut_rep_972.init = 16'h6666;
    PFUMX i25300 (.BLUT(n40555), .ALUT(n40556), .C0(i[1]), .Z(n40560));
    LUT4 div_4016_i3072_1_lut (.A(n104_adj_216), .Z(n4683)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3072_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_1658_i53_2_lut_rep_1028 (.A(n2563), .B(n124_adj_229), 
         .Z(n42727)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i53_2_lut_rep_1028.init = 16'h6666;
    LUT4 i25912_3_lut_4_lut (.A(n4324), .B(n117), .C(n37_adj_594), .D(n42542), 
         .Z(n38948)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25912_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_LessThan_2841_i43_2_lut_rep_842 (.A(n4323), .B(n116_adj_224), 
         .Z(n42541)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i43_2_lut_rep_842.init = 16'h6666;
    LUT4 i23930_3_lut_4_lut (.A(n4563), .B(n129), .C(n130_adj_233), .D(n4564), 
         .Z(n39190)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23930_3_lut_4_lut.init = 16'h9009;
    LUT4 i25859_4_lut (.A(n42662), .B(n42663), .C(n42665), .D(n38034), 
         .Z(n38050)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25859_4_lut.init = 16'hfffe;
    LUT4 div_4016_i3071_1_lut (.A(n103_adj_215), .Z(n4682)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3071_1_lut.init = 16'h5555;
    LUT4 i22725_3_lut_4_lut (.A(n3304), .B(n125_adj_230), .C(n37_adj_384), 
         .D(n42673), .Z(n37985)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22725_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2841_i22_3_lut_3_lut (.A(n4323), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n22_adj_584)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i22_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i23941_2_lut_3_lut_4_lut (.A(n4560), .B(n126), .C(n127_adj_231), 
         .D(n4561), .Z(n39201)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23941_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_i2849_1_lut (.A(n106_adj_217), .Z(n4352)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2849_1_lut.init = 16'h5555;
    PFUMX i25103 (.BLUT(n40356), .ALUT(n40357), .C0(i[1]), .Z(n40363));
    LUT4 div_4016_LessThan_1658_i44_3_lut_3_lut (.A(n2563), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n44_adj_303)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24975_3_lut (.A(\U[2] [8]), .B(\U[3] [8]), .C(i[0]), .Z(n40235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24975_3_lut.init = 16'hcaca;
    PFUMX i25104 (.BLUT(n40358), .ALUT(n40359), .C0(i[1]), .Z(n40364));
    LUT4 div_4016_i2925_1_lut (.A(n105), .Z(n4465)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2925_1_lut.init = 16'h5555;
    LUT4 i24974_3_lut (.A(\U[0] [8]), .B(\U[1] [8]), .C(i[0]), .Z(n40234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24974_3_lut.init = 16'hcaca;
    LUT4 i22774_4_lut (.A(n42664), .B(n42666), .C(n53_adj_393), .D(n37985), 
         .Z(n38034)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22774_4_lut.init = 16'h0001;
    LUT4 div_4016_LessThan_1658_i49_2_lut_rep_1029 (.A(n2565), .B(n126), 
         .Z(n42728)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i49_2_lut_rep_1029.init = 16'h6666;
    LUT4 div_4016_LessThan_2153_i43_2_lut_rep_973 (.A(n3303), .B(n124_adj_229), 
         .Z(n42672)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i43_2_lut_rep_973.init = 16'h6666;
    LUT4 mux_4010_i27_4_lut (.A(n85), .B(n36692), .C(n15805), .D(i[1]), 
         .Z(n5330)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i27_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_2153_i34_3_lut_3_lut (.A(n3303), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n34_adj_382)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i34_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_116 (.A(i[0]), .B(\y[3] [26]), .Z(n36692)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_116.init = 16'h8888;
    LUT4 div_4016_LessThan_3137_i34_3_lut_3_lut (.A(n4762), .B(n113_adj_222), 
         .C(n114), .Z(n34_adj_722)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i34_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25105 (.BLUT(n40360), .ALUT(n40361), .C0(i[1]), .Z(n40365));
    LUT4 mux_4010_i24_4_lut (.A(n94), .B(n36690), .C(n15805), .D(i[1]), 
         .Z(n5333)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i24_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_2841_i39_2_lut_rep_843 (.A(n4325), .B(n118_adj_225), 
         .Z(n42542)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i39_2_lut_rep_843.init = 16'h6666;
    LUT4 i24966_3_lut (.A(\U[14] [7]), .B(\U[15] [7]), .C(i[0]), .Z(n40226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24966_3_lut.init = 16'hcaca;
    LUT4 i25868_4_lut (.A(n42667), .B(n42668), .C(n42670), .D(n37998), 
         .Z(n38012)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25868_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_117 (.A(i[0]), .B(\y[3] [23]), .Z(n36690)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_117.init = 16'h8888;
    LUT4 i25880_4_lut (.A(n42568), .B(n38723), .C(n42569), .D(n38721), 
         .Z(n40102)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25880_4_lut.init = 16'hfbff;
    LUT4 i25818_4_lut (.A(n42635), .B(n42636), .C(n42638), .D(n38239), 
         .Z(n38257)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25818_4_lut.init = 16'hfffe;
    LUT4 div_4016_i2772_1_lut (.A(n108), .Z(n4117)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2772_1_lut.init = 16'h5555;
    LUT4 i23461_4_lut (.A(n42570), .B(n42579), .C(n42578), .D(n38641), 
         .Z(n38721)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23461_4_lut.init = 16'h5455;
    LUT4 i24965_3_lut (.A(\U[12] [7]), .B(\U[13] [7]), .C(i[0]), .Z(n40225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24965_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1658_i46_3_lut_3_lut (.A(n2565), .B(n126), .C(n127_adj_231), 
         .Z(n46_adj_305)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1658_i43_2_lut_rep_1030 (.A(n2568), .B(n129), 
         .Z(n42729)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i43_2_lut_rep_1030.init = 16'h6666;
    LUT4 div_4016_i2850_1_lut (.A(n107_adj_218), .Z(n4236)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2850_1_lut.init = 16'h5555;
    PFUMX i25117 (.BLUT(n40369), .ALUT(n40370), .C0(i[1]), .Z(n40377));
    LUT4 div_4016_i2525_1_lut (.A(n110_adj_220), .Z(n3870)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2525_1_lut.init = 16'h5555;
    LUT4 div_4016_i2609_1_lut (.A(n109_adj_219), .Z(n3995)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2609_1_lut.init = 16'h5555;
    LUT4 i24964_3_lut (.A(\U[10] [7]), .B(\U[11] [7]), .C(i[0]), .Z(n40224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24964_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2153_i39_2_lut_rep_974 (.A(n3305), .B(n126), 
         .Z(n42673)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i39_2_lut_rep_974.init = 16'h6666;
    LUT4 div_4016_i2351_1_lut (.A(n112_adj_221), .Z(n3611)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2351_1_lut.init = 16'h5555;
    PFUMX i25312 (.BLUT(n40564), .ALUT(n40565), .C0(i[1]), .Z(n40572));
    LUT4 div_4016_i2439_1_lut (.A(n111), .Z(n3871)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2439_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_2841_i24_3_lut_3_lut (.A(n4325), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n24_adj_585)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i24_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i2262_1_lut (.A(n114), .Z(n3340)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2262_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_2153_i36_3_lut_3_lut (.A(n3305), .B(n126), .C(n127_adj_231), 
         .Z(n36_adj_383)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i36_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25118 (.BLUT(n40371), .ALUT(n40372), .C0(i[1]), .Z(n40378));
    LUT4 div_4016_LessThan_2841_i33_2_lut_rep_844 (.A(n4328), .B(n121_adj_227), 
         .Z(n42543)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i33_2_lut_rep_844.init = 16'h6666;
    LUT4 mux_4010_i25_4_lut (.A(n91), .B(n36688), .C(n15805), .D(i[1]), 
         .Z(n5332)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i25_4_lut.init = 16'hca0a;
    PFUMX i25119 (.BLUT(n40373), .ALUT(n40374), .C0(i[1]), .Z(n40379));
    LUT4 div_4016_i2352_1_lut (.A(n113_adj_222), .Z(n3477)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2352_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_2153_i33_2_lut_rep_975 (.A(n3308), .B(n129), 
         .Z(n42674)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i33_2_lut_rep_975.init = 16'h6666;
    LUT4 div_4016_i2076_1_lut (.A(n116_adj_224), .Z(n3057)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2076_1_lut.init = 16'h5555;
    LUT4 div_4016_i2170_1_lut (.A(n115_adj_223), .Z(n3479)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i2170_1_lut.init = 16'h5555;
    LUT4 i24963_3_lut (.A(\U[8] [7]), .B(\U[9] [7]), .C(i[0]), .Z(n40223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24963_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i28_3_lut_3_lut (.A(n4328), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n28_adj_588)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i28_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_118 (.A(i[0]), .B(\y[3] [24]), .Z(n36688)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_118.init = 16'h8888;
    LUT4 div_4016_i1781_1_lut (.A(n118_adj_225), .Z(n2762)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1781_1_lut.init = 16'h5555;
    LUT4 mux_4010_i22_4_lut (.A(n100), .B(n36686), .C(n15805), .D(i[1]), 
         .Z(n5335)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i22_4_lut.init = 16'hca0a;
    LUT4 div_4016_i1881_1_lut (.A(n117), .Z(n2911)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1881_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_119 (.A(i[0]), .B(\y[3] [21]), .Z(n36686)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_119.init = 16'h8888;
    LUT4 div_4016_LessThan_1658_i42_3_lut_3_lut (.A(n2568), .B(n129), .C(n130_adj_233), 
         .Z(n42_adj_302)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1658_i42_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i1575_1_lut (.A(n120), .Z(n2455)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1575_1_lut.init = 16'h5555;
    LUT4 mux_4010_i23_4_lut (.A(n97), .B(n36684), .C(n15805), .D(i[1]), 
         .Z(n5334)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i23_4_lut.init = 16'hca0a;
    LUT4 i23381_4_lut (.A(n35_adj_533), .B(n42580), .C(n42581), .D(n23_adj_525), 
         .Z(n38641)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23381_4_lut.init = 16'h5554;
    PFUMX i25120 (.BLUT(n40375), .ALUT(n40376), .C0(i[1]), .Z(n40380));
    LUT4 i25575_4_lut_4_lut (.A(n42730), .B(n37632), .C(n58_adj_298), 
         .D(n44_adj_290), .Z(n60_adj_299)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25575_4_lut_4_lut.init = 16'hf4b0;
    PFUMX i25313 (.BLUT(n40566), .ALUT(n40567), .C0(i[1]), .Z(n40573));
    LUT4 i25917_3_lut_4_lut (.A(n4328), .B(n121_adj_227), .C(n31_adj_590), 
         .D(n42544), .Z(n38926)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25917_3_lut_4_lut.init = 16'hfff6;
    LUT4 div_4016_mux_3_i12_3_lut (.A(n5345), .B(n22_adj_182), .C(n5325), 
         .Z(n883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 div_4016_i1679_1_lut (.A(n119_adj_226), .Z(n3060)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1679_1_lut.init = 16'h5555;
    LUT4 i24962_3_lut (.A(\U[6] [7]), .B(\U[7] [7]), .C(i[0]), .Z(n40222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24962_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2153_i32_3_lut_3_lut (.A(n3308), .B(n129), .C(n130_adj_233), 
         .Z(n32_adj_381)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2153_i32_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1553_i63_2_lut_rep_1031 (.A(n2402), .B(n120), 
         .Z(n42730)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i63_2_lut_rep_1031.init = 16'h6666;
    L6MUX21 div_4016_LessThan_1446_i64 (.D0(n54_adj_284), .D1(n62_adj_288), 
            .SD(n37586), .Z(n64_adj_289));
    LUT4 div_4016_i1361_1_lut (.A(n122_adj_228), .Z(n2298)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1361_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_120 (.A(i[0]), .B(\y[3] [22]), .Z(n36684)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_120.init = 16'h8888;
    LUT4 div_4016_i1469_1_lut (.A(n121_adj_227), .Z(n2456)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1469_1_lut.init = 16'h5555;
    LUT4 div_4016_i1139_1_lut (.A(n124_adj_229), .Z(n1805)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1139_1_lut.init = 16'h5555;
    LUT4 i24961_3_lut (.A(\U[4] [7]), .B(\U[5] [7]), .C(i[0]), .Z(n40221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24961_3_lut.init = 16'hcaca;
    LUT4 div_4016_i1251_1_lut (.A(n123), .Z(n2137)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1251_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_2058_i63_2_lut_rep_976 (.A(n3152), .B(n115_adj_223), 
         .Z(n42675)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i63_2_lut_rep_976.init = 16'h6666;
    LUT4 div_4016_i1026_1_lut (.A(n126), .Z(n1462)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1026_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_1553_i58_3_lut_3_lut (.A(n2402), .B(n120), .C(n56_adj_297), 
         .Z(n58_adj_298)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i58_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24761_2_lut (.A(n49_adj_782), .B(n47_adj_780), .Z(n40021)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24761_2_lut.init = 16'h1111;
    LUT4 div_4016_LessThan_1553_i61_2_lut_rep_1032 (.A(n2403), .B(n121_adj_227), 
         .Z(n42731)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i61_2_lut_rep_1032.init = 16'h6666;
    PFUMX i25132 (.BLUT(n40384), .ALUT(n40385), .C0(i[1]), .Z(n40392));
    LUT4 div_4016_i1140_1_lut (.A(n125_adj_230), .Z(n1635)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i1140_1_lut.init = 16'h5555;
    LUT4 div_4016_i911_1_lut (.A(n128_adj_232), .Z(n2142)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i911_1_lut.init = 16'h5555;
    LUT4 i25204_3_lut (.A(\U[10] [23]), .B(\U[11] [23]), .C(i[0]), .Z(n40464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25204_3_lut.init = 16'hcaca;
    LUT4 div_4016_i910_1_lut (.A(n127_adj_231), .Z(n2141)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i910_1_lut.init = 16'h5555;
    LUT4 div_4016_LessThan_2993_i12_3_lut_3_lut (.A(n4563), .B(n129), .C(n130_adj_233), 
         .Z(n12_adj_642)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24960_3_lut (.A(\U[2] [7]), .B(\U[3] [7]), .C(i[0]), .Z(n40220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24960_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i49_4_lut (.A(n4758), .B(n108), .C(n22248), 
         .D(n4783), .Z(n49_adj_782)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i49_4_lut.init = 16'h663c;
    LUT4 mux_4010_i20_4_lut (.A(n106), .B(n36680), .C(n15805), .D(i[1]), 
         .Z(n5337)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i20_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_121 (.A(i[0]), .B(\y[3] [19]), .Z(n36680)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_121.init = 16'h8888;
    LUT4 div_4016_LessThan_2058_i60_3_lut_3_lut (.A(n3152), .B(n115_adj_223), 
         .C(n58_adj_375), .Z(n60_adj_376)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_4010_i21_4_lut (.A(n103), .B(n36682), .C(n15805), .D(i[1]), 
         .Z(n5336)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i21_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_3137_i6_4_lut (.A(n132), .B(n131_adj_234), .C(n4780), 
         .D(n893), .Z(n6_adj_704)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i6_4_lut.init = 16'h0c8e;
    LUT4 i25604_4_lut_4_lut (.A(n42677), .B(n37949), .C(n54_adj_373), 
         .D(n32_adj_361), .Z(n56_adj_374)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25604_4_lut_4_lut.init = 16'hf4b0;
    PFUMX i25133 (.BLUT(n40386), .ALUT(n40387), .C0(i[1]), .Z(n40393));
    LUT4 div_4016_LessThan_3206_i47_4_lut (.A(n4759), .B(n109_adj_219), 
         .C(n22249), .D(n4783), .Z(n47_adj_780)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i47_4_lut.init = 16'h663c;
    LUT4 i1_2_lut_adj_122 (.A(i[0]), .B(\y[3] [20]), .Z(n36682)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_122.init = 16'h8888;
    LUT4 i24959_3_lut (.A(\U[0] [7]), .B(\U[1] [7]), .C(i[0]), .Z(n40219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24959_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i24_3_lut (.A(n5468), .B(n76_adj_199), .C(n5460), 
         .Z(n109_adj_219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i24_3_lut.init = 16'hcaca;
    LUT4 i25897_4_lut_4_lut (.A(n42677), .B(n37947), .C(n42676), .D(n42675), 
         .Z(n37963)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25897_4_lut_4_lut.init = 16'hfff4;
    PFUMX i25134 (.BLUT(n40388), .ALUT(n40389), .C0(i[1]), .Z(n40394));
    PFUMX i25314 (.BLUT(n40568), .ALUT(n40569), .C0(i[1]), .Z(n40574));
    LUT4 div_4016_LessThan_2993_i15_2_lut_rep_809 (.A(n4562), .B(n128_adj_232), 
         .Z(n42508)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2993_i15_2_lut_rep_809.init = 16'h6666;
    LUT4 i25899_4_lut_4_lut (.A(n42677), .B(n37940), .C(n42676), .D(n42675), 
         .Z(n37961)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25899_4_lut_4_lut.init = 16'hfffb;
    LUT4 mux_4010_i18_4_lut (.A(n112), .B(n36676), .C(n15805), .D(i[1]), 
         .Z(n5339)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i18_4_lut.init = 16'hca0a;
    PFUMX i25135 (.BLUT(n40390), .ALUT(n40391), .C0(i[1]), .Z(n40395));
    LUT4 i25203_3_lut (.A(\U[8] [23]), .B(\U[9] [23]), .C(i[0]), .Z(n40463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25203_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i35_2_lut_rep_845 (.A(n4327), .B(n120), 
         .Z(n42544)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i35_2_lut_rep_845.init = 16'h6666;
    LUT4 div_4016_LessThan_1553_i56_3_lut_3_lut (.A(n2403), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n56_adj_297)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i56_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_123 (.A(i[0]), .B(\y[3] [17]), .Z(n36676)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_123.init = 16'h8888;
    LUT4 i24951_3_lut (.A(\U[14] [6]), .B(\U[15] [6]), .C(i[0]), .Z(n40211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24951_3_lut.init = 16'hcaca;
    LUT4 mux_4010_i19_4_lut (.A(n109), .B(n36678), .C(n15805), .D(i[1]), 
         .Z(n5338)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i19_4_lut.init = 16'hca0a;
    LUT4 i22687_4_lut (.A(n42679), .B(n42678), .C(n42685), .D(n37900), 
         .Z(n37947)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22687_4_lut.init = 16'h1011;
    LUT4 div_4016_LessThan_3137_i43_2_lut_rep_753 (.A(n4761), .B(n112_adj_221), 
         .Z(n42452)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i43_2_lut_rep_753.init = 16'h6666;
    LUT4 i23954_2_lut_3_lut_4_lut (.A(n4562), .B(n128_adj_232), .C(n124_adj_229), 
         .D(n4558), .Z(n39214)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23954_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2058_i61_2_lut_rep_977 (.A(n3153), .B(n116_adj_224), 
         .Z(n42676)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i61_2_lut_rep_977.init = 16'h6666;
    LUT4 div_4016_LessThan_2841_i30_3_lut_3_lut (.A(n4327), .B(n120), .C(n28_adj_588), 
         .Z(n30_adj_589)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2058_i40_3_lut_3_lut (.A(n3153), .B(n116_adj_224), 
         .C(n125_adj_230), .Z(n40_adj_366)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i40_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2918_i63_2_lut_rep_810 (.A(n4427), .B(n105), 
         .Z(n42509)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i63_2_lut_rep_810.init = 16'h6666;
    LUT4 i1_2_lut_adj_124 (.A(i[0]), .B(\y[3] [18]), .Z(n36678)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_124.init = 16'h8888;
    LUT4 mux_4010_i16_4_lut (.A(n118), .B(n36674), .C(n15805), .D(i[1]), 
         .Z(n5341)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i16_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_2058_i59_2_lut_rep_978 (.A(n3154), .B(n117), 
         .Z(n42677)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i59_2_lut_rep_978.init = 16'h6666;
    LUT4 div_4016_mux_3_i15_3_lut (.A(n5342), .B(n19_adj_179), .C(n5325), 
         .Z(n880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_125 (.A(i[0]), .B(\y[3] [15]), .Z(n36674)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_125.init = 16'h8888;
    LUT4 mux_4010_i17_4_lut (.A(n115), .B(n36672), .C(n15805), .D(i[1]), 
         .Z(n5340)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i17_4_lut.init = 16'hca0a;
    PFUMX i25147 (.BLUT(n40399), .ALUT(n40400), .C0(i[1]), .Z(n40407));
    LUT4 div_4016_LessThan_3206_i18_3_lut (.A(n122_adj_228), .B(n121_adj_227), 
         .C(n23_adj_757), .Z(n18_adj_752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i18_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_126 (.A(i[0]), .B(\y[3] [16]), .Z(n36672)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_126.init = 16'h8888;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 div_4016_LessThan_2918_i60_3_lut_3_lut (.A(n4427), .B(n105), .C(n58_adj_637), 
         .Z(n60_adj_638)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i60_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i25923_4_lut (.A(n42438), .B(n39_adj_773), .C(n37_adj_771), .D(n39796), 
         .Z(n39989)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25923_4_lut.init = 16'hfeff;
    LUT4 i24536_4_lut (.A(n35_adj_769), .B(n33_adj_767), .C(n31_adj_765), 
         .D(n39780), .Z(n39796)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24536_4_lut.init = 16'h1011;
    VLO i1 (.Z(GND_net));
    LUT4 mux_4010_i14_4_lut (.A(n124), .B(n36670), .C(n15805), .D(i[1]), 
         .Z(n5343)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i14_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_2058_i54_3_lut_3_lut (.A(n3154), .B(n117), .C(n42_adj_367), 
         .Z(n54_adj_373)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24520_4_lut (.A(n29_adj_763), .B(n27_adj_761), .C(n15_adj_749), 
         .D(n39733), .Z(n39780)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24520_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_adj_127 (.A(i[0]), .B(\y[3] [13]), .Z(n36670)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_127.init = 16'h8888;
    LUT4 mux_4010_i15_4_lut (.A(n121), .B(n36668), .C(n15805), .D(i[1]), 
         .Z(n5342)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i15_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_128 (.A(i[0]), .B(\y[3] [14]), .Z(n36668)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_128.init = 16'h8888;
    LUT4 i25691_4_lut_4_lut (.A(n42511), .B(n39168), .C(n52_adj_634), 
         .D(n16_adj_612), .Z(n54_adj_635)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25691_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i24950_3_lut (.A(\U[12] [6]), .B(\U[13] [6]), .C(i[0]), .Z(n40210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24950_3_lut.init = 16'hcaca;
    PFUMX i25315 (.BLUT(n40570), .ALUT(n40571), .C0(i[1]), .Z(n40575));
    LUT4 i25833_4_lut (.A(n42643), .B(n42642), .C(n42645), .D(n38185), 
         .Z(n38199)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25833_4_lut.init = 16'hfffe;
    LUT4 div_4016_LessThan_2681_i61_2_lut (.A(n4077), .B(n109_adj_219), 
         .Z(n38723)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i61_2_lut.init = 16'h9999;
    LUT4 i25600_4_lut_4_lut (.A(n42680), .B(n37927), .C(n48_adj_370), 
         .D(n34_adj_363), .Z(n50_adj_371)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25600_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i24949_3_lut (.A(\U[10] [6]), .B(\U[11] [6]), .C(i[0]), .Z(n40209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24949_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i36_3_lut_3_lut (.A(n4761), .B(n112_adj_221), 
         .C(n34_adj_722), .Z(n36_adj_723)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i36_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_4010_i12_4_lut (.A(n130), .B(n36666), .C(n15805), .D(i[1]), 
         .Z(n5345)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i12_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_2841_i29_2_lut_rep_846 (.A(n4330), .B(n123), 
         .Z(n42545)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i29_2_lut_rep_846.init = 16'h6666;
    PFUMX i25148 (.BLUT(n40401), .ALUT(n40402), .C0(i[1]), .Z(n40408));
    LUT4 i25855_4_lut_4_lut (.A(n42511), .B(n39164), .C(n42510), .D(n42509), 
         .Z(n39184)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25855_4_lut_4_lut.init = 16'hfff4;
    LUT4 div_4016_LessThan_1553_i59_2_lut_rep_1033 (.A(n2404), .B(n122_adj_228), 
         .Z(n42732)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i59_2_lut_rep_1033.init = 16'h6666;
    LUT4 i25904_4_lut (.A(n42680), .B(n42681), .C(n42682), .D(n37918), 
         .Z(n37932)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25904_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_129 (.A(i[0]), .B(\y[3] [11]), .Z(n36666)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_129.init = 16'h8888;
    LUT4 div_4016_LessThan_2058_i37_2_lut (.A(n3165), .B(n128_adj_232), 
         .Z(n37)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i37_2_lut.init = 16'h6666;
    PFUMX i25149 (.BLUT(n40403), .ALUT(n40404), .C0(i[1]), .Z(n40409));
    LUT4 i1_4_lut_adj_130 (.A(n160_adj_156), .B(i[1]), .C(done_N_1932), 
         .D(n13381), .Z(n30845)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(40[7] 135[14])
    defparam i1_4_lut_adj_130.init = 16'heca0;
    LUT4 i22372_2_lut_3_lut_4_lut (.A(n2404), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n2403), .Z(n37632)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22372_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i22680_4_lut_4_lut (.A(n42680), .B(n37923), .C(n42678), .D(n42679), 
         .Z(n37940)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22680_4_lut_4_lut.init = 16'h000b;
    LUT4 div_4016_LessThan_2058_i55_2_lut_rep_979 (.A(n3156), .B(n119_adj_226), 
         .Z(n42678)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i55_2_lut_rep_979.init = 16'h6666;
    LUT4 i24948_3_lut (.A(\U[8] [6]), .B(\U[9] [6]), .C(i[0]), .Z(n40208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24948_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1553_i57_2_lut_rep_1034 (.A(n2405), .B(n123), 
         .Z(n42733)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i57_2_lut_rep_1034.init = 16'h6666;
    LUT4 mux_4010_i13_4_lut (.A(n127), .B(n36664), .C(n15805), .D(i[1]), 
         .Z(n5344)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i13_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_3206_i24_3_lut (.A(n16_adj_750), .B(n110_adj_220), 
         .C(n45_adj_778), .Z(n24_adj_758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i24_3_lut.init = 16'hcaca;
    LUT4 div_4016_i3340_4_lut (.A(n64_adj_703), .B(n22304), .C(n42786), 
         .D(n30950), .Z(n5523)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3340_4_lut.init = 16'hc0c5;
    LUT4 div_4016_i3339_4_lut (.A(n64_adj_670), .B(n22303), .C(n42786), 
         .D(n42792), .Z(n5522)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3339_4_lut.init = 16'hc0c5;
    PFUMX i25327 (.BLUT(n40579), .ALUT(n40580), .C0(i[1]), .Z(n40587));
    LUT4 div_4016_i3338_4_lut (.A(n64_adj_640), .B(n22302), .C(n42786), 
         .D(n35961), .Z(n5521)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3338_4_lut.init = 16'hc0c5;
    PFUMX i25150 (.BLUT(n40405), .ALUT(n40406), .C0(i[1]), .Z(n40410));
    LUT4 i24947_3_lut (.A(\U[6] [6]), .B(\U[7] [6]), .C(i[0]), .Z(n40207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24947_3_lut.init = 16'hcaca;
    LUT4 div_4016_i3337_4_lut (.A(n64_adj_608), .B(n22301), .C(n42786), 
         .D(n42794), .Z(n5520)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3337_4_lut.init = 16'hc0c5;
    LUT4 div_4016_LessThan_2058_i57_2_lut_rep_980 (.A(n3155), .B(n118_adj_225), 
         .Z(n42679)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i57_2_lut_rep_980.init = 16'h6666;
    LUT4 div_4016_LessThan_1553_i54_3_lut_3_lut (.A(n2405), .B(n123), .C(n46_adj_291), 
         .Z(n54_adj_296)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i54_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_i3336_4_lut (.A(n64_adj_578), .B(n22300), .C(n42786), 
         .D(n35955), .Z(n5519)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3336_4_lut.init = 16'hc0c5;
    LUT4 i23739_2_lut_3_lut_4_lut (.A(n4330), .B(n123), .C(n111), .D(n4318), 
         .Z(n38999)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23739_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i24473_2_lut (.A(n13_adj_747), .B(n11_adj_745), .Z(n39733)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24473_2_lut.init = 16'h1111;
    LUT4 i24946_3_lut (.A(\U[4] [6]), .B(\U[5] [6]), .C(i[0]), .Z(n40206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24946_3_lut.init = 16'hcaca;
    LUT4 div_4016_i3335_4_lut (.A(n64_adj_549), .B(n22299), .C(n42786), 
         .D(n42790), .Z(n5518)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3335_4_lut.init = 16'hc0c5;
    LUT4 div_4016_i3334_4_lut (.A(n64_adj_520), .B(n22298), .C(n42786), 
         .D(n35919), .Z(n5517)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3334_4_lut.init = 16'hc0c5;
    LUT4 i23911_4_lut_4_lut (.A(n42511), .B(n39146), .C(n42513), .D(n42510), 
         .Z(n39171)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23911_4_lut_4_lut.init = 16'h0004;
    LUT4 div_4016_i3333_4_lut (.A(n64_adj_493), .B(n22297), .C(n42786), 
         .D(n30929), .Z(n5516)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3333_4_lut.init = 16'hc0c5;
    PFUMX i25328 (.BLUT(n40581), .ALUT(n40582), .C0(i[1]), .Z(n40588));
    LUT4 div_4016_i3316_4_lut (.A(n37282), .B(n22280), .C(n42786), .D(n64_adj_241), 
         .Z(n5499)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3316_4_lut.init = 16'hc0c5;
    PFUMX i25162 (.BLUT(n40414), .ALUT(n40415), .C0(i[1]), .Z(n40422));
    LUT4 i1_4_lut_adj_131 (.A(n37274), .B(n35922), .C(n37276), .D(n37272), 
         .Z(n37282)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_131.init = 16'hfffe;
    LUT4 i1_2_lut_adj_132 (.A(i[0]), .B(\y[3] [12]), .Z(n36664)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_132.init = 16'h8888;
    LUT4 i1_2_lut_adj_133 (.A(i[0]), .B(\y[3] [9]), .Z(n36662)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_133.init = 16'h8888;
    LUT4 mux_4010_i11_4_lut (.A(n133), .B(n36660), .C(n15805), .D(i[1]), 
         .Z(n5346)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i11_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_134 (.A(n37258), .B(n42820), .C(n37256), .D(n37252), 
         .Z(n37276)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_134.init = 16'hfffe;
    LUT4 i25693_4_lut_4_lut (.A(n42511), .B(n39166), .C(n54_adj_635), 
         .D(n32_adj_623), .Z(n56_adj_636)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25693_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_adj_135 (.A(n119_adj_226), .B(n121_adj_227), .Z(n37258)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_135.init = 16'heeee;
    LUT4 div_4016_LessThan_2058_i42_3_lut_3_lut (.A(n3155), .B(n118_adj_225), 
         .C(n119_adj_226), .Z(n42_adj_367)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i42_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i25163 (.BLUT(n40416), .ALUT(n40417), .C0(i[1]), .Z(n40423));
    LUT4 i1_2_lut_adj_136 (.A(n64), .B(n30872), .Z(n1078)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_136.init = 16'heeee;
    LUT4 div_4016_LessThan_3206_i26_3_lut (.A(n14_adj_748), .B(n117), .C(n31_adj_765), 
         .Z(n26_adj_760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i26_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2681_i35_2_lut (.A(n4090), .B(n122_adj_228), 
         .Z(n35_adj_533)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2681_i35_2_lut.init = 16'h6666;
    LUT4 i24945_3_lut (.A(\U[2] [6]), .B(\U[3] [6]), .C(i[0]), .Z(n40205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24945_3_lut.init = 16'hcaca;
    PFUMX i25164 (.BLUT(n40418), .ALUT(n40419), .C0(i[1]), .Z(n40424));
    LUT4 i22363_3_lut_4_lut (.A(n2405), .B(n123), .C(n47), .D(n42735), 
         .Z(n37623)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22363_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_2918_i61_2_lut_rep_811 (.A(n4428), .B(n106_adj_217), 
         .Z(n42510)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i61_2_lut_rep_811.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i4_4_lut (.A(n132), .B(n131_adj_234), .C(n4883), 
         .D(n708), .Z(n4_adj_738)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i4_4_lut.init = 16'h0c8e;
    LUT4 i1_4_lut_adj_137 (.A(n36500), .B(n64_adj_797), .C(n35925), .D(n36498), 
         .Z(n36422)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_137.init = 16'hfffe;
    LUT4 i1_4_lut_adj_138 (.A(n113_adj_222), .B(n37172), .C(n42815), .D(n115_adj_223), 
         .Z(n36500)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_138.init = 16'hfffe;
    PFUMX i25165 (.BLUT(n40420), .ALUT(n40421), .C0(i[1]), .Z(n40425));
    LUT4 i1_4_lut_adj_139 (.A(n36492), .B(n42821), .C(n126), .D(n128_adj_232), 
         .Z(n36498)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_139.init = 16'hfffe;
    LUT4 i22689_2_lut_3_lut_4_lut (.A(n3155), .B(n118_adj_225), .C(n119_adj_226), 
         .D(n3156), .Z(n37949)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22689_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_3206_i34_3_lut (.A(n32_adj_766), .B(n112_adj_221), 
         .C(n42438), .Z(n34_adj_768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i34_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i10_3_lut (.A(n127_adj_231), .B(n126), .C(n13_adj_747), 
         .Z(n10_adj_744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i10_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2058_i53_2_lut_rep_981 (.A(n3157), .B(n120), 
         .Z(n42680)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i53_2_lut_rep_981.init = 16'h6666;
    PFUMX i25329 (.BLUT(n40583), .ALUT(n40584), .C0(i[1]), .Z(n40589));
    LUT4 div_4016_LessThan_2058_i48_3_lut_3_lut (.A(n3157), .B(n120), .C(n46_adj_369), 
         .Z(n48_adj_370)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i48_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_1553_i53_2_lut_rep_1035 (.A(n2407), .B(n125_adj_230), 
         .Z(n42734)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i53_2_lut_rep_1035.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i11_4_lut (.A(n4777), .B(n127_adj_231), 
         .C(n22267), .D(n4783), .Z(n11_adj_745)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i11_4_lut.init = 16'h663c;
    LUT4 i24944_3_lut (.A(\U[0] [6]), .B(\U[1] [6]), .C(i[0]), .Z(n40204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24944_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_140 (.A(i[0]), .B(\y[3] [10]), .Z(n36660)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_140.init = 16'h8888;
    LUT4 div_4016_i3311_4_lut (.A(n37284), .B(n22275), .C(n42786), .D(n42778), 
         .Z(n5494)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_i3311_4_lut.init = 16'hc0c5;
    LUT4 i23650_3_lut_4_lut (.A(n4330), .B(n123), .C(n19_adj_582), .D(n42546), 
         .Z(n38910)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i23650_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_LessThan_1553_i50_3_lut_3_lut (.A(n2407), .B(n125_adj_230), 
         .C(n48_adj_292), .Z(n50_adj_294)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i50_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_141 (.A(n35916), .B(n131_adj_234), .Z(n37284)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_141.init = 16'heeee;
    LUT4 mux_4010_i8_4_lut (.A(n142), .B(n36656), .C(n15805), .D(i[1]), 
         .Z(n5349)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i8_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_142 (.A(i[0]), .B(\y[3] [7]), .Z(n36656)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_142.init = 16'h8888;
    LUT4 mux_4010_i9_4_lut (.A(n139), .B(n36658), .C(n15805), .D(i[1]), 
         .Z(n5348)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i9_4_lut.init = 16'hca0a;
    LUT4 div_4016_LessThan_3206_i44_3_lut (.A(n42_adj_775), .B(n107_adj_218), 
         .C(n42439), .Z(n44_adj_777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i44_3_lut.init = 16'hcaca;
    LUT4 i25826_3_lut_4_lut (.A(n2407), .B(n125_adj_230), .C(n49_adj_293), 
         .D(n42736), .Z(n37610)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25826_3_lut_4_lut.init = 16'hfff6;
    LUT4 i24936_3_lut (.A(\U[14] [5]), .B(\U[15] [5]), .C(i[0]), .Z(n40196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24936_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2058_i51_2_lut_rep_982 (.A(n3158), .B(n121_adj_227), 
         .Z(n42681)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i51_2_lut_rep_982.init = 16'h6666;
    PFUMX i25177 (.BLUT(n40429), .ALUT(n40430), .C0(i[1]), .Z(n40437));
    LUT4 i25202_3_lut (.A(\U[6] [23]), .B(\U[7] [23]), .C(i[0]), .Z(n40462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25202_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i26_3_lut (.A(n5466), .B(n74_adj_198), .C(n5460), 
         .Z(n107_adj_218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i26_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i8_3_lut (.A(n128_adj_232), .B(n124_adj_229), 
         .C(n17_adj_751), .Z(n8_adj_742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i8_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_5_i25_3_lut (.A(n5467), .B(n75), .C(n5460), .Z(n108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i25_3_lut.init = 16'hcaca;
    LUT4 i25201_3_lut (.A(\U[4] [23]), .B(\U[5] [23]), .C(i[0]), .Z(n40461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25201_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2058_i46_3_lut_3_lut (.A(n3158), .B(n121_adj_227), 
         .C(n122_adj_228), .Z(n46_adj_369)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i46_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2058_i49_2_lut_rep_983 (.A(n3159), .B(n122_adj_228), 
         .Z(n42682)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i49_2_lut_rep_983.init = 16'h6666;
    LUT4 i22667_2_lut_3_lut_4_lut (.A(n3159), .B(n122_adj_228), .C(n121_adj_227), 
         .D(n3158), .Z(n37927)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22667_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_4016_LessThan_2058_i47_2_lut_rep_984 (.A(n3160), .B(n123), 
         .Z(n42683)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i47_2_lut_rep_984.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i50_3_lut (.A(n22_adj_756), .B(n104_adj_216), 
         .C(n57_adj_789), .Z(n50_adj_783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i50_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i64_4_lut (.A(n40_adj_774), .B(n37376), 
         .C(n42437), .D(n40057), .Z(n4885)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i64_4_lut.init = 16'hcacc;
    PFUMX i25330 (.BLUT(n40585), .ALUT(n40586), .C0(i[1]), .Z(n40590));
    PFUMX i25178 (.BLUT(n40431), .ALUT(n40432), .C0(i[1]), .Z(n40438));
    L6MUX21 div_4016_LessThan_1337_i64 (.D0(n56_adj_274), .D1(n62_adj_277), 
            .SD(n37544), .Z(n64_adj_278));
    LUT4 div_4016_LessThan_3206_i35_4_lut (.A(n4765), .B(n115_adj_223), 
         .C(n22255), .D(n4783), .Z(n35_adj_769)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i35_4_lut.init = 16'h663c;
    LUT4 div_4016_LessThan_2918_i30_3_lut_3_lut (.A(n4428), .B(n106_adj_217), 
         .C(n14_adj_611), .Z(n30_adj_622)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2918_i30_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_2058_i44_3_lut_3_lut (.A(n3160), .B(n123), .C(n36_adj_364), 
         .Z(n44_adj_368)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2058_i44_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_4016_LessThan_3206_i6_3_lut (.A(n130_adj_233), .B(n129), .C(n7_adj_741), 
         .Z(n6_adj_740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i6_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i62_rep_16_4_lut (.A(n48_adj_781), .B(n37377), 
         .C(n42437), .D(n40059), .Z(n37376)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i62_rep_16_4_lut.init = 16'hcacc;
    LUT4 i24797_4_lut (.A(n61_adj_793), .B(n59_adj_791), .C(n57_adj_789), 
         .D(n40033), .Z(n40057)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24797_4_lut.init = 16'h0100;
    LUT4 div_4016_LessThan_3206_i60_rep_17_4_lut (.A(n52_adj_784), .B(n37378), 
         .C(n42437), .D(n40061), .Z(n37377)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i60_rep_17_4_lut.init = 16'hcacc;
    LUT4 div_4016_LessThan_3206_i54_rep_20_3_lut (.A(n20_adj_754), .B(n102), 
         .C(n61_adj_793), .Z(n37380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i54_rep_20_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_143 (.A(i[0]), .B(\y[3] [8]), .Z(n36658)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_143.init = 16'h8888;
    LUT4 i24747_4_lut (.A(n49_adj_782), .B(n47_adj_780), .C(n45_adj_778), 
         .D(n39995), .Z(n40007)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24747_4_lut.init = 16'h0100;
    LUT4 div_4016_LessThan_1553_i55_2_lut_rep_1036 (.A(n2406), .B(n124_adj_229), 
         .Z(n42735)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i55_2_lut_rep_1036.init = 16'h6666;
    LUT4 i24735_2_lut (.A(n43_adj_776), .B(n39987), .Z(n39995)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i24735_2_lut.init = 16'h1111;
    LUT4 div_4016_mux_5_i5_3_lut (.A(n5487), .B(n95_adj_212), .C(n5460), 
         .Z(n128_adj_232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i5_3_lut.init = 16'hcaca;
    LUT4 mux_4010_i7_4_lut (.A(n145), .B(n36654), .C(n15805), .D(i[1]), 
         .Z(n5350)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i7_4_lut.init = 16'hca0a;
    LUT4 div_4016_mux_5_i9_3_lut (.A(n5483), .B(n91_adj_209), .C(n5460), 
         .Z(n124_adj_229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_5_i9_3_lut.init = 16'hcaca;
    PFUMX i25179 (.BLUT(n40433), .ALUT(n40434), .C0(i[1]), .Z(n40439));
    LUT4 mux_4010_i10_4_lut (.A(n136), .B(n36662), .C(n15805), .D(i[1]), 
         .Z(n5347)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(105[14] 112[8])
    defparam mux_4010_i10_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_144 (.A(i[0]), .B(\y[3] [6]), .Z(n36654)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(99[19:20])
    defparam i1_2_lut_adj_144.init = 16'h8888;
    LUT4 i24935_3_lut (.A(\U[12] [5]), .B(\U[13] [5]), .C(i[0]), .Z(n40195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24935_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_3_i16_3_lut (.A(n5341), .B(n18_adj_178), .C(n5325), 
         .Z(n879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i16_3_lut.init = 16'hcaca;
    LUT4 i25843_4_lut (.A(n42650), .B(n38136), .C(n42651), .D(n38127), 
         .Z(n38148)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i25843_4_lut.init = 16'hfbff;
    LUT4 div_4016_LessThan_3206_i30_3_lut (.A(n12_adj_746), .B(n115_adj_223), 
         .C(n35_adj_769), .Z(n30_adj_764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i30_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_3_i17_3_lut (.A(n5340), .B(n17_adj_177), .C(n5325), 
         .Z(n878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i17_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3137_i37_2_lut_rep_754 (.A(n4764), .B(n115_adj_223), 
         .Z(n42453)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3137_i37_2_lut_rep_754.init = 16'h6666;
    LUT4 div_4016_LessThan_3206_i15_4_lut (.A(n4775), .B(n125_adj_230), 
         .C(n22265), .D(n4783), .Z(n15_adj_749)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i15_4_lut.init = 16'h663c;
    LUT4 i22658_3_lut_4_lut (.A(n3160), .B(n123), .C(n37), .D(n42684), 
         .Z(n37918)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam i22658_3_lut_4_lut.init = 16'h0009;
    LUT4 div_4016_mux_3_i18_3_lut (.A(n5339), .B(n16_adj_176), .C(n5325), 
         .Z(n877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i18_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_3206_i16_3_lut (.A(n123), .B(n111), .C(n43_adj_776), 
         .Z(n16_adj_750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_3206_i16_3_lut.init = 16'hcaca;
    LUT4 div_4016_mux_3_i19_3_lut (.A(n5338), .B(n15_adj_175), .C(n5325), 
         .Z(n876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_mux_3_i19_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_2841_i27_2_lut_rep_847 (.A(n4331), .B(n124_adj_229), 
         .Z(n42546)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i27_2_lut_rep_847.init = 16'h6666;
    LUT4 div_4016_LessThan_2841_i18_3_lut_3_lut (.A(n4331), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n18_adj_581)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_2841_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24934_3_lut (.A(\U[10] [5]), .B(\U[11] [5]), .C(i[0]), .Z(n40194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24934_3_lut.init = 16'hcaca;
    LUT4 div_4016_LessThan_1553_i46_3_lut_3_lut (.A(n2406), .B(n124_adj_229), 
         .C(n128_adj_232), .Z(n46_adj_291)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/matrix_inv/backward.v(116[21:37])
    defparam div_4016_LessThan_1553_i46_3_lut_3_lut.init = 16'hd4d4;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

