// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Tue Sep 23 20:22:52 2025
//
// Verilog Description of module FFT
//

module FFT (clk, rst_n, in_valid, din_r, din_i, out_valid, dout_r, 
            dout_i) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(12[8:11])
    input clk;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    input rst_n;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(14[7:12])
    input in_valid;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(15[7:15])
    input [11:0]din_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    input [11:0]din_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    output out_valid;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(18[8:17])
    output [15:0]dout_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    output [15:0]dout_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire GND_net, VCC_net, rst_n_c, in_valid_c, din_r_c_11, din_r_c_10, 
        din_r_c_9, din_r_c_8, din_r_c_7, din_r_c_6, din_r_c_5, din_r_c_4, 
        din_r_c_3, din_r_c_2, din_r_c_1, din_r_c_0, din_i_c_11, din_i_c_10, 
        din_i_c_9, din_i_c_8, din_i_c_7, din_i_c_6, din_i_c_5, din_i_c_4, 
        din_i_c_3, din_i_c_2, din_i_c_1, din_i_c_0, out_valid_c, dout_r_c_15, 
        dout_r_c_14, dout_r_c_13, dout_r_c_12, dout_r_c_11, dout_r_c_10, 
        dout_r_c_9, dout_r_c_8, dout_r_c_7, dout_r_c_6, dout_r_c_5, 
        dout_r_c_4, dout_r_c_3, dout_r_c_2, dout_r_c_1, dout_r_c_0, 
        dout_i_c_15, dout_i_c_14, dout_i_c_13, dout_i_c_12, dout_i_c_11, 
        dout_i_c_10, dout_i_c_9, dout_i_c_8, dout_i_c_7, dout_i_c_6, 
        dout_i_c_5, dout_i_c_4, dout_i_c_3, dout_i_c_2, dout_i_c_1, 
        dout_i_c_0;
    wire [15:0]\result_r[0] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[1] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[2] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[3] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[4] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[5] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[6] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[7] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[8] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[9] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[10] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[11] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[12] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[13] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[14] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[15] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[16] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[17] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[18] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[19] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[20] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[21] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[22] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[23] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[24] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[25] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[26] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[27] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[28] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[29] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[30] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_r[31] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(24[20:28])
    wire [15:0]\result_i[0] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[1] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[2] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[3] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[4] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[5] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[6] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[7] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[8] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[9] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[10] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[11] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[12] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[13] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[14] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[15] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[16] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[17] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[18] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[19] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[20] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[21] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[22] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[23] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[24] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[25] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[26] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[27] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[28] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[29] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[30] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [15:0]\result_i[31] ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(25[20:28])
    wire [5:0]count_y;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(30[21:28])
    
    wire n33616, n12334, n12333;
    wire [23:0]din_r_reg;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(33[19:28])
    wire [23:0]op_r_23__N_1106;
    wire [23:0]din_i_reg;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(33[29:38])
    
    wire in_valid_reg, r4_valid, n34076;
    wire [1:0]no5_state;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(35[11:20])
    
    wire s5_count, over, next_out_valid;
    wire [4:0]y_1_delay;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(40[10:19])
    wire [23:0]out_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(42[13:18])
    wire [23:0]out_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(42[19:24])
    
    wire n34843, n34075, n8958, n8952, n8956, n8966, n8954, n8953;
    wire [23:0]rom16_w_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(52[12:21])
    
    wire n10735, n10734, n9099, n9098;
    wire [23:0]rom16_w_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(52[22:31])
    wire [23:0]shift_16_dout_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(53[12:27])
    wire [23:0]shift_16_dout_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(53[28:43])
    
    wire n8962, n8955;
    wire [1:0]rom8_state;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(56[12:22])
    wire [23:0]rom8_w_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(57[12:20])
    
    wire n9096, n11130;
    wire [23:0]rom8_w_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(57[21:29])
    
    wire n8577;
    wire [23:0]shift_8_dout_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(58[12:26])
    wire [23:0]shift_8_dout_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(58[27:41])
    
    wire n8591, n8576;
    wire [23:0]radix_no1_op_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(60[12:26])
    wire [23:0]radix_no1_op_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(60[27:41])
    wire [1:0]rom4_state;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(64[12:22])
    
    wire n34074, n32133, n12291, n11137;
    wire [23:0]rom4_w_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(65[12:20])
    
    wire n33699, n11132, n11138, n11134;
    wire [23:0]rom4_w_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(65[21:29])
    
    wire n11131, n11557, n8582;
    wire [23:0]shift_4_dout_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(66[12:26])
    wire [23:0]shift_4_dout_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(66[27:41])
    
    wire n10733, n8575, n9089, n33313;
    wire [23:0]rom2_w_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(72[12:20])
    
    wire n12172, n12065, n12066, n12067, n12068, n12069, n12070, 
        n12071, n12072, n12073, n12074, n12075, n12077;
    wire [23:0]shift_2_dout_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(73[12:26])
    wire [23:0]shift_2_dout_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(73[27:41])
    
    wire n11141, n11140, n11136, n34073, n33698, n34072, n34071, 
        n34070, n33259, n33615, n34069, n33697, n34068, n34067, 
        n34066, n33332, n33333, n34065, n33696, n34064, n34063, 
        n34061, n33266, n33288, n34060, n33695, n34059, n34058;
    wire [23:0]shift_1_dout_r;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(78[12:26])
    wire [23:0]shift_1_dout_i;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(78[27:41])
    
    wire n11129, n11128;
    wire [15:0]next_dout_r_15__N_1029;
    wire [15:0]next_dout_i_15__N_1045;
    
    wire rst_n_N_2;
    wire [511:0]result_r_ns_0__15__N_3;
    wire [511:0]result_i_ns_0__15__N_517;
    
    wire next_over_N_1081;
    wire [23:0]op_i_23__N_1154;
    wire [23:0]delay_r_23__N_1178;
    wire [23:0]delay_i_23__N_1202;
    
    wire n12453, n12452, n12451, n12450, n12449, n12448;
    wire [48:0]op_r_23__N_1268;
    
    wire n12447, n12344, n12345, n12346, n12347, n12348, n12349, 
        n12350, n12351, n12352, n12353, n32132;
    wire [48:0]op_r_23__N_1226;
    wire [41:0]op_r_23__N_1082;
    
    wire n319;
    wire [65:0]op_i_23__N_1310;
    wire [41:0]op_i_23__N_1130;
    
    wire n10728, n8977, n10727, n10730, n8973, n10718, n8967, 
        n65, n8976, n10721, n9088, n9102, n9090, n9105, n8972, 
        n9100, n10725, n9084, n10729, n8969, n9104, n9092, n8957, 
        n12446, n12368, n12445, n65_adj_6358, n12444, n66, n69, 
        n73, n68, n70, n77, n71, n8959, n72, n74, n75, n9103, 
        n76, n78, n81, n79, n80, n82, n85, n83, n84, n86, 
        n87, n11171, n8964, n88, n89, n9101, n8963, n9087, n8960, 
        n8961, n8965;
    wire [383:0]dout_r_23__N_2506;
    wire [383:0]dout_i_23__N_3274;
    
    wire n33614, n32131, n34057, n33457, n33613, n33694, n33693, 
        n33692, n34056, n33691, n33344, n34055, n33689, n33688, 
        n33612, n33687, n34631, n33456, n33611, n34054, n33455, 
        n33610, n33686, n34053, n34052, n33685, n33343, n34051, 
        n34050, n33684, n33609, n33608, n33683, n33454, n34049, 
        n34048, n33682, n34047, n33681, n34046, n33680, n33679, 
        n34045, n33678, n34044, n34043, n33677, n34042, n34041, 
        n33676, n33675, n33453, n34040, n33607, n34039, n33674, 
        n33673, n33342, n34038, n33672, n33671, n33606, n33331, 
        n34037, n33605, n34036, n33670, n33669, n33452, n34035, 
        n33668, n34034, n34033, n33667, n33666, n33451, n33341, 
        n33299, n33665, n33604, n34032, n33603, n33602, n34030, 
        n34029, n33664, n33663, n33450, n33601, n33662, n33661, 
        n33600, n34028, n34027, n33660, n33449, n34026, n33658, 
        n33657, n33656, n33599, n34025, n33655, n33448, n33654, 
        n34024, n33653, n33598, n34023, n33652, n34022, n33447, 
        n34021, n33651, n33596, n33650, n33446, n33595, n33594, 
        n33649, n8574, n8573, n33327, n33593, n8572, n8703, n8706, 
        n8708, n8571, n8570, n8569, n8568, n8580, n8701, n34020, 
        n34019, n33648, n34018, n33647, n33646, n33645, n33644, 
        n34017, n33445, n33592, n34016, n33444, n33591, n34630, 
        n33643, n34015, n34014, n34013, n8705, n33321, n33265, 
        n8707, n8585, n8587, n34012, n33590, n33589, n34629, n33642, 
        n34011, n33443, n33588, n33641, n33324, n34010, n33587, 
        n33586, n33640, n34009, n33441, n33328, n33585, n33639, 
        n34008, n33584, n33638, n34007, n33637, n34006, n33636, 
        n33635, n33634, n33633, n34005, n33440, n34628, n33583, 
        n34004, n33582;
    wire [5:0]count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(11[11:16])
    
    wire n34575, n33581, n33632, n34003, n34002, n34627, n12292, 
        n12264;
    wire [23:0]op_r_23__N_1106_adj_7319;
    wire [23:0]op_i_23__N_1154_adj_7320;
    
    wire n9097, n8589, n34589, n8590, n3, n119;
    wire [48:0]op_r_23__N_1268_adj_7324;
    
    wire n12321, n12300, n12301, n12302, n12303, n12304, n12305, 
        n12306, n12307, n12308, n12309, n12322, n12323, n12324, 
        n12325, n12326, n12327, n12328, n12329, n12330, n12331;
    wire [48:0]op_r_23__N_1226_adj_7326;
    wire [41:0]op_r_23__N_1082_adj_7327;
    
    wire n319_adj_6495;
    wire [65:0]op_i_23__N_1310_adj_7329;
    wire [41:0]op_i_23__N_1130_adj_7330;
    
    wire n9091, n67, n10722, n8588, n10726, n9080, n89_adj_6552, 
        n88_adj_6553, n87_adj_6554, n86_adj_6555, n85_adj_6556, n84_adj_6557, 
        n83_adj_6558, n82_adj_6559, n81_adj_6560, n80_adj_6561, n9093, 
        n79_adj_6562, n78_adj_6563, n77_adj_6564, n76_adj_6565, n75_adj_6566, 
        n74_adj_6567, n73_adj_6568, n72_adj_6569, n71_adj_6570, n70_adj_6571, 
        n9081, n69_adj_6572, n68_adj_6573, n9082, n67_adj_6574, n11142, 
        n9095, n66_adj_6575, n10720, n65_adj_6576, n9094, n10724, 
        n9085, n10719, n9083, n10723, n10732, valid;
    wire [191:0]dout_r_23__N_4286;
    wire [191:0]dout_i_23__N_4670;
    
    wire n34626, n34001, n8696, n8697, n8698, n8699, n33580, n8586, 
        n8593, n8711, n8712, n8713, n8714, n8715, n8716, n8717, 
        n8718, n8719, n8720, n8721, n33999, n33631, n33311, n29782, 
        n8824, n8825, n12082, n8826, n8827, n8828, n8829, n8830, 
        n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, 
        n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, 
        n8847, n8848, n8849, n11564, n12087, n11561, n12175, n11570, 
        n33998, n11567, n12086, n11575, n11573, n12085, n12083, 
        n12084, n33301;
    wire [3:0]s_count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(12[11:18])
    
    wire n33997, n8709, n12078, n28591, n28589, n34625, n34588;
    wire [23:0]op_r_23__N_1106_adj_7370;
    wire [23:0]op_i_23__N_1154_adj_7371;
    
    wire n8968, n8975, n34624, n119_adj_6625, n12314, n12315, n12316, 
        n12317, n12318, n12319, n12320;
    wire [48:0]op_r_23__N_1268_adj_7375;
    
    wire n12332, n12270, n12271, n12272, n12273, n12274, n12275, 
        n12276, n12277, n12278, n12279, n12280, n12281, n12282, 
        n12283, n12284, n12285, n12286, n12287, n12288, n12289, 
        n12290;
    wire [48:0]op_r_23__N_1226_adj_7377;
    wire [41:0]op_r_23__N_1082_adj_7378;
    
    wire n319_adj_6714;
    wire [65:0]op_i_23__N_1310_adj_7380;
    wire [41:0]op_i_23__N_1130_adj_7381;
    
    wire n11143, n9086, n11135, valid_adj_6771;
    wire [95:0]dout_r_23__N_5203;
    wire [95:0]dout_i_23__N_5395;
    
    wire n33439, n11562, n11560, n11559, n11568, n11566, n11565, 
        n11574, n11572, n11571, n11577, n11576, n11563, n65_adj_6772, 
        n11569, n32130, n32129, n11133, n12336, n12294, n12293, 
        n12263, n12262, n12335, n8583, n8704, n12261;
    wire [2:0]s_count_adj_7402;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(12[11:18])
    
    wire n8710, state_1__N_5502, n33630, n33996, n34623, n33995, 
        n34622, n8702;
    wire [23:0]op_r_23__N_1106_adj_7425;
    wire [23:0]op_i_23__N_1154_adj_7426;
    wire [23:0]delay_r_23__N_1178_adj_7427;
    wire [23:0]delay_i_23__N_1202_adj_7428;
    wire [48:0]op_r_23__N_1268_adj_7430;
    
    wire n12240, n12241, n12242, n12243, n12244, n12245, n12246, 
        n12247, n12248, n12249, n12250, n12251, n12252, n12253, 
        n12254, n12255, n12256, n12257, n12258, n12259;
    wire [48:0]op_r_23__N_1226_adj_7432;
    wire [41:0]op_r_23__N_1082_adj_7433;
    
    wire n319_adj_6944, n11148, n11149, n11150, n11151, n11152, 
        n11153, n11154, n11155, n11156, n11157, n11158, n11159, 
        n11160, n11161, n11162, n11163, n11164, n11165, n11166, 
        n11167, n11168, n11169, n11170;
    wire [65:0]op_i_23__N_1310_adj_7435;
    wire [41:0]op_i_23__N_1130_adj_7436;
    
    wire n8579, n11126, valid_adj_7001;
    wire [47:0]dout_r_23__N_5681;
    wire [47:0]dout_i_23__N_5777;
    
    wire n8592, n8581, n34621, n8700;
    wire [5:0]count_adj_7456;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(11[11:16])
    
    wire n33629, n11127, n10006;
    wire [1:0]s_count_adj_7458;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(12[11:18])
    
    wire n11578, n10005, n10004;
    wire [1:0]state_1__N_5843;
    
    wire n10003, n12076, n10002, n12173, n12088, n12089, n12260, 
        n12174;
    wire [23:0]op_r_23__N_1106_adj_7481;
    
    wire n10001, n34620, n33579, n32128, n32127;
    wire [23:0]op_i_23__N_1154_adj_7482;
    
    wire n32126, n32125, n12176, n10000, n12080;
    wire [23:0]delay_r_23__N_1178_adj_7483;
    wire [23:0]delay_i_23__N_1202_adj_7484;
    
    wire n12081, n12079, n9999, n7614, n7613, n7612, n7611, n7610;
    wire [48:0]op_r_23__N_1268_adj_7486;
    
    wire n12152, n12153, n12154, n12155, n12156, n12157, n12158, 
        n12159, n12160, n12161, n12162, n12163, n12164, n12165, 
        n12166, n12167, n12168, n12169, n12170, n12171;
    wire [48:0]op_r_23__N_1226_adj_7488;
    wire [41:0]op_r_23__N_1082_adj_7489;
    
    wire n7609, n7608, n7607, n7606, n7605, n7604, n7603, n7602, 
        n11139, n11579, n319_adj_7163, n89_adj_7164, n88_adj_7165, 
        n87_adj_7166;
    wire [65:0]op_i_23__N_1310_adj_7491;
    wire [41:0]op_i_23__N_1130_adj_7492;
    
    wire n7601, n7600, n7599, n7598, n7597, n7596, n7595, n7594, 
        n7593, valid_adj_7215, n7592;
    wire [23:0]dout_r_23__N_5926;
    wire [23:0]dout_i_23__N_5974;
    
    wire n7591, n33320, n33578, n33994, n33627, n33993, n33992, 
        n33991, n33317, n33319, n33990, n33626, n33989, n33988, 
        n7561, n7560, n7559, n7558, n7557, n7556, n7555, n7554, 
        n7553, n7552, n7551, n7550, n7549, n7548, n7547, n7546, 
        n7545, n7544, n7543, n7542, n7541, n7540, n7539, n7538, 
        n33987, n33316, n32925, n33986, n33625, n33985, n33984, 
        n33983, n33314, n33982, n33624, n33981, n7508, n7507, 
        n7506, n7505, n7504, n7503, n7502, n7501, n7500, n7499, 
        n7498, n7497, n7496, n7495, n7494, n7493, n7492, n7491, 
        n7490, n7489, n7488, n7487, n7486, n7485, n33980, n33979, 
        n33312, n34619, n33978, n33623, n33977, n33976, n33975, 
        n33310, n33974, n7455, n7454, n7453, n7452, n7451, n7450, 
        n7449, n7448, n7447, n7446, n7445, n7444, n7443, n7442, 
        n7441, n7440, n7439, n7438, n7437, n7436, n7435, n7434, 
        n7433, n7432, n33622, n33973, n33972, n33971, n33309, 
        n33970, n33621, n33968, n33967, n33966, n33308, n86_adj_7216, 
        n85_adj_7217, n8974, n9998, n84_adj_7218, n83_adj_7219, n9997, 
        n82_adj_7220, n81_adj_7221, n11558, n80_adj_7222, n79_adj_7223, 
        n78_adj_7224, n77_adj_7225, n8970, n76_adj_7226, n75_adj_7227, 
        n74_adj_7228, n33965, n33620, n33619, n11556, n73_adj_7229, 
        n72_adj_7230, n9983, n71_adj_7231, n9984, n70_adj_7232, n33577, 
        n69_adj_7233, n68_adj_7234, n9985, n9986, n10731, n9987, 
        n9988, n33964, n31572, n33618, n31574, n33963, n31576, 
        n31578, n33962, n31580, n33961, n31582, n31584, n31586, 
        n33307, n31588, n33576, n31590, n31592, n31594, n67_adj_7235, 
        n66_adj_7236, n9989, n65_adj_7237, n8584, n12338, n33960, 
        n33617, n33959, n33958, n33957, n33306, n33956, n33575, 
        n33955, n33954, n33953, n33305, n12337, n31670, n31672, 
        n31674, n33952, n31676, n33438, n31678, n33951, n31680, 
        n31682, n33950, n31684, n32124, n9990, n9991, n33949, 
        n31474, n31476, n31478, n33286, n31480, n31482, n31484, 
        n31486, n31488, n33948, n31490, n33574, n31492, n33947, 
        n31494, n31496, n8971, n33946, n9992, n33945, n33285, 
        n33944, n33437, n33943, n33942, n33941, n33284, n33264, 
        n33940, n33573, n33939, n32123, n9993, n31703, n33937, 
        n31705, n33936, n31707, n31709, n31711, n33282, n31713, 
        n33572, n31715, n31717, n9994, n6514, n31425, n31427, 
        n33935, n31429, n33436, n31431, n33934, n31433, n34618, 
        n31435, n33933, n31437, n33932, n31439, n31441, n31443, 
        n33281, n31445, n31447, n8578, n9995, n31376, n31378, 
        n31380, n33931, n31382, n33571, n31384, n33930, n31386, 
        n34617, n31388, n33929, n31390, n33928, n31392, n31394, 
        n31396, n33280, n31398, n9996, n34802, n34801, n29815, 
        n34800, n33927, n32122, n32392, n33435, n32120, n33926, 
        n17, n32119, n32391, n32390, n32118, n32117, n32116, n32115, 
        n32114, n32113, n34799, n32112, n32111, n33925, clk_c_enable_2310, 
        n32386, n32110, n32109, n32108, n32107, n29828, n33570, 
        n34795, n32385, n34794, n34587, clk_c_enable_2259, n34616, 
        n33924, n35, n34, n33, n32, n31, n30, n32106, n33923, 
        n32105, n32384, n32104, n32103, n19995, n34615, n33434, 
        n33922, n33569, n34614, n29827, n29826, n33921, n29824, 
        n29823, n29822, n33920, n29820, n29819, n29816, n66_adj_7238, 
        n67_adj_7239, n68_adj_7240, n69_adj_7241, n70_adj_7242, n71_adj_7243, 
        n72_adj_7244, n73_adj_7245, n74_adj_7246, n75_adj_7247, n76_adj_7248, 
        n77_adj_7249, n78_adj_7250, n79_adj_7251, n80_adj_7252, n81_adj_7253, 
        n82_adj_7254, n83_adj_7255, n84_adj_7256, n85_adj_7257, n86_adj_7258, 
        n87_adj_7259, n88_adj_7260, n89_adj_7261, n111, n114, n117, 
        n120, n123, n126, n111_adj_7262, n114_adj_7263, n117_adj_7264, 
        n120_adj_7265, n123_adj_7266, n126_adj_7267, n66_adj_7268, n67_adj_7269, 
        n68_adj_7270, n69_adj_7271, n70_adj_7272, n71_adj_7273, n72_adj_7274, 
        n73_adj_7275, n74_adj_7276, n75_adj_7277, n76_adj_7278, n77_adj_7279, 
        n78_adj_7280, n79_adj_7281, n80_adj_7282, n81_adj_7283, n82_adj_7284, 
        n83_adj_7285, n84_adj_7286, n85_adj_7287, n86_adj_7288, n87_adj_7289, 
        n88_adj_7290, n89_adj_7291, n34841, n33919, n34789, n34788, 
        n33918, n33917, n33433, n34787, n33916, n34839, n33915, 
        n34612, n34785, n33914, n34613, n33913, n33912, n33911, 
        n33568, n34611, n33910, n33432, n33909, n33908, n33431, 
        n33340, n33567, n33906, n33905, n34610, n34609, n33430, 
        n33904, n33429, n33903, n33902, n34779, n34778, n33901, 
        n34608, n33565, n34777, n33900, n34607, n33261, n34776, 
        n33899, n33428, n33898, n33564, n33897, n33427, clk_c_enable_2285, 
        n33426, n33896, n33563, n33425, n33895, n34606, n33894, 
        n33893, n33562, n33424, n33260, n34771, n33561, n33892, 
        n33891, n33890, n34770, n34769, n33889, n34586, n33888, 
        clk_c_enable_2299, n33303, n33423, clk_c_enable_1419, n33560, 
        clk_c_enable_2305, n34762, n34761, n34760, n34759, n34757, 
        n34756, n34755, n34754, n34753, n34752, n34751, clk_c_enable_2300, 
        clk_c_enable_1396, clk_c_enable_1373, n33559, n34742, n34741, 
        n34740, n34739, n34738, n34737, n34736, n34735, n34734, 
        n34733, n34731, n34730, n34729, n34727, n34726, n34725, 
        n34724, n34723, n33051, n33422, n33558, n33887, n34585, 
        n33886, n33885, n33263, n33557, n33884, n33556, n33883, 
        n34247, n33882, n33881, n33304, n34605, n34246, n33880, 
        n33421, n33879, n34245, n33878, n33877, n33296, n34244, 
        n33875, n33420, n33874, n34243, n33873, n33872, n34720, 
        n33294, n33262, n34242, n33871, n33555, n33870, n34241, 
        n33869, n33868, n33292, n34240, n33867, n33419, n33866, 
        n34239, n33865, n33864, n33270, n34238, n33863, n33554, 
        n33862, n34237, n33861, n33553, n34520, n33552, n34604, 
        n33551, n34812, n33295, n34578, n34584, n34717, n33550, 
        n34603, n33549, n33548, n34602, n33547, n34601, n33326, 
        n33546, n33289, n33545, n33544, n33543, n33323, n33542, 
        n34600, n33541, n34599, n33540, n33300, n33539, n34716, 
        n33538, n33537, n34715, n33536, n34714, n33534, n34713, 
        n34236, n33418, n33860, n33859, n34712, n33858, n33417, 
        n33298, n30503, n30499, n33857, n34711, n34710, n34709, 
        n34708, n34707, n34706, n34705, n34704, n34703, n34702, 
        n30207, n34701, n30203, n30197, n30191, n30179, n34235, 
        n33856, n33533, n34700, n30041, n30040, n34699, n34698, 
        n33293, n34697, n28598, n34234, n33855, n33854, n34233, 
        n33853, n33416, n33339, n33532, n33415, n33531, n33852, 
        n34232, n33851, n33414, n33530, n33850, n34231, n33315, 
        n33849, n33529, n34230, n33413, n33412, n33528, n33848, 
        n33410, n33527, n34696, n34598, n33526, n34597, n33013, 
        n33525, n33030, n33847, n34229, n34228, n34227, n34226, 
        n34225, n34224, n34223, n34222, n34221, n34220, n34219, 
        n34218, n34216, n34215, n34214, n34213, n34212, n34211, 
        n34210, n34209, n34208, n34207, n33846, n34206, n34205, 
        n34204, n34203, n34202, n34201, n34200, n34199, n34198, 
        n34197, n34196, n34195, n34194, n34193, n34192, n34191, 
        n34190, n34189, n34188, n34187, n34185, n34184, n33844, 
        n34695, n33302, n34694, n34183, n34693, n33843, n34182, 
        n6, n34692, n33409, n33842, n33841, n34691, n34690, n33269, 
        n34689, n33268, n34688, n33524, n33329, n33330, n33840, 
        n34811, n34181, n33839, n33408, n33838, n33523, n6_adj_7292, 
        n5, n34180, n33522, n34179, n34687, n34686, n34178, n33837, 
        n34685, n33407, n33836, n34177, n33835, n32928, n34684, 
        n34683, n34176, n34682, n33834, n34681, n33267, n33521, 
        n34175, n34174, n33833, n34680, n32944, n34679, n34678, 
        n33406, n34677, n34676, n34173, n34675, n20103, n33520, 
        n34577, n33519, n33405, n34576, n20095, n34583, n34582, 
        n20089, n34581, n34580, n34674, n32102, n32101, n32383, 
        n32100, n32099, n32382, n32098, n32097, n32381, n33832, 
        n32094, n32380, n34673, n32093, n32092, n32379, n32091, 
        n32090, n32378, n32089, n32088, n32377, n32087, n32086, 
        n32376, n32085, n32084, n32375, n32083, n32082, n32374, 
        n33258, n32081, n32080, n32373, n32079, n32078, n32372, 
        n33831, n32077, n32076, n32371, n32075, n32074, n32370, 
        n32073, n32072, n32369, n32071, n32070, n32368, n33830, 
        n34172, n32069, n32068, n32367, n32067, n32066, n32366, 
        n33518, n32065, n32064, n32365, n32063, n32062, n32364, 
        n33829, n34171, n32061, n32060, n32363, n32059, n32058, 
        n33404, n34170, n32057, n32056, n32360, n33517, n32053, 
        n32359, n33403, n33828, n32052, n32051, n32358, n32050, 
        n32049, n32357, n33516, n32048, n32047, n32356, n32046, 
        n32045, n32355, n33297, n33827, n32044, n32043, n32354, 
        n32042, n32041, n32353, n33515, n32040, n32039, n32352, 
        n33514, n32037, n32351, n33826, n32036, n32035, n32350, 
        n32034, n32033, n32349, n33513, n32032, n32031, n32347, 
        n32030, n32029, n32346, n33512, n32028, n32027, n32345, 
        n32026, n33511, n32344, n33402, n33401, n32022, n32343, 
        n32021, n32020, n32342, n33510, n32019, n32018, n32341, 
        n32017, n32016, n32340, n32015, n32014, n34169, n32013, 
        n32012, n32338, n32011, n32337, n32008, n32007, n32336, 
        n33825, n32006, n32005, n32335, n32004, n32003, n32334, 
        n34168, n34167, n32002, n32001, n32333, n32000, n31999, 
        n32332, n33400, n31998, n31997, n32331, n33399, n33509, 
        n32330, n33508, n33824, n33507, n31992, n32329, n31991, 
        n31990, n32328, n33398, n31989, n31988, n32327, n31987, 
        n31986, n32326, n33283, n33397, n31985, n31984, n32325, 
        n31983, n31982, n32324, n33506, n31981, n31980, n31979, 
        n31978, n32322, n33823, n33822, n31977, n31976, n32321, 
        n31975, n31974, n32320, n33505, n31973, n31972, n32319, 
        n31971, n31970, n32318, n33396, n33503, n31969, n31968, 
        n32317, n31967, n31966, n32316, n33395, n31964, n32315, 
        n31963, n31962, n32314, n33394, n33502, n31961, n31960, 
        n32313, n31959, n31958, n32312, n33501, n31957, n31956, 
        n32311, n31955, n31954, n34672, n31953, n33393, n32308, 
        n34166, n31949, n32307, n31948, n31947, n32306, n31946, 
        n31945, n32305, n34165, n33500, n31944, n31943, n32304, 
        n31942, n31941, n32303, n33821, n31940, n31939, n32302, 
        n31938, n31936, n32301, n34164, n33392, n31935, n31934, 
        n32300, n31933, n31932, n32299, n33820, n31931, n31930, 
        n32298, n31929, n31928, n32297, n33819, n33499, n31927, 
        n31926, n33818, n31925, n33391, n32294, n33817, n31923, 
        n31922, n32293, n31921, n31920, n32292, n33390, n31919, 
        n34163, n32291, n31917, n31916, n32290, n31915, n31914, 
        n32289, n31913, n31912, n32288, n33816, n31911, n31910, 
        n32287, n31909, n31908, n32286, n33498, n31907, n31906, 
        n32285, n33389, n33815, n32284, n33813, n31901, n32283, 
        n31900, n31899, n33388, n31898, n31897, n32280, n31896, 
        n31895, n32279, n33497, n33496, n31894, n31893, n32278, 
        n31892, n31891, n32277, n33387, n31890, n34162, n32276, 
        n31888, n31887, n32275, n34161, n34160, n31886, n31885, 
        n32274, n31884, n31883, n32273, n33495, n31882, n31881, 
        n32272, n31880, n31879, n32271, n33386, n33385, n31878, 
        n31877, n32270, n31876, n31875, n32269, n33384, n31874, 
        n33812, n33383, n31872, n31871, n32266, n33494, n31870, 
        n31869, n32265, n31868, n31867, n32264, n31866, n31865, 
        n32263, n31864, n31863, n32262, n33811, n31862, n31861, 
        n32261, n33810, n31859, n32260, n33493, n31858, n31857, 
        n32259, n31856, n31855, n32258, n32464, n33492, n31854, 
        n31853, n32257, n31852, n31851, n32256, n32463, n31850, 
        n31849, n32255, n31848, n33382, n32254, n32462, n33491, 
        n33809, n33381, n32253, n31843, n31842, n32252, n32461, 
        n31841, n31840, n33379, n31839, n31838, n32250, n32460, 
        n33490, n31837, n31836, n32249, n31835, n31834, n32248, 
        n32459, n31833, n31832, n32247, n31831, n31830, n32246, 
        n32458, n31829, n33489, n32245, n31827, n31826, n32244, 
        n32457, n31825, n31824, n32243, n31823, n33488, n32242, 
        n32456, n33808, n31821, n31820, n32241, n31819, n31818, 
        n32240, n32455, n31817, n31816, n32239, n31815, n31814, 
        n32238, n32454, n34671, n31813, n31812, n32237, n31811, 
        n31805, n32236, n32453, n33378, n33334, n32235, n31810, 
        n31803, n32234, n34670, n31808, n32233, n31804, n31807, 
        n32232, n33807, n31733, n32231, n34159, n31731, n33806, 
        n33805, n33377, n33804, n31729, n32229, n31727, n32228, 
        n32448, n31725, n32227, n33279, n31723, n32226, n32447, 
        n33376, n33325, n31721, n32225, n31719, n32224, n32446, 
        n34158, n32223, n31700, n33803, n32222, n32445, n31698, 
        n33487, n32221, n31696, n33802, n32220, n32444, n31694, 
        n34157, n32219, n31692, n33801, n32218, n32443, n31690, 
        n33800, n32217, n31688, n32216, n32442, n31686, n34669, 
        n32215, n33278, n33290, n32441, n34156, n34154, n32213, 
        n33799, n33375, n32212, n32440, n33798, n34153, n32211, 
        n33797, n33796, n32210, n32439, n33374, n32209, n33277, 
        n33486, n32208, n32438, n32207, n34152, n33795, n32206, 
        n32437, n33794, n33485, n33793, n34151, n34150, n33792, 
        n33791, n33373, n33790, n32202, n34668, n33276, n32201, 
        n34149, n33484, n31618, n32200, n31616, n32199, n31614, 
        n34148, n32198, n31612, n33789, n32197, n32432, n34667, 
        n31610, n33372, n32196, n31608, n33788, n32195, n32431, 
        n31606, n34147, n32194, n31604, n33787, n32193, n32430, 
        n33786, n31602, n33785, n32192, n31600, n32191, n32429, 
        n31598, n34666, n33275, n31596, n33483, n32189, n32428, 
        n33482, clk_c_enable_2283, n34596, n32188, n34146, n33784, 
        n32187, n32427, n33371, n33782, n32186, n34145, n33781, 
        n32185, n32426, n33780, n34595, n32184, n33322, n32183, 
        n32425, n34579, n32182, n34594, n34144, n33481, n32424, 
        n34665, n33779, n33370, n34664, n33778, n34143, n32178, 
        n32423, n33777, n33776, n32177, n31410, n31400, n32176, 
        n32422, n33775, n34663, n32175, n33274, n31809, n32174, 
        n32421, n31802, n31801, n32173, n31402, n32172, n34662, 
        n34142, n31408, n34661, n32171, n31406, n34660, n32170, 
        n34141, n31404, n34659, n32169, n34140, n33774, n32168, 
        n33369, n33480, n33773, n34139, n32167, n31520, n33772, 
        n33771, n32416, n31518, n33770, n32165, n31516, n34658, 
        n32164, n32415, n33479, n31514, n34657, n32163, n31512, 
        n33273, n32162, n32414, n31510, n33257, n32161, n31508, 
        n34656, n32160, n32413, n33291, n31506, n34655, n32159, 
        n31504, n34138, n32158, n32412, n31502, n33769, n32157, 
        n31500, n33368, n32156, n32411, n33478, n31498, n33768, 
        n32155, n34137, n31471, n32154, n32410, n33767, n31469, 
        n32153, n33766, n31467, n32152, n32409, n33367, n34654, 
        n31465, n32151, n34653, n31463, n33272, n32408, n31461, 
        n32149, n34652, n31459, n32148, n32407, n33477, n34651, 
        n31457, n32147, n34136, n31455, n32146, n32406, n33765, 
        n31453, n32145, n33366, n31451, n32144, n32405, n33476, 
        n33764, n31449, n32143, n34135, n33763, n32142, n33475, 
        n31422, n33762, n32141, n31420, n34650, n32140, n33365, 
        n34593, n31418, n34649, n32139, n31416, n33271, n32138, 
        n31414, n33474, n31412, n34648, n33364, n33472, n34134, 
        n33761, n34133, n33760, n34132, n33759, n34131, n33758, 
        n34130, n33757, n34129, n33756, n34128, n33755, n34127, 
        n33754, n34126, n33753, n34125, n33751, n34123, n33750, 
        n34122, n33749, n34121, n33748, n34120, n33747, n34119, 
        n33746, n34118, n33745, n34117, n33744, n34116, n33743, 
        n34115, n33742, n34114, n33741, n34113, n33740, n34112, 
        n33739, n34111, n33738, n34110, n33737, n34109, n33736, 
        n34108, n33735, n34107, n33734, n34106, n33733, n34105, 
        n33732, n34104, n33731, n34103, n33730, n34102, n33729, 
        n34101, n33728, n34100, n33727, n34099, n33726, n34098, 
        n33725, n34097, n33724, n34096, n33723, n34095, n33722, 
        n34094, n33720, n34092, n33719, n34091, n33718, n34090, 
        n33717, n34089, n33471, n33470, n33716, n33363, n34647, 
        n33362, n34842, n33469, n33715, n33361, n34088, n34592, 
        n33338, n34532, n33360, n34087, n33359, n33714, n33468, 
        n33713, n33712, n34086, n33467, n34591, n33358, n33357, 
        n34085, n34646, n33711, n34645, n33710, n33709, n33708, 
        n34084, n34083, n33356, n34644, n33355, n34643, n33337, 
        n33707, n33706, n34642, n34590, n33466, n34082, n33354, 
        n33465, n33353, n33464, n34641, n33352, n34640, n33463, 
        n33351, n33350, n34081, n33462, n33705, n33704, n33336, 
        n34639, n33461, n34638, n33703, n34080, n34637, n34079, 
        n34636, n34635, n34078, n34634, n33702, n33701, n33700, 
        n33348, n33347, n34077, n33346, n33460, n34633, n33335, 
        n33459, n33458, n33345, n34632;
    
    VHI i2 (.Z(VCC_net));
    LUT4 i15227_3_lut (.A(\result_i[26] [6]), .B(\result_i[27] [6]), .C(y_1_delay[0]), 
         .Z(n33611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15227_3_lut.init = 16'hcaca;
    LUT4 i15032_3_lut (.A(\result_i[8] [12]), .B(\result_i[9] [12]), .C(y_1_delay[0]), 
         .Z(n33416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15032_3_lut.init = 16'hcaca;
    PFUMX i15604 (.BLUT(n33974), .ALUT(n33975), .C0(y_1_delay[1]), .Z(n33988));
    PFUMX i14955 (.BLUT(n33327), .ALUT(n33328), .C0(y_1_delay[1]), .Z(n33339));
    LUT4 i15135_3_lut (.A(\result_i[28] [9]), .B(\result_i[29] [9]), .C(y_1_delay[0]), 
         .Z(n33519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15135_3_lut.init = 16'hcaca;
    CCU2C _add_1_1110_add_4_18 (.A0(shift_2_dout_i[15]), .B0(shift_2_dout_r[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[16]), .B1(shift_2_dout_r[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32116), .COUT(n32117), .S0(n12167), 
          .S1(n12168));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_18.INJECT1_1 = "NO";
    LUT4 i2831_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[468])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2831_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1110_add_4_16 (.A0(shift_2_dout_i[13]), .B0(shift_2_dout_r[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[14]), .B1(shift_2_dout_r[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32115), .COUT(n32116), .S0(n12165), 
          .S1(n12166));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_16.INJECT1_1 = "NO";
    LUT4 i2823_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[469])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2823_3_lut_4_lut.init = 16'hf2d0;
    FD1P3AX result_i_31___i1 (.D(result_i_ns_0__15__N_517[0]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i1.GSR = "ENABLED";
    PFUMX i15423 (.BLUT(n33798), .ALUT(n33799), .C0(y_1_delay[1]), .Z(n33807));
    FD1S3AX in_valid_reg_48 (.D(in_valid_c), .CK(clk_c), .Q(in_valid_reg));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam in_valid_reg_48.GSR = "ENABLED";
    FD1S3AX r4_valid_50 (.D(clk_c_enable_2300), .CK(clk_c), .Q(r4_valid));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam r4_valid_50.GSR = "ENABLED";
    FD1S3AX assign_out_52 (.D(next_out_valid), .CK(clk_c), .Q(out_valid_c));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam assign_out_52.GSR = "ENABLED";
    LUT4 i2815_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[470])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2815_3_lut_4_lut.init = 16'hf2d0;
    FD1S3AX y_1_delay_i0 (.D(n34740), .CK(clk_c), .Q(y_1_delay[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam y_1_delay_i0.GSR = "ENABLED";
    FD1S3AX din_r_reg_i1 (.D(din_r_c_0), .CK(clk_c), .Q(din_r_reg[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i1.GSR = "ENABLED";
    PFUMX i15605 (.BLUT(n33976), .ALUT(n33977), .C0(y_1_delay[1]), .Z(n33989));
    FD1P3AX result_i_31___i86 (.D(result_i_ns_0__15__N_517[85]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i86.GSR = "ENABLED";
    LUT4 i2807_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[471])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2807_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15733 (.BLUT(n34108), .ALUT(n34109), .C0(y_1_delay[1]), .Z(n34117));
    LUT4 i2799_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[472])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2799_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i14956 (.BLUT(n33329), .ALUT(n33330), .C0(y_1_delay[1]), .Z(n33340));
    LUT4 i2791_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[473])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2791_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15031_3_lut (.A(\result_i[6] [12]), .B(\result_i[7] [12]), .C(y_1_delay[0]), 
         .Z(n33415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15031_3_lut.init = 16'hcaca;
    CCU2C _add_1_1078_add_4_13 (.A0(shift_1_dout_i[11]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[11]), .A1(shift_1_dout_i[12]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[12]), .CIN(n31971), 
          .COUT(n31972), .S0(op_i_23__N_1154_adj_7482[11]), .S1(op_i_23__N_1154_adj_7482[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_13.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_13.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_13.INJECT1_1 = "NO";
    LUT4 i2783_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[474])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2783_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15291_3_lut (.A(\result_i[30] [4]), .B(\result_i[31] [4]), .C(y_1_delay[0]), 
         .Z(n33675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15291_3_lut.init = 16'hcaca;
    LUT4 i6737_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[491])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6737_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2775_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[475])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2775_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15107 (.BLUT(n33476), .ALUT(n33477), .C0(y_1_delay[1]), .Z(n33491));
    LUT4 i6729_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[492])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6729_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2767_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[476])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2767_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15226_3_lut (.A(\result_i[24] [6]), .B(\result_i[25] [6]), .C(y_1_delay[0]), 
         .Z(n33610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15226_3_lut.init = 16'hcaca;
    LUT4 i2759_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[477])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2759_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2751_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[478])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2751_3_lut_4_lut.init = 16'hf2d0;
    FD1P3AX result_i_31___i85 (.D(result_i_ns_0__15__N_517[84]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i85.GSR = "ENABLED";
    PFUMX i14957 (.BLUT(n33331), .ALUT(n33332), .C0(y_1_delay[1]), .Z(n33341));
    LUT4 i2743_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[479])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2743_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6953_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[464])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6953_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6945_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[465])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6945_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6937_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[466])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6937_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15030_3_lut (.A(\result_i[4] [12]), .B(\result_i[5] [12]), .C(y_1_delay[0]), 
         .Z(n33414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15030_3_lut.init = 16'hcaca;
    LUT4 i6721_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[493])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6721_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6713_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[494])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6713_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15033_3_lut (.A(\result_i[10] [12]), .B(\result_i[11] [12]), .C(y_1_delay[0]), 
         .Z(n33417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15033_3_lut.init = 16'hcaca;
    LUT4 i6929_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[467])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6929_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6921_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[468])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6921_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6705_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[495])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6705_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2863_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[464])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2863_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15108 (.BLUT(n33478), .ALUT(n33479), .C0(y_1_delay[1]), .Z(n33492));
    PFUMX i15606 (.BLUT(n33978), .ALUT(n33979), .C0(y_1_delay[1]), .Z(n33990));
    LUT4 i6913_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[469])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6913_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6905_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[470])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6905_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6897_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[471])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6897_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2855_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[465])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2855_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2847_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[466])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2847_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2839_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[2] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[467])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2839_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6889_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[472])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6889_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15225_3_lut (.A(\result_i[22] [6]), .B(\result_i[23] [6]), .C(y_1_delay[0]), 
         .Z(n33609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15225_3_lut.init = 16'hcaca;
    LUT4 i6881_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[473])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6881_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6873_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[474])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6873_3_lut_4_lut.init = 16'hf2d0;
    FD1P3AX result_i_31___i84 (.D(result_i_ns_0__15__N_517[83]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i84.GSR = "ENABLED";
    FD1P3AX result_i_31___i83 (.D(result_i_ns_0__15__N_517[82]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i83.GSR = "ENABLED";
    LUT4 i6865_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[475])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6865_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15109 (.BLUT(n33480), .ALUT(n33481), .C0(y_1_delay[1]), .Z(n33493));
    LUT4 i6857_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[476])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6857_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15607 (.BLUT(n33980), .ALUT(n33981), .C0(y_1_delay[1]), .Z(n33991));
    LUT4 i6849_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[477])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6849_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15224_3_lut (.A(\result_i[20] [6]), .B(\result_i[21] [6]), .C(y_1_delay[0]), 
         .Z(n33608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15224_3_lut.init = 16'hcaca;
    LUT4 i6841_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[478])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6841_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6833_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[2] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[479])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6833_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2992_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[448])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2992_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15110 (.BLUT(n33482), .ALUT(n33483), .C0(y_1_delay[1]), .Z(n33494));
    PFUMX i15237 (.BLUT(n33612), .ALUT(n33613), .C0(y_1_delay[1]), .Z(n33621));
    LUT4 i2984_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[449])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2984_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15223_3_lut (.A(\result_i[18] [6]), .B(\result_i[19] [6]), .C(y_1_delay[0]), 
         .Z(n33607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15223_3_lut.init = 16'hcaca;
    LUT4 i2976_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[450])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2976_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i14958 (.BLUT(n33333), .ALUT(n33334), .C0(y_1_delay[1]), .Z(n33342));
    FD1P3AX result_i_31___i82 (.D(result_i_ns_0__15__N_517[81]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i82.GSR = "ENABLED";
    LUT4 i2968_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[451])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2968_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15222_3_lut (.A(\result_i[16] [6]), .B(\result_i[17] [6]), .C(y_1_delay[0]), 
         .Z(n33606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15222_3_lut.init = 16'hcaca;
    CCU2C _add_1_1078_add_4_11 (.A0(shift_1_dout_i[9]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[9]), .A1(shift_1_dout_i[10]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[10]), .CIN(n31970), 
          .COUT(n31971), .S0(op_i_23__N_1154_adj_7482[9]), .S1(op_i_23__N_1154_adj_7482[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_11.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_11.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_11.INJECT1_1 = "NO";
    OB dout_r_pad_5 (.I(dout_r_c_5), .O(dout_r[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    LUT4 i2960_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[452])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2960_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2952_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[453])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2952_3_lut_4_lut.init = 16'hf1e0;
    OB dout_r_pad_6 (.I(dout_r_c_6), .O(dout_r[6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    LUT4 i2944_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[454])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2944_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15111 (.BLUT(n33484), .ALUT(n33485), .C0(y_1_delay[1]), .Z(n33495));
    LUT4 i15589_3_lut (.A(\result_r[6] [9]), .B(\result_r[7] [9]), .C(y_1_delay[0]), 
         .Z(n33973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15589_3_lut.init = 16'hcaca;
    LUT4 i15588_3_lut (.A(\result_r[4] [9]), .B(\result_r[5] [9]), .C(y_1_delay[0]), 
         .Z(n33972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15588_3_lut.init = 16'hcaca;
    OB dout_r_pad_7 (.I(dout_r_c_7), .O(dout_r[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    LUT4 i2936_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[455])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2936_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i14954 (.BLUT(n33325), .ALUT(n33326), .C0(y_1_delay[1]), .Z(n33338));
    PFUMX i15665 (.BLUT(n34034), .ALUT(n34035), .C0(y_1_delay[1]), .Z(n34049));
    PFUMX i15112 (.BLUT(n33486), .ALUT(n33487), .C0(y_1_delay[1]), .Z(n33496));
    CCU2C _add_1_1078_add_4_9 (.A0(shift_1_dout_i[7]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[7]), .A1(shift_1_dout_i[8]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[8]), .CIN(n31969), 
          .COUT(n31970), .S1(op_i_23__N_1154_adj_7482[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_9.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_9.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_9.INJECT1_1 = "NO";
    PFUMX i15416 (.BLUT(n33784), .ALUT(n33785), .C0(y_1_delay[1]), .Z(n33800));
    PFUMX i15417 (.BLUT(n33786), .ALUT(n33787), .C0(y_1_delay[1]), .Z(n33801));
    CCU2C _add_1_1078_add_4_7 (.A0(shift_1_dout_i[5]), .B0(n34769), .C0(count_adj_7456[1]), 
          .D0(op_i_23__N_1154_adj_7426[5]), .A1(shift_1_dout_i[6]), .B1(n34769), 
          .C1(count_adj_7456[1]), .D1(op_i_23__N_1154_adj_7426[6]), .CIN(n31968), 
          .COUT(n31969));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_7.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_7.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_7.INJECT1_1 = "NO";
    PFUMX i15013 (.BLUT(n33381), .ALUT(n33382), .C0(y_1_delay[1]), .Z(n33397));
    PFUMX i15730 (.BLUT(n34102), .ALUT(n34103), .C0(y_1_delay[1]), .Z(n34114));
    PFUMX i15014 (.BLUT(n33383), .ALUT(n33384), .C0(y_1_delay[1]), .Z(n33398));
    PFUMX i15015 (.BLUT(n33385), .ALUT(n33386), .C0(y_1_delay[1]), .Z(n33399));
    LUT4 i15587_3_lut (.A(\result_r[2] [9]), .B(\result_r[3] [9]), .C(y_1_delay[0]), 
         .Z(n33971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15587_3_lut.init = 16'hcaca;
    PFUMX i15016 (.BLUT(n33387), .ALUT(n33388), .C0(y_1_delay[1]), .Z(n33400));
    CCU2C _add_1_1078_add_4_5 (.A0(shift_1_dout_i[3]), .B0(n34769), .C0(count_adj_7456[1]), 
          .D0(op_i_23__N_1154_adj_7426[3]), .A1(shift_1_dout_i[4]), .B1(n34769), 
          .C1(count_adj_7456[1]), .D1(op_i_23__N_1154_adj_7426[4]), .CIN(n31967), 
          .COUT(n31968));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_5.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_5.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_5.INJECT1_1 = "NO";
    PFUMX i15418 (.BLUT(n33788), .ALUT(n33789), .C0(y_1_delay[1]), .Z(n33802));
    CCU2C _add_1_1078_add_4_3 (.A0(shift_1_dout_i[1]), .B0(n34769), .C0(count_adj_7456[1]), 
          .D0(op_i_23__N_1154_adj_7426[1]), .A1(shift_1_dout_i[2]), .B1(n34769), 
          .C1(count_adj_7456[1]), .D1(op_i_23__N_1154_adj_7426[2]), .CIN(n31966), 
          .COUT(n31967));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_3.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_3.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_3.INJECT1_1 = "NO";
    LUT4 i2928_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[456])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2928_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15586_3_lut (.A(\result_r[0] [9]), .B(\result_r[1] [9]), .C(y_1_delay[0]), 
         .Z(n33970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15586_3_lut.init = 16'hcaca;
    LUT4 i2920_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[457])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2920_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2912_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[458])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2912_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15221_3_lut (.A(\result_i[14] [6]), .B(\result_i[15] [6]), .C(y_1_delay[0]), 
         .Z(n33605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15221_3_lut.init = 16'hcaca;
    LUT4 i2904_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[459])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2904_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15220_3_lut (.A(\result_i[12] [6]), .B(\result_i[13] [6]), .C(y_1_delay[0]), 
         .Z(n33604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15220_3_lut.init = 16'hcaca;
    LUT4 i2896_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[460])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2896_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2888_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[461])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2888_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15017 (.BLUT(n33389), .ALUT(n33390), .C0(y_1_delay[1]), .Z(n33401));
    LUT4 i15029_3_lut (.A(\result_i[2] [12]), .B(\result_i[3] [12]), .C(y_1_delay[0]), 
         .Z(n33413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15029_3_lut.init = 16'hcaca;
    PFUMX i15419 (.BLUT(n33790), .ALUT(n33791), .C0(y_1_delay[1]), .Z(n33803));
    PFUMX i15420 (.BLUT(n33792), .ALUT(n33793), .C0(y_1_delay[1]), .Z(n33804));
    LUT4 i2880_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[462])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2880_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15447 (.BLUT(n33815), .ALUT(n33816), .C0(y_1_delay[1]), .Z(n33831));
    LUT4 i15028_3_lut (.A(\result_i[0] [12]), .B(\result_i[1] [12]), .C(y_1_delay[0]), 
         .Z(n33412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15028_3_lut.init = 16'hcaca;
    LUT4 i2872_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_i[3] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[463])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2872_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7081_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[448])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7081_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15608 (.BLUT(n33982), .ALUT(n33983), .C0(y_1_delay[1]), .Z(n33992));
    LUT4 i15219_3_lut (.A(\result_i[10] [6]), .B(\result_i[11] [6]), .C(y_1_delay[0]), 
         .Z(n33603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15219_3_lut.init = 16'hcaca;
    LUT4 i7073_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[449])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7073_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15218_3_lut (.A(\result_i[8] [6]), .B(\result_i[9] [6]), .C(y_1_delay[0]), 
         .Z(n33602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15218_3_lut.init = 16'hcaca;
    LUT4 i7065_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[450])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7065_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15731 (.BLUT(n34104), .ALUT(n34105), .C0(y_1_delay[1]), .Z(n34115));
    PFUMX i15018 (.BLUT(n33391), .ALUT(n33392), .C0(y_1_delay[1]), .Z(n33402));
    PFUMX i15421 (.BLUT(n33794), .ALUT(n33795), .C0(y_1_delay[1]), .Z(n33805));
    PFUMX i15732 (.BLUT(n34106), .ALUT(n34107), .C0(y_1_delay[1]), .Z(n34116));
    PFUMX i15422 (.BLUT(n33796), .ALUT(n33797), .C0(y_1_delay[1]), .Z(n33806));
    PFUMX i15019 (.BLUT(n33393), .ALUT(n33394), .C0(y_1_delay[1]), .Z(n33403));
    PFUMX i15106 (.BLUT(n33474), .ALUT(n33475), .C0(y_1_delay[1]), .Z(n33490));
    FD1P3AX result_i_31___i81 (.D(result_i_ns_0__15__N_517[80]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i81.GSR = "ENABLED";
    PFUMX i15113 (.BLUT(n33488), .ALUT(n33489), .C0(y_1_delay[1]), .Z(n33497));
    LUT4 i12103_1_lut (.A(over), .Z(clk_c_enable_2259)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam i12103_1_lut.init = 16'h5555;
    LUT4 i15217_3_lut (.A(\result_i[6] [6]), .B(\result_i[7] [6]), .C(y_1_delay[0]), 
         .Z(n33601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15217_3_lut.init = 16'hcaca;
    LUT4 i15216_3_lut (.A(\result_i[4] [6]), .B(\result_i[5] [6]), .C(y_1_delay[0]), 
         .Z(n33600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15216_3_lut.init = 16'hcaca;
    LUT4 i15215_3_lut (.A(\result_i[2] [6]), .B(\result_i[3] [6]), .C(y_1_delay[0]), 
         .Z(n33599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15215_3_lut.init = 16'hcaca;
    LUT4 i12103_1_lut_rep_448 (.A(over), .Z(clk_c_enable_2283)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam i12103_1_lut_rep_448.init = 16'h5555;
    LUT4 i15214_3_lut (.A(\result_i[0] [6]), .B(\result_i[1] [6]), .C(y_1_delay[0]), 
         .Z(n33598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15214_3_lut.init = 16'hcaca;
    PFUMX i15609 (.BLUT(n33984), .ALUT(n33985), .C0(y_1_delay[1]), .Z(n33993));
    PFUMX i15448 (.BLUT(n33817), .ALUT(n33818), .C0(y_1_delay[1]), .Z(n33832));
    FD1P3AX result_i_31___i80 (.D(result_i_ns_0__15__N_517[79]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i80.GSR = "ENABLED";
    FD1P3AX result_i_31___i79 (.D(result_i_ns_0__15__N_517[78]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i79.GSR = "ENABLED";
    FD1P3AX result_i_31___i78 (.D(result_i_ns_0__15__N_517[77]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i78.GSR = "ENABLED";
    FD1P3AX result_i_31___i77 (.D(result_i_ns_0__15__N_517[76]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i77.GSR = "ENABLED";
    FD1P3AX result_i_31___i76 (.D(result_i_ns_0__15__N_517[75]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i76.GSR = "ENABLED";
    FD1P3AX result_i_31___i75 (.D(result_i_ns_0__15__N_517[74]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i75.GSR = "ENABLED";
    FD1P3AX result_i_31___i74 (.D(result_i_ns_0__15__N_517[73]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i74.GSR = "ENABLED";
    FD1P3AX result_i_31___i73 (.D(result_i_ns_0__15__N_517[72]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i73.GSR = "ENABLED";
    FD1P3AX result_i_31___i72 (.D(result_i_ns_0__15__N_517[71]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i72.GSR = "ENABLED";
    FD1P3AX result_i_31___i71 (.D(result_i_ns_0__15__N_517[70]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i71.GSR = "ENABLED";
    FD1P3AX result_i_31___i70 (.D(result_i_ns_0__15__N_517[69]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i70.GSR = "ENABLED";
    FD1P3AX result_i_31___i69 (.D(result_i_ns_0__15__N_517[68]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i69.GSR = "ENABLED";
    FD1P3AX result_i_31___i68 (.D(result_i_ns_0__15__N_517[67]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i68.GSR = "ENABLED";
    FD1P3AX result_i_31___i67 (.D(result_i_ns_0__15__N_517[66]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i67.GSR = "ENABLED";
    FD1P3AX result_i_31___i66 (.D(result_i_ns_0__15__N_517[65]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i66.GSR = "ENABLED";
    FD1P3AX over_53 (.D(VCC_net), .SP(next_over_N_1081), .CK(clk_c), .Q(over));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam over_53.GSR = "ENABLED";
    LUT4 i15570_3_lut (.A(\result_r[30] [10]), .B(\result_r[31] [10]), .C(y_1_delay[0]), 
         .Z(n33954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15570_3_lut.init = 16'hcaca;
    LUT4 i7057_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[451])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7057_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15569_3_lut (.A(\result_r[28] [10]), .B(\result_r[29] [10]), .C(y_1_delay[0]), 
         .Z(n33953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15569_3_lut.init = 16'hcaca;
    PFUMX i15020 (.BLUT(n33395), .ALUT(n33396), .C0(y_1_delay[1]), .Z(n33404));
    PFUMX i15047 (.BLUT(n33418), .ALUT(n33419), .C0(y_1_delay[1]), .Z(n33431));
    PFUMX i15449 (.BLUT(n33819), .ALUT(n33820), .C0(y_1_delay[1]), .Z(n33833));
    LUT4 i15568_3_lut (.A(\result_r[26] [10]), .B(\result_r[27] [10]), .C(y_1_delay[0]), 
         .Z(n33952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15568_3_lut.init = 16'hcaca;
    LUT4 i15567_3_lut (.A(\result_r[24] [10]), .B(\result_r[25] [10]), .C(y_1_delay[0]), 
         .Z(n33951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15567_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(count_y[1]), .B(count_y[4]), .C(count_y[2]), .D(count_y[5]), 
         .Z(n32925)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hfffe;
    PFUMX i15450 (.BLUT(n33821), .ALUT(n33822), .C0(y_1_delay[1]), .Z(n33834));
    LUT4 i15566_3_lut (.A(\result_r[22] [10]), .B(\result_r[23] [10]), .C(y_1_delay[0]), 
         .Z(n33950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15566_3_lut.init = 16'hcaca;
    PFUMX i15048 (.BLUT(n33420), .ALUT(n33421), .C0(y_1_delay[1]), .Z(n33432));
    LUT4 i15565_3_lut (.A(\result_r[20] [10]), .B(\result_r[21] [10]), .C(y_1_delay[0]), 
         .Z(n33949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15565_3_lut.init = 16'hcaca;
    PFUMX i15451 (.BLUT(n33823), .ALUT(n33824), .C0(y_1_delay[1]), .Z(n33835));
    LUT4 i15564_3_lut (.A(\result_r[18] [10]), .B(\result_r[19] [10]), .C(y_1_delay[0]), 
         .Z(n33948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15564_3_lut.init = 16'hcaca;
    LUT4 i15563_3_lut (.A(\result_r[16] [10]), .B(\result_r[17] [10]), .C(y_1_delay[0]), 
         .Z(n33947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15563_3_lut.init = 16'hcaca;
    CCU2C _add_1_1110_add_4_14 (.A0(shift_2_dout_i[11]), .B0(shift_2_dout_r[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[12]), .B1(shift_2_dout_r[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32114), .COUT(n32115), .S0(n12163), 
          .S1(n12164));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_12 (.A0(shift_2_dout_i[9]), .B0(shift_2_dout_r[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[10]), .B1(shift_2_dout_r[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32113), .COUT(n32114), .S0(n12161), 
          .S1(n12162));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_10 (.A0(shift_2_dout_i[7]), .B0(shift_2_dout_r[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[8]), .B1(shift_2_dout_r[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32112), .COUT(n32113), .S0(n12159), 
          .S1(n12160));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_8 (.A0(shift_2_dout_i[5]), .B0(shift_2_dout_r[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[6]), .B1(shift_2_dout_r[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32111), .COUT(n32112), .S0(n12157), 
          .S1(n12158));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_6 (.A0(shift_2_dout_i[3]), .B0(shift_2_dout_r[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[4]), .B1(shift_2_dout_r[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32110), .COUT(n32111), .S0(n12155), 
          .S1(n12156));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_4 (.A0(shift_2_dout_i[1]), .B0(shift_2_dout_r[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[2]), .B1(shift_2_dout_r[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32109), .COUT(n32110), .S0(n12153), 
          .S1(n12154));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(shift_2_dout_i[0]), .B1(shift_2_dout_r[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32109), .S1(n12152));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1110_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_26 (.A0(shift_8_dout_i[23]), .B0(shift_8_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n32108), .S0(n319_adj_6495));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1048_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_24 (.A0(shift_8_dout_i[22]), .B0(shift_8_dout_r[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[23]), .B1(shift_8_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32107), .COUT(n32108), .S0(n11170), 
          .S1(n11171));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_22 (.A0(shift_8_dout_i[20]), .B0(shift_8_dout_r[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[21]), .B1(shift_8_dout_r[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32106), .COUT(n32107), .S0(n11168), 
          .S1(n11169));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_20 (.A0(shift_8_dout_i[18]), .B0(shift_8_dout_r[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[19]), .B1(shift_8_dout_r[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32105), .COUT(n32106), .S0(n11166), 
          .S1(n11167));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_18 (.A0(shift_8_dout_i[16]), .B0(shift_8_dout_r[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[17]), .B1(shift_8_dout_r[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32104), .COUT(n32105), .S0(n11164), 
          .S1(n11165));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_16 (.A0(shift_8_dout_i[14]), .B0(shift_8_dout_r[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[15]), .B1(shift_8_dout_r[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32103), .COUT(n32104), .S0(n11162), 
          .S1(n11163));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_14 (.A0(shift_8_dout_i[12]), .B0(shift_8_dout_r[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[13]), .B1(shift_8_dout_r[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32102), .COUT(n32103), .S0(n11160), 
          .S1(n11161));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_12 (.A0(shift_8_dout_i[10]), .B0(shift_8_dout_r[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[11]), .B1(shift_8_dout_r[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32101), .COUT(n32102), .S0(n11158), 
          .S1(n11159));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_10 (.A0(shift_8_dout_i[8]), .B0(shift_8_dout_r[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[9]), .B1(shift_8_dout_r[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32100), .COUT(n32101), .S0(n11156), 
          .S1(n11157));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_8 (.A0(shift_8_dout_i[6]), .B0(shift_8_dout_r[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[7]), .B1(shift_8_dout_r[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32099), .COUT(n32100), .S0(n11154), 
          .S1(n11155));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_6 (.A0(shift_8_dout_i[4]), .B0(shift_8_dout_r[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[5]), .B1(shift_8_dout_r[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32098), .COUT(n32099), .S0(n11152), 
          .S1(n11153));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_4 (.A0(shift_8_dout_i[2]), .B0(shift_8_dout_r[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[3]), .B1(shift_8_dout_r[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32097), .COUT(n32098), .S0(n11150), 
          .S1(n11151));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1048_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1048_add_4_2 (.A0(shift_8_dout_i[0]), .B0(shift_8_dout_r[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[1]), .B1(shift_8_dout_r[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32097), .S1(n11149));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1048_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1048_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1048_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1048_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_32 (.A0(op_r_23__N_1268[30]), .B0(op_i_23__N_1310[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[31]), .B1(op_i_23__N_1310[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32094), .S0(op_i_23__N_1130[30]), 
          .S1(op_i_23__N_1130[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_30 (.A0(op_r_23__N_1268[28]), .B0(op_i_23__N_1310[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[29]), .B1(op_i_23__N_1310[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32093), .COUT(n32094), .S0(op_i_23__N_1130[28]), 
          .S1(op_i_23__N_1130[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_28 (.A0(op_r_23__N_1268[26]), .B0(op_i_23__N_1310[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[27]), .B1(op_i_23__N_1310[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32092), .COUT(n32093), .S0(op_i_23__N_1130[26]), 
          .S1(op_i_23__N_1130[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_26 (.A0(op_r_23__N_1268[24]), .B0(op_i_23__N_1310[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[25]), .B1(op_i_23__N_1310[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32091), .COUT(n32092), .S0(op_i_23__N_1130[24]), 
          .S1(op_i_23__N_1130[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_24 (.A0(op_r_23__N_1268[22]), .B0(op_i_23__N_1310[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[23]), .B1(op_i_23__N_1310[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32090), .COUT(n32091), .S0(op_i_23__N_1130[22]), 
          .S1(op_i_23__N_1130[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_22 (.A0(op_r_23__N_1268[20]), .B0(op_i_23__N_1310[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[21]), .B1(op_i_23__N_1310[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32089), .COUT(n32090), .S0(op_i_23__N_1130[20]), 
          .S1(op_i_23__N_1130[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_20 (.A0(op_r_23__N_1268[18]), .B0(op_i_23__N_1310[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[19]), .B1(op_i_23__N_1310[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32088), .COUT(n32089), .S0(op_i_23__N_1130[18]), 
          .S1(op_i_23__N_1130[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_18 (.A0(op_r_23__N_1268[16]), .B0(op_i_23__N_1310[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[17]), .B1(op_i_23__N_1310[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32087), .COUT(n32088), .S0(op_i_23__N_1130[16]), 
          .S1(op_i_23__N_1130[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_16 (.A0(op_r_23__N_1268[14]), .B0(op_i_23__N_1310[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[15]), .B1(op_i_23__N_1310[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32086), .COUT(n32087), .S0(op_i_23__N_1130[14]), 
          .S1(op_i_23__N_1130[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_16.INJECT1_1 = "NO";
    LUT4 i15562_3_lut (.A(\result_r[14] [10]), .B(\result_r[15] [10]), .C(y_1_delay[0]), 
         .Z(n33946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15562_3_lut.init = 16'hcaca;
    PFUMX i15452 (.BLUT(n33825), .ALUT(n33826), .C0(y_1_delay[1]), .Z(n33836));
    LUT4 i15561_3_lut (.A(\result_r[12] [10]), .B(\result_r[13] [10]), .C(y_1_delay[0]), 
         .Z(n33945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15561_3_lut.init = 16'hcaca;
    LUT4 i15560_3_lut (.A(\result_r[10] [10]), .B(\result_r[11] [10]), .C(y_1_delay[0]), 
         .Z(n33944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15560_3_lut.init = 16'hcaca;
    LUT4 i12448_2_lut (.A(out_valid_c), .B(over), .Z(next_out_valid)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(309[10:38])
    defparam i12448_2_lut.init = 16'heeee;
    LUT4 i15559_3_lut (.A(\result_r[8] [10]), .B(\result_r[9] [10]), .C(y_1_delay[0]), 
         .Z(n33943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15559_3_lut.init = 16'hcaca;
    LUT4 i15849_3_lut (.A(\result_r[30] [1]), .B(\result_r[31] [1]), .C(y_1_delay[0]), 
         .Z(n34233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15849_3_lut.init = 16'hcaca;
    LUT4 i15848_3_lut (.A(\result_r[28] [1]), .B(\result_r[29] [1]), .C(y_1_delay[0]), 
         .Z(n34232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15848_3_lut.init = 16'hcaca;
    LUT4 i15558_3_lut (.A(\result_r[6] [10]), .B(\result_r[7] [10]), .C(y_1_delay[0]), 
         .Z(n33942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15558_3_lut.init = 16'hcaca;
    LUT4 i7049_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[452])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7049_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15049 (.BLUT(n33422), .ALUT(n33423), .C0(y_1_delay[1]), .Z(n33433));
    PFUMX i15453 (.BLUT(n33827), .ALUT(n33828), .C0(y_1_delay[1]), .Z(n33837));
    PFUMX i15050 (.BLUT(n33424), .ALUT(n33425), .C0(y_1_delay[1]), .Z(n33434));
    LUT4 i15290_3_lut (.A(\result_i[28] [4]), .B(\result_i[29] [4]), .C(y_1_delay[0]), 
         .Z(n33674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15290_3_lut.init = 16'hcaca;
    PFUMX i15454 (.BLUT(n33829), .ALUT(n33830), .C0(y_1_delay[1]), .Z(n33838));
    PFUMX i15137 (.BLUT(n33505), .ALUT(n33506), .C0(y_1_delay[1]), .Z(n33521));
    LUT4 i15557_3_lut (.A(\result_r[4] [10]), .B(\result_r[5] [10]), .C(y_1_delay[0]), 
         .Z(n33941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15557_3_lut.init = 16'hcaca;
    LUT4 i7041_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[453])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7041_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7033_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[454])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7033_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15556_3_lut (.A(\result_r[2] [10]), .B(\result_r[3] [10]), .C(y_1_delay[0]), 
         .Z(n33940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15556_3_lut.init = 16'hcaca;
    FD1S3AX s5_count_49 (.D(n19995), .CK(clk_c), .Q(s5_count));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam s5_count_49.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i1 (.D(next_dout_i_15__N_1045[0]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_0));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i1.GSR = "ENABLED";
    LUT4 i15555_3_lut (.A(\result_r[0] [10]), .B(\result_r[1] [10]), .C(y_1_delay[0]), 
         .Z(n33939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15555_3_lut.init = 16'hcaca;
    PFUMX i15168 (.BLUT(n33536), .ALUT(n33537), .C0(y_1_delay[1]), .Z(n33552));
    LUT4 i7025_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[455])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7025_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1078_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(shift_1_dout_i[0]), .B1(n34769), .C1(count_adj_7456[1]), 
          .D1(op_i_23__N_1154_adj_7426[0]), .COUT(n31966));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1078_add_4_1.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_1.INJECT1_1 = "NO";
    LUT4 i15289_3_lut (.A(\result_i[26] [4]), .B(\result_i[27] [4]), .C(y_1_delay[0]), 
         .Z(n33673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15289_3_lut.init = 16'hcaca;
    LUT4 i7017_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[456])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7017_3_lut_4_lut.init = 16'hf1e0;
    OB dout_r_pad_8 (.I(dout_r_c_8), .O(dout_r[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    LUT4 i15847_3_lut (.A(\result_r[26] [1]), .B(\result_r[27] [1]), .C(y_1_delay[0]), 
         .Z(n34231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15847_3_lut.init = 16'hcaca;
    PFUMX i15169 (.BLUT(n33538), .ALUT(n33539), .C0(y_1_delay[1]), .Z(n33553));
    OB dout_r_pad_9 (.I(dout_r_c_9), .O(dout_r[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_10 (.I(dout_r_c_10), .O(dout_r[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_11 (.I(dout_r_c_11), .O(dout_r[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_12 (.I(dout_r_c_12), .O(dout_r[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    PFUMX i15051 (.BLUT(n33426), .ALUT(n33427), .C0(y_1_delay[1]), .Z(n33435));
    PFUMX i15757 (.BLUT(n34125), .ALUT(n34126), .C0(y_1_delay[1]), .Z(n34141));
    LUT4 i15846_3_lut (.A(\result_r[24] [1]), .B(\result_r[25] [1]), .C(y_1_delay[0]), 
         .Z(n34230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15846_3_lut.init = 16'hcaca;
    LUT4 i7009_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[457])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7009_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15288_3_lut (.A(\result_i[24] [4]), .B(\result_i[25] [4]), .C(y_1_delay[0]), 
         .Z(n33672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15288_3_lut.init = 16'hcaca;
    FD1P3AX result_r_31___i1 (.D(result_r_ns_0__15__N_3[0]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i1.GSR = "ENABLED";
    LUT4 i7001_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[458])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7001_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6993_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[459])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6993_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6985_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[460])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6985_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15649_3_lut (.A(\result_r[2] [7]), .B(\result_r[3] [7]), .C(y_1_delay[0]), 
         .Z(n34033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15649_3_lut.init = 16'hcaca;
    PFUMX i15138 (.BLUT(n33507), .ALUT(n33508), .C0(y_1_delay[1]), .Z(n33522));
    FD1P3AX result_i_31___i65 (.D(result_i_ns_0__15__N_517[64]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[27] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i65.GSR = "ENABLED";
    CCU2C _add_1_1031_add_4_25 (.A0(n31476), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[22]), .A1(n31474), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[23]), .CIN(n31964), .S0(op_i_23__N_1154_adj_7371[22]), 
          .S1(op_i_23__N_1154_adj_7371[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_25.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_25.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_25.INJECT1_1 = "NO";
    FD1P3AX dout_r_i0_i1 (.D(next_dout_r_15__N_1029[0]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_0));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_1031_add_4_23 (.A0(n31480), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[20]), .A1(n31478), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[21]), .CIN(n31963), .COUT(n31964), .S0(op_i_23__N_1154_adj_7371[20]), 
          .S1(op_i_23__N_1154_adj_7371[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_23.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_23.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_23.INJECT1_1 = "NO";
    LUT4 i6977_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[461])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6977_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15170 (.BLUT(n33540), .ALUT(n33541), .C0(y_1_delay[1]), .Z(n33554));
    LUT4 r4_valid_I_0_65_2_lut (.A(r4_valid), .B(s5_count), .Z(no5_state[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(247[8:36])
    defparam r4_valid_I_0_65_2_lut.init = 16'h2222;
    LUT4 i6969_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[462])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6969_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6961_3_lut_4_lut (.A(n34716), .B(n34704), .C(\result_r[3] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[463])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6961_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14081_2_lut (.A(shift_1_dout_i[0]), .B(shift_1_dout_r[0]), .Z(n11556)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14081_2_lut.init = 16'h6666;
    LUT4 i3120_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[432])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14068_2_lut (.A(op_i_23__N_1154[0]), .B(op_r_23__N_1106[0]), .Z(n9983)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14068_2_lut.init = 16'h6666;
    LUT4 i3112_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[433])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3112_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15633 (.BLUT(n34001), .ALUT(n34002), .C0(y_1_delay[1]), .Z(n34017));
    LUT4 i3104_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[434])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3096_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[435])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3096_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3088_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[436])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3088_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3080_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[437])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3080_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3072_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[438])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3072_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3064_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[439])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3064_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15171 (.BLUT(n33542), .ALUT(n33543), .C0(y_1_delay[1]), .Z(n33555));
    LUT4 i3056_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[440])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3056_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15261 (.BLUT(n33629), .ALUT(n33630), .C0(y_1_delay[1]), .Z(n33645));
    LUT4 i3048_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[441])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3048_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3040_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[442])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3040_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3032_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[443])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3032_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3024_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[444])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3024_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3016_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[445])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3016_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3008_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[446])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3008_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3000_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_i[4] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[447])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3000_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7209_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[432])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7209_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7201_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[433])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7201_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7193_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[434])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7193_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7185_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[435])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7177_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[436])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7177_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7169_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[437])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7169_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7161_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[438])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7161_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15758 (.BLUT(n34127), .ALUT(n34128), .C0(y_1_delay[1]), .Z(n34142));
    FD1P3AX result_i_31___i64 (.D(result_i_ns_0__15__N_517[63]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i64.GSR = "ENABLED";
    LUT4 i7153_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[439])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7153_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7145_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[440])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7145_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7137_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[441])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7137_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX din_i_reg_i1 (.D(din_i_c_0), .CK(clk_c), .Q(din_i_reg[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i1.GSR = "ENABLED";
    GSR GSR_INST (.GSR(rst_n_c));
    LUT4 i7129_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[442])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7129_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7121_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[443])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7113_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[444])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7113_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15172 (.BLUT(n33544), .ALUT(n33545), .C0(y_1_delay[1]), .Z(n33556));
    LUT4 i7105_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[445])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7105_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i63 (.D(result_i_ns_0__15__N_517[62]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i63.GSR = "ENABLED";
    PFUMX i15634 (.BLUT(n34003), .ALUT(n34004), .C0(y_1_delay[1]), .Z(n34018));
    PFUMX i15635 (.BLUT(n34005), .ALUT(n34006), .C0(y_1_delay[1]), .Z(n34019));
    PFUMX i15636 (.BLUT(n34007), .ALUT(n34008), .C0(y_1_delay[1]), .Z(n34020));
    PFUMX i15637 (.BLUT(n34009), .ALUT(n34010), .C0(y_1_delay[1]), .Z(n34021));
    PFUMX i15638 (.BLUT(n34011), .ALUT(n34012), .C0(y_1_delay[1]), .Z(n34022));
    PFUMX i15639 (.BLUT(n34013), .ALUT(n34014), .C0(y_1_delay[1]), .Z(n34023));
    PFUMX i15262 (.BLUT(n33631), .ALUT(n33632), .C0(y_1_delay[1]), .Z(n33646));
    PFUMX i15263 (.BLUT(n33633), .ALUT(n33634), .C0(y_1_delay[1]), .Z(n33647));
    PFUMX i15640 (.BLUT(n34015), .ALUT(n34016), .C0(y_1_delay[1]), .Z(n34024));
    PFUMX i15264 (.BLUT(n33635), .ALUT(n33636), .C0(y_1_delay[1]), .Z(n33648));
    PFUMX i15265 (.BLUT(n33637), .ALUT(n33638), .C0(y_1_delay[1]), .Z(n33649));
    PFUMX i15266 (.BLUT(n33639), .ALUT(n33640), .C0(y_1_delay[1]), .Z(n33650));
    PFUMX i15267 (.BLUT(n33641), .ALUT(n33642), .C0(y_1_delay[1]), .Z(n33651));
    PFUMX i15268 (.BLUT(n33643), .ALUT(n33644), .C0(y_1_delay[1]), .Z(n33652));
    LUT4 i7097_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[446])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7097_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15139 (.BLUT(n33509), .ALUT(n33510), .C0(y_1_delay[1]), .Z(n33523));
    LUT4 i7089_3_lut_4_lut (.A(n34716), .B(n34705), .C(\result_r[4] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[447])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7089_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3248_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[416])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3248_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3240_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[417])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3240_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3232_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[418])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3232_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3224_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[419])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3224_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15173 (.BLUT(n33546), .ALUT(n33547), .C0(y_1_delay[1]), .Z(n33557));
    LUT4 i3216_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[420])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3216_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3208_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[421])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3208_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3200_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[422])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3200_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15140 (.BLUT(n33511), .ALUT(n33512), .C0(y_1_delay[1]), .Z(n33524));
    LUT4 i3192_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[423])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3184_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[424])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3184_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15666 (.BLUT(n34036), .ALUT(n34037), .C0(y_1_delay[1]), .Z(n34050));
    PFUMX i15478 (.BLUT(n33846), .ALUT(n33847), .C0(y_1_delay[1]), .Z(n33862));
    LUT4 i3176_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[425])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3176_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3168_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[426])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3168_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3160_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[427])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3160_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3152_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[428])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3152_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3144_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[429])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3144_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15759 (.BLUT(n34129), .ALUT(n34130), .C0(y_1_delay[1]), .Z(n34143));
    LUT4 i3136_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[430])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3136_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15141 (.BLUT(n33513), .ALUT(n33514), .C0(y_1_delay[1]), .Z(n33525));
    LUT4 i3128_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_i[5] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[431])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7337_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[416])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7337_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i62 (.D(result_i_ns_0__15__N_517[61]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i62.GSR = "ENABLED";
    FD1P3AX result_i_31___i61 (.D(result_i_ns_0__15__N_517[60]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i61.GSR = "ENABLED";
    FD1P3AX result_i_31___i60 (.D(result_i_ns_0__15__N_517[59]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i60.GSR = "ENABLED";
    FD1P3AX result_i_31___i59 (.D(result_i_ns_0__15__N_517[58]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i59.GSR = "ENABLED";
    FD1P3AX result_i_31___i58 (.D(result_i_ns_0__15__N_517[57]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i58.GSR = "ENABLED";
    FD1P3AX result_i_31___i57 (.D(result_i_ns_0__15__N_517[56]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i57.GSR = "ENABLED";
    FD1P3AX result_i_31___i56 (.D(result_i_ns_0__15__N_517[55]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i56.GSR = "ENABLED";
    FD1P3AX result_i_31___i55 (.D(result_i_ns_0__15__N_517[54]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i55.GSR = "ENABLED";
    FD1P3AX result_i_31___i54 (.D(result_i_ns_0__15__N_517[53]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i54.GSR = "ENABLED";
    FD1P3AX result_i_31___i53 (.D(result_i_ns_0__15__N_517[52]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i53.GSR = "ENABLED";
    FD1P3AX result_i_31___i52 (.D(result_i_ns_0__15__N_517[51]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i52.GSR = "ENABLED";
    FD1P3AX result_i_31___i51 (.D(result_i_ns_0__15__N_517[50]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i51.GSR = "ENABLED";
    FD1P3AX result_i_31___i50 (.D(result_i_ns_0__15__N_517[49]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i50.GSR = "ENABLED";
    FD1P3AX result_i_31___i49 (.D(result_i_ns_0__15__N_517[48]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[28] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i49.GSR = "ENABLED";
    FD1P3AX result_i_31___i48 (.D(result_i_ns_0__15__N_517[47]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i48.GSR = "ENABLED";
    FD1P3AX result_i_31___i47 (.D(result_i_ns_0__15__N_517[46]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i47.GSR = "ENABLED";
    LUT4 i7329_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[417])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7329_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7321_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[418])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7321_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7313_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[419])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7313_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7305_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[420])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7305_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15479 (.BLUT(n33848), .ALUT(n33849), .C0(y_1_delay[1]), .Z(n33863));
    LUT4 i7297_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[421])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7297_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7289_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[422])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7289_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7281_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[423])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7281_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7273_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[424])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7273_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7265_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[425])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7265_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7257_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[426])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7257_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7249_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[427])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7249_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7241_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[428])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7241_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7233_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[429])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7233_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7225_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[430])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7225_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7217_3_lut_4_lut (.A(n34716), .B(n34706), .C(\result_r[5] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[431])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7217_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3376_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[400])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3376_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15480 (.BLUT(n33850), .ALUT(n33851), .C0(y_1_delay[1]), .Z(n33864));
    LUT4 i3368_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[401])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3368_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15142 (.BLUT(n33515), .ALUT(n33516), .C0(y_1_delay[1]), .Z(n33526));
    LUT4 i3360_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[402])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3360_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3352_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[403])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3352_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3344_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[404])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3344_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3336_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[405])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3336_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3328_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[406])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3328_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3320_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[407])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3320_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3312_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[408])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3312_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15481 (.BLUT(n33852), .ALUT(n33853), .C0(y_1_delay[1]), .Z(n33865));
    LUT4 i3304_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[409])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3304_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3296_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[410])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3296_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3288_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[411])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3288_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3280_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[412])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3280_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3272_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[413])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3272_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3264_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[414])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3264_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i46 (.D(result_i_ns_0__15__N_517[45]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i46.GSR = "ENABLED";
    FD1P3AX result_i_31___i45 (.D(result_i_ns_0__15__N_517[44]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i45.GSR = "ENABLED";
    FD1P3AX result_i_31___i44 (.D(result_i_ns_0__15__N_517[43]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i44.GSR = "ENABLED";
    LUT4 i3256_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_i[6] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[415])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3256_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i43 (.D(result_i_ns_0__15__N_517[42]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i43.GSR = "ENABLED";
    FD1P3AX result_i_31___i42 (.D(result_i_ns_0__15__N_517[41]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i42.GSR = "ENABLED";
    FD1P3AX result_i_31___i41 (.D(result_i_ns_0__15__N_517[40]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i41.GSR = "ENABLED";
    FD1P3AX result_i_31___i40 (.D(result_i_ns_0__15__N_517[39]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i40.GSR = "ENABLED";
    FD1P3AX result_i_31___i39 (.D(result_i_ns_0__15__N_517[38]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i39.GSR = "ENABLED";
    FD1P3AX result_i_31___i38 (.D(result_i_ns_0__15__N_517[37]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i38.GSR = "ENABLED";
    FD1P3AX result_i_31___i37 (.D(result_i_ns_0__15__N_517[36]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i37.GSR = "ENABLED";
    FD1P3AX result_i_31___i36 (.D(result_i_ns_0__15__N_517[35]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i36.GSR = "ENABLED";
    FD1P3AX result_i_31___i35 (.D(result_i_ns_0__15__N_517[34]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i35.GSR = "ENABLED";
    FD1P3AX result_i_31___i34 (.D(result_i_ns_0__15__N_517[33]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i34.GSR = "ENABLED";
    FD1P3AX count_y_689__i0 (.D(n35), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(count_y[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689__i0.GSR = "ENABLED";
    FD1P3AX result_i_31___i33 (.D(result_i_ns_0__15__N_517[32]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[29] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i33.GSR = "ENABLED";
    OB dout_r_pad_13 (.I(dout_r_c_13), .O(dout_r[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_14 (.I(dout_r_c_14), .O(dout_r[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    FD1P3AX result_i_31___i32 (.D(result_i_ns_0__15__N_517[31]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i32.GSR = "ENABLED";
    FD1P3AX result_i_31___i31 (.D(result_i_ns_0__15__N_517[30]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i31.GSR = "ENABLED";
    FD1P3AX result_i_31___i30 (.D(result_i_ns_0__15__N_517[29]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i30.GSR = "ENABLED";
    LUT4 i7465_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[400])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7465_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i29 (.D(result_i_ns_0__15__N_517[28]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i29.GSR = "ENABLED";
    FD1P3AX result_i_31___i28 (.D(result_i_ns_0__15__N_517[27]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i28.GSR = "ENABLED";
    FD1P3AX result_i_31___i27 (.D(result_i_ns_0__15__N_517[26]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i27.GSR = "ENABLED";
    FD1P3AX result_i_31___i26 (.D(result_i_ns_0__15__N_517[25]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i26.GSR = "ENABLED";
    FD1P3AX result_i_31___i25 (.D(result_i_ns_0__15__N_517[24]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i25.GSR = "ENABLED";
    CCU2C _add_1_1012_add_4_2 (.A0(op_r_23__N_1268_adj_7324[0]), .B0(op_i_23__N_1310_adj_7329[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[1]), 
          .B1(op_i_23__N_1310_adj_7329[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n31807));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1012_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_2.INJECT1_1 = "NO";
    FD1P3AX result_i_31___i24 (.D(result_i_ns_0__15__N_517[23]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i24.GSR = "ENABLED";
    FD1P3AX result_i_31___i23 (.D(result_i_ns_0__15__N_517[22]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i23.GSR = "ENABLED";
    FD1P3AX result_i_31___i22 (.D(result_i_ns_0__15__N_517[21]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i22.GSR = "ENABLED";
    FD1P3AX result_i_31___i21 (.D(result_i_ns_0__15__N_517[20]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i21.GSR = "ENABLED";
    FD1P3AX result_i_31___i20 (.D(result_i_ns_0__15__N_517[19]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i20.GSR = "ENABLED";
    FD1P3AX result_i_31___i19 (.D(result_i_ns_0__15__N_517[18]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i19.GSR = "ENABLED";
    FD1P3AX result_i_31___i18 (.D(result_i_ns_0__15__N_517[17]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i18.GSR = "ENABLED";
    FD1P3AX result_i_31___i17 (.D(result_i_ns_0__15__N_517[16]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[30] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i17.GSR = "ENABLED";
    FD1P3AX result_i_31___i16 (.D(result_i_ns_0__15__N_517[15]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i16.GSR = "ENABLED";
    FD1P3AX result_i_31___i15 (.D(result_i_ns_0__15__N_517[14]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i15.GSR = "ENABLED";
    CCU2C _add_1_1131_add_4_9 (.A0(n30197), .B0(n34736), .C0(count[5]), 
          .D0(n17), .A1(n28598), .B1(count[5]), .C1(n32928), .D1(n33013), 
          .CIN(n31804), .COUT(n31805), .S0(n12351), .S1(n12352));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1131_add_4_9.INIT0 = 16'h8878;
    defparam _add_1_1131_add_4_9.INIT1 = 16'h4bbb;
    defparam _add_1_1131_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1131_add_4_9.INJECT1_1 = "NO";
    FD1P3AX result_i_31___i14 (.D(result_i_ns_0__15__N_517[13]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i14.GSR = "ENABLED";
    FD1P3AX result_i_31___i13 (.D(result_i_ns_0__15__N_517[12]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i13.GSR = "ENABLED";
    FD1P3AX result_i_31___i12 (.D(result_i_ns_0__15__N_517[11]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i12.GSR = "ENABLED";
    FD1P3AX result_i_31___i11 (.D(result_i_ns_0__15__N_517[10]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i11.GSR = "ENABLED";
    FD1P3AX result_i_31___i10 (.D(result_i_ns_0__15__N_517[9]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i10.GSR = "ENABLED";
    LUT4 i7457_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[401])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7457_3_lut_4_lut.init = 16'hf1e0;
    OB dout_r_pad_4 (.I(dout_r_c_4), .O(dout_r[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    FD1P3AX result_i_31___i9 (.D(result_i_ns_0__15__N_517[8]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i9.GSR = "ENABLED";
    OB dout_r_pad_15 (.I(dout_r_c_15), .O(dout_r[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB out_valid_pad (.I(out_valid_c), .O(out_valid));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(18[8:17])
    LUT4 i7449_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[402])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7449_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7441_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[403])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7441_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15760 (.BLUT(n34131), .ALUT(n34132), .C0(y_1_delay[1]), .Z(n34144));
    LUT4 i7433_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[404])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7433_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i8 (.D(result_i_ns_0__15__N_517[7]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i8.GSR = "ENABLED";
    FD1P3AX result_i_31___i7 (.D(result_i_ns_0__15__N_517[6]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i7.GSR = "ENABLED";
    FD1P3AX result_i_31___i6 (.D(result_i_ns_0__15__N_517[5]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i6.GSR = "ENABLED";
    FD1P3AX result_i_31___i5 (.D(result_i_ns_0__15__N_517[4]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i5.GSR = "ENABLED";
    FD1P3AX result_i_31___i4 (.D(result_i_ns_0__15__N_517[3]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i4.GSR = "ENABLED";
    FD1P3AX result_i_31___i3 (.D(result_i_ns_0__15__N_517[2]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i3.GSR = "ENABLED";
    FD1P3AX result_i_31___i2 (.D(result_i_ns_0__15__N_517[1]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[31] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i2.GSR = "ENABLED";
    FD1S3AX din_i_reg_i12 (.D(din_i_c_11), .CK(clk_c), .Q(din_i_reg[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i12.GSR = "ENABLED";
    FD1S3AX din_i_reg_i11 (.D(din_i_c_10), .CK(clk_c), .Q(din_i_reg[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i11.GSR = "ENABLED";
    FD1S3AX din_i_reg_i10 (.D(din_i_c_9), .CK(clk_c), .Q(din_i_reg[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i10.GSR = "ENABLED";
    FD1S3AX din_i_reg_i9 (.D(din_i_c_8), .CK(clk_c), .Q(din_i_reg[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i9.GSR = "ENABLED";
    FD1S3AX din_i_reg_i8 (.D(din_i_c_7), .CK(clk_c), .Q(din_i_reg[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i8.GSR = "ENABLED";
    FD1S3AX din_i_reg_i7 (.D(din_i_c_6), .CK(clk_c), .Q(din_i_reg[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i7.GSR = "ENABLED";
    FD1S3AX din_i_reg_i6 (.D(din_i_c_5), .CK(clk_c), .Q(din_i_reg[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i6.GSR = "ENABLED";
    FD1S3AX din_i_reg_i5 (.D(din_i_c_4), .CK(clk_c), .Q(din_i_reg[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i5.GSR = "ENABLED";
    FD1S3AX din_i_reg_i4 (.D(din_i_c_3), .CK(clk_c), .Q(din_i_reg[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i4.GSR = "ENABLED";
    FD1S3AX din_i_reg_i3 (.D(din_i_c_2), .CK(clk_c), .Q(din_i_reg[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i3.GSR = "ENABLED";
    FD1S3AX din_i_reg_i2 (.D(din_i_c_1), .CK(clk_c), .Q(din_i_reg[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_i_reg_i2.GSR = "ENABLED";
    FD1P3AX result_i_31___i87 (.D(result_i_ns_0__15__N_517[86]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i87.GSR = "ENABLED";
    PFUMX i15174 (.BLUT(n33548), .ALUT(n33549), .C0(y_1_delay[1]), .Z(n33558));
    PFUMX i15143 (.BLUT(n33517), .ALUT(n33518), .C0(y_1_delay[1]), .Z(n33527));
    LUT4 i7425_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[405])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7425_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1070_add_4_20 (.A0(shift_1_dout_i[18]), .B0(shift_1_dout_r[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[19]), .B1(shift_1_dout_r[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32371), .COUT(n32372), .S0(n11574), 
          .S1(n11575));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_14 (.A0(op_r_23__N_1268[12]), .B0(op_i_23__N_1310[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[13]), .B1(op_i_23__N_1310[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32085), .COUT(n32086), .S0(op_i_23__N_1130[12]), 
          .S1(op_i_23__N_1130[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_12 (.A0(op_r_23__N_1268[10]), .B0(op_i_23__N_1310[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[11]), .B1(op_i_23__N_1310[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32084), .COUT(n32085), .S0(op_i_23__N_1130[10]), 
          .S1(op_i_23__N_1130[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_18 (.A0(shift_1_dout_i[16]), .B0(shift_1_dout_r[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[17]), .B1(shift_1_dout_r[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32370), .COUT(n32371), .S0(n11572), 
          .S1(n11573));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_10 (.A0(op_r_23__N_1268[8]), .B0(op_i_23__N_1310[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[9]), .B1(op_i_23__N_1310[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32083), .COUT(n32084), .S0(op_i_23__N_1130[8]), 
          .S1(op_i_23__N_1130[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_8 (.A0(op_r_23__N_1268[6]), .B0(op_i_23__N_1310[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[7]), .B1(op_i_23__N_1310[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32082), .COUT(n32083));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_8.INJECT1_1 = "NO";
    PFUMX i15482 (.BLUT(n33854), .ALUT(n33855), .C0(y_1_delay[1]), .Z(n33866));
    CCU2C _add_1_1070_add_4_16 (.A0(shift_1_dout_i[14]), .B0(shift_1_dout_r[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[15]), .B1(shift_1_dout_r[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32369), .COUT(n32370), .S0(n11570), 
          .S1(n11571));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_6 (.A0(op_r_23__N_1268[4]), .B0(op_i_23__N_1310[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[5]), .B1(op_i_23__N_1310[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32081), .COUT(n32082));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_4 (.A0(op_r_23__N_1268[2]), .B0(op_i_23__N_1310[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[3]), .B1(op_i_23__N_1310[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32080), .COUT(n32081));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_14 (.A0(shift_1_dout_i[12]), .B0(shift_1_dout_r[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[13]), .B1(shift_1_dout_r[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32368), .COUT(n32369), .S0(n11568), 
          .S1(n11569));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_2 (.A0(op_r_23__N_1268[0]), .B0(op_i_23__N_1310[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[1]), .B1(op_i_23__N_1310[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32080));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_993_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_993_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_26 (.A0(op_i_23__N_1154_adj_7371[23]), .B0(n34841), 
          .C0(shift_2_dout_i[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n32079), .S0(delay_i_23__N_1202_adj_7428[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_26.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1113_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_26.INJECT1_1 = "NO";
    LUT4 i7417_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[406])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7417_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7409_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[407])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7409_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1070_add_4_12 (.A0(shift_1_dout_i[10]), .B0(shift_1_dout_r[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[11]), .B1(shift_1_dout_r[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32367), .COUT(n32368), .S0(n11566), 
          .S1(n11567));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_24 (.A0(op_i_23__N_1154_adj_7371[21]), .B0(n34841), 
          .C0(shift_2_dout_i[21]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[22]), 
          .B1(n34841), .C1(shift_2_dout_i[22]), .D1(VCC_net), .CIN(n32078), 
          .COUT(n32079), .S0(delay_i_23__N_1202_adj_7428[21]), .S1(delay_i_23__N_1202_adj_7428[22]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_24.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_24.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_22 (.A0(op_i_23__N_1154_adj_7371[19]), .B0(n34841), 
          .C0(shift_2_dout_i[19]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[20]), 
          .B1(n34841), .C1(shift_2_dout_i[20]), .D1(VCC_net), .CIN(n32077), 
          .COUT(n32078), .S0(delay_i_23__N_1202_adj_7428[19]), .S1(delay_i_23__N_1202_adj_7428[20]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_22.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_22.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_10 (.A0(shift_1_dout_i[8]), .B0(shift_1_dout_r[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[9]), .B1(shift_1_dout_r[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32366), .COUT(n32367), .S0(n11564), 
          .S1(n11565));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_20 (.A0(op_i_23__N_1154_adj_7371[17]), .B0(n34841), 
          .C0(shift_2_dout_i[17]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[18]), 
          .B1(n34841), .C1(shift_2_dout_i[18]), .D1(VCC_net), .CIN(n32076), 
          .COUT(n32077), .S0(delay_i_23__N_1202_adj_7428[17]), .S1(delay_i_23__N_1202_adj_7428[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_20.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_20.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_18 (.A0(op_i_23__N_1154_adj_7371[15]), .B0(n34841), 
          .C0(shift_2_dout_i[15]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[16]), 
          .B1(n34841), .C1(shift_2_dout_i[16]), .D1(VCC_net), .CIN(n32075), 
          .COUT(n32076), .S0(delay_i_23__N_1202_adj_7428[15]), .S1(delay_i_23__N_1202_adj_7428[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_18.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_18.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_18.INJECT1_1 = "NO";
    LUT4 i7401_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[408])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7401_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1070_add_4_8 (.A0(shift_1_dout_i[6]), .B0(shift_1_dout_r[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[7]), .B1(shift_1_dout_r[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32365), .COUT(n32366), .S0(n11562), 
          .S1(n11563));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_16 (.A0(op_i_23__N_1154_adj_7371[13]), .B0(n34841), 
          .C0(shift_2_dout_i[13]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[14]), 
          .B1(n34841), .C1(shift_2_dout_i[14]), .D1(VCC_net), .CIN(n32074), 
          .COUT(n32075), .S0(delay_i_23__N_1202_adj_7428[13]), .S1(delay_i_23__N_1202_adj_7428[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_16.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_16.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_14 (.A0(op_i_23__N_1154_adj_7371[11]), .B0(n34841), 
          .C0(shift_2_dout_i[11]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[12]), 
          .B1(n34841), .C1(shift_2_dout_i[12]), .D1(VCC_net), .CIN(n32073), 
          .COUT(n32074), .S0(delay_i_23__N_1202_adj_7428[11]), .S1(delay_i_23__N_1202_adj_7428[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_14.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_14.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_6 (.A0(shift_1_dout_i[4]), .B0(shift_1_dout_r[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[5]), .B1(shift_1_dout_r[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32364), .COUT(n32365), .S0(n11560), 
          .S1(n11561));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_12 (.A0(op_i_23__N_1154_adj_7371[9]), .B0(n34841), 
          .C0(shift_2_dout_i[9]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[10]), 
          .B1(n34841), .C1(shift_2_dout_i[10]), .D1(VCC_net), .CIN(n32072), 
          .COUT(n32073), .S0(delay_i_23__N_1202_adj_7428[9]), .S1(delay_i_23__N_1202_adj_7428[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_12.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_12.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_12.INJECT1_1 = "NO";
    LUT4 i7393_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[409])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7393_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7385_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[410])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7385_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7377_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[411])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7377_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7369_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[412])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7369_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1070_add_4_4 (.A0(shift_1_dout_i[2]), .B0(shift_1_dout_r[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[3]), .B1(shift_1_dout_r[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32363), .COUT(n32364), .S0(n11558), 
          .S1(n11559));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_10 (.A0(op_i_23__N_1154_adj_7371[7]), .B0(n34841), 
          .C0(shift_2_dout_i[7]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[8]), 
          .B1(n34841), .C1(shift_2_dout_i[8]), .D1(VCC_net), .CIN(n32071), 
          .COUT(n32072), .S0(delay_i_23__N_1202_adj_7428[7]), .S1(delay_i_23__N_1202_adj_7428[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_10.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_10.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_8 (.A0(op_i_23__N_1154_adj_7371[5]), .B0(n34841), 
          .C0(shift_2_dout_i[5]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[6]), 
          .B1(n34841), .C1(shift_2_dout_i[6]), .D1(VCC_net), .CIN(n32070), 
          .COUT(n32071), .S0(delay_i_23__N_1202_adj_7428[5]), .S1(delay_i_23__N_1202_adj_7428[6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_8.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_8.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_2 (.A0(shift_1_dout_i[0]), .B0(shift_1_dout_r[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[1]), .B1(shift_1_dout_r[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32363), .S1(n11557));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1070_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_6 (.A0(op_i_23__N_1154_adj_7371[3]), .B0(n34841), 
          .C0(shift_2_dout_i[3]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[4]), 
          .B1(n34841), .C1(shift_2_dout_i[4]), .D1(VCC_net), .CIN(n32069), 
          .COUT(n32070), .S0(delay_i_23__N_1202_adj_7428[3]), .S1(delay_i_23__N_1202_adj_7428[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_6.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_6.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1113_add_4_4 (.A0(op_i_23__N_1154_adj_7371[1]), .B0(n34841), 
          .C0(shift_2_dout_i[1]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[2]), 
          .B1(n34841), .C1(shift_2_dout_i[2]), .D1(VCC_net), .CIN(n32068), 
          .COUT(n32069), .S0(delay_i_23__N_1202_adj_7428[1]), .S1(delay_i_23__N_1202_adj_7428[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_4.INIT0 = 16'h8787;
    defparam _add_1_1113_add_4_4.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_4.INJECT1_1 = "NO";
    LUT4 i7361_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[413])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7361_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1113_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(op_i_23__N_1154_adj_7371[0]), .B1(n34841), 
          .C1(shift_2_dout_i[0]), .D1(VCC_net), .COUT(n32068), .S1(delay_i_23__N_1202_adj_7428[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1113_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1113_add_4_2.INIT1 = 16'h8787;
    defparam _add_1_1113_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1113_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_26 (.A0(shift_16_dout_i[23]), .B0(shift_16_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n32067), .S0(n319));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_990_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_26 (.A0(n9081), .B0(n65_adj_6576), .C0(GND_net), 
          .D0(VCC_net), .A1(n9080), .B1(n65_adj_6576), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32360), .S0(op_i_23__N_1310_adj_7491[30]), 
          .S1(op_i_23__N_1310_adj_7491[31]));
    defparam _add_1_1086_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_24 (.A0(shift_16_dout_i[22]), .B0(shift_16_dout_r[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[23]), .B1(shift_16_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32066), .COUT(n32067), .S0(n10005), 
          .S1(n10006));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_22 (.A0(shift_16_dout_i[20]), .B0(shift_16_dout_r[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[21]), .B1(shift_16_dout_r[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32065), .COUT(n32066), .S0(n10003), 
          .S1(n10004));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_22.INJECT1_1 = "NO";
    LUT4 i7353_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[414])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7353_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7345_3_lut_4_lut (.A(n34716), .B(n34707), .C(\result_r[6] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[415])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7345_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1086_add_4_24 (.A0(n9083), .B0(n67_adj_6574), .C0(GND_net), 
          .D0(VCC_net), .A1(n9082), .B1(n66_adj_6575), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32359), .COUT(n32360), .S0(op_i_23__N_1310_adj_7491[28]), 
          .S1(op_i_23__N_1310_adj_7491[29]));
    defparam _add_1_1086_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_20 (.A0(shift_16_dout_i[18]), .B0(shift_16_dout_r[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[19]), .B1(shift_16_dout_r[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32064), .COUT(n32065), .S0(n10001), 
          .S1(n10002));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_18 (.A0(shift_16_dout_i[16]), .B0(shift_16_dout_r[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[17]), .B1(shift_16_dout_r[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32063), .COUT(n32064), .S0(n9999), 
          .S1(n10000));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_22 (.A0(n9085), .B0(n69_adj_6572), .C0(GND_net), 
          .D0(VCC_net), .A1(n9084), .B1(n68_adj_6573), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32358), .COUT(n32359), .S0(op_i_23__N_1310_adj_7491[26]), 
          .S1(op_i_23__N_1310_adj_7491[27]));
    defparam _add_1_1086_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_16 (.A0(shift_16_dout_i[14]), .B0(shift_16_dout_r[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[15]), .B1(shift_16_dout_r[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32062), .COUT(n32063), .S0(n9997), 
          .S1(n9998));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_14 (.A0(shift_16_dout_i[12]), .B0(shift_16_dout_r[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[13]), .B1(shift_16_dout_r[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32061), .COUT(n32062), .S0(n9995), 
          .S1(n9996));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_14.INJECT1_1 = "NO";
    LUT4 i3505_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[384])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3505_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1086_add_4_20 (.A0(n9087), .B0(n71_adj_6570), .C0(GND_net), 
          .D0(VCC_net), .A1(n9086), .B1(n70_adj_6571), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32357), .COUT(n32358), .S0(op_i_23__N_1310_adj_7491[24]), 
          .S1(op_i_23__N_1310_adj_7491[25]));
    defparam _add_1_1086_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_12 (.A0(shift_16_dout_i[10]), .B0(shift_16_dout_r[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[11]), .B1(shift_16_dout_r[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32060), .COUT(n32061), .S0(n9993), 
          .S1(n9994));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_10 (.A0(shift_16_dout_i[8]), .B0(shift_16_dout_r[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[9]), .B1(shift_16_dout_r[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32059), .COUT(n32060), .S0(n9991), 
          .S1(n9992));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_18 (.A0(n9089), .B0(n73_adj_6568), .C0(GND_net), 
          .D0(VCC_net), .A1(n9088), .B1(n72_adj_6569), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32356), .COUT(n32357), .S0(op_i_23__N_1310_adj_7491[22]), 
          .S1(op_i_23__N_1310_adj_7491[23]));
    defparam _add_1_1086_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_8 (.A0(op_i_23__N_1154[6]), .B0(op_r_23__N_1106[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[7]), .B1(op_r_23__N_1106[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32058), .COUT(n32059), .S0(n9989), 
          .S1(n9990));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_8.INJECT1_1 = "NO";
    LUT4 i3497_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[385])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3497_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3489_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[386])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3489_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3481_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[387])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3481_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3473_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[388])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3473_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15845_3_lut (.A(\result_r[22] [1]), .B(\result_r[23] [1]), .C(y_1_delay[0]), 
         .Z(n34229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15845_3_lut.init = 16'hcaca;
    OB dout_r_pad_3 (.I(dout_r_c_3), .O(dout_r[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_2 (.I(dout_r_c_2), .O(dout_r[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_1 (.I(dout_r_c_1), .O(dout_r[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_r_pad_0 (.I(dout_r_c_0), .O(dout_r[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(19[26:32])
    OB dout_i_pad_15 (.I(dout_i_c_15), .O(dout_i[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_14 (.I(dout_i_c_14), .O(dout_i[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_13 (.I(dout_i_c_13), .O(dout_i[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_12 (.I(dout_i_c_12), .O(dout_i[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_11 (.I(dout_i_c_11), .O(dout_i[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_10 (.I(dout_i_c_10), .O(dout_i[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_9 (.I(dout_i_c_9), .O(dout_i[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_8 (.I(dout_i_c_8), .O(dout_i[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_7 (.I(dout_i_c_7), .O(dout_i[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_6 (.I(dout_i_c_6), .O(dout_i[6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_5 (.I(dout_i_c_5), .O(dout_i[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_4 (.I(dout_i_c_4), .O(dout_i[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_3 (.I(dout_i_c_3), .O(dout_i[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_2 (.I(dout_i_c_2), .O(dout_i[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_1 (.I(dout_i_c_1), .O(dout_i[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    OB dout_i_pad_0 (.I(dout_i_c_0), .O(dout_i[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(20[26:32])
    IB clk_pad (.I(clk), .O(clk_c));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(14[7:12])
    IB in_valid_pad (.I(in_valid), .O(in_valid_c));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(15[7:15])
    IB din_r_pad_11 (.I(din_r[11]), .O(din_r_c_11));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_10 (.I(din_r[10]), .O(din_r_c_10));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_9 (.I(din_r[9]), .O(din_r_c_9));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_8 (.I(din_r[8]), .O(din_r_c_8));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_7 (.I(din_r[7]), .O(din_r_c_7));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_6 (.I(din_r[6]), .O(din_r_c_6));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_5 (.I(din_r[5]), .O(din_r_c_5));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_4 (.I(din_r[4]), .O(din_r_c_4));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_3 (.I(din_r[3]), .O(din_r_c_3));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_2 (.I(din_r[2]), .O(din_r_c_2));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_1 (.I(din_r[1]), .O(din_r_c_1));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_r_pad_0 (.I(din_r[0]), .O(din_r_c_0));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(16[21:26])
    IB din_i_pad_11 (.I(din_i[11]), .O(din_i_c_11));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_10 (.I(din_i[10]), .O(din_i_c_10));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_9 (.I(din_i[9]), .O(din_i_c_9));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_8 (.I(din_i[8]), .O(din_i_c_8));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_7 (.I(din_i[7]), .O(din_i_c_7));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_6 (.I(din_i[6]), .O(din_i_c_6));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_5 (.I(din_i[5]), .O(din_i_c_5));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_4 (.I(din_i[4]), .O(din_i_c_4));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_3 (.I(din_i[3]), .O(din_i_c_3));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_2 (.I(din_i[2]), .O(din_i_c_2));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_1 (.I(din_i[1]), .O(din_i_c_1));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    IB din_i_pad_0 (.I(din_i[0]), .O(din_i_c_0));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(17[21:26])
    LUT4 i3465_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[389])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3465_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14941_3_lut (.A(\result_i[12] [15]), .B(\result_i[13] [15]), .C(y_1_delay[0]), 
         .Z(n33325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14941_3_lut.init = 16'hcaca;
    LUT4 i3457_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[390])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3457_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX result_i_31___i88 (.D(result_i_ns_0__15__N_517[87]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i88.GSR = "ENABLED";
    FD1P3AX result_i_31___i89 (.D(result_i_ns_0__15__N_517[88]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i89.GSR = "ENABLED";
    FD1P3AX result_i_31___i90 (.D(result_i_ns_0__15__N_517[89]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i90.GSR = "ENABLED";
    FD1P3AX result_i_31___i91 (.D(result_i_ns_0__15__N_517[90]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i91.GSR = "ENABLED";
    FD1P3AX result_i_31___i92 (.D(result_i_ns_0__15__N_517[91]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i92.GSR = "ENABLED";
    FD1P3AX result_i_31___i93 (.D(result_i_ns_0__15__N_517[92]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i93.GSR = "ENABLED";
    FD1P3AX result_i_31___i94 (.D(result_i_ns_0__15__N_517[93]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i94.GSR = "ENABLED";
    FD1P3AX result_i_31___i95 (.D(result_i_ns_0__15__N_517[94]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i95.GSR = "ENABLED";
    FD1P3AX result_i_31___i96 (.D(result_i_ns_0__15__N_517[95]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[26] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i96.GSR = "ENABLED";
    FD1P3AX result_i_31___i97 (.D(result_i_ns_0__15__N_517[96]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i97.GSR = "ENABLED";
    FD1P3AX result_i_31___i98 (.D(result_i_ns_0__15__N_517[97]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i98.GSR = "ENABLED";
    FD1P3AX result_i_31___i99 (.D(result_i_ns_0__15__N_517[98]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i99.GSR = "ENABLED";
    FD1P3AX result_i_31___i100 (.D(result_i_ns_0__15__N_517[99]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i100.GSR = "ENABLED";
    FD1P3AX result_i_31___i101 (.D(result_i_ns_0__15__N_517[100]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i101.GSR = "ENABLED";
    FD1P3AX result_i_31___i102 (.D(result_i_ns_0__15__N_517[101]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i102.GSR = "ENABLED";
    FD1P3AX result_i_31___i103 (.D(result_i_ns_0__15__N_517[102]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i103.GSR = "ENABLED";
    FD1P3AX result_i_31___i104 (.D(result_i_ns_0__15__N_517[103]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i104.GSR = "ENABLED";
    FD1P3AX result_i_31___i105 (.D(result_i_ns_0__15__N_517[104]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i105.GSR = "ENABLED";
    FD1P3AX result_i_31___i106 (.D(result_i_ns_0__15__N_517[105]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i106.GSR = "ENABLED";
    FD1P3AX result_i_31___i107 (.D(result_i_ns_0__15__N_517[106]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i107.GSR = "ENABLED";
    FD1P3AX result_i_31___i108 (.D(result_i_ns_0__15__N_517[107]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i108.GSR = "ENABLED";
    FD1P3AX result_i_31___i109 (.D(result_i_ns_0__15__N_517[108]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i109.GSR = "ENABLED";
    FD1P3AX result_i_31___i110 (.D(result_i_ns_0__15__N_517[109]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i110.GSR = "ENABLED";
    FD1P3AX result_i_31___i111 (.D(result_i_ns_0__15__N_517[110]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i111.GSR = "ENABLED";
    FD1P3AX result_i_31___i112 (.D(result_i_ns_0__15__N_517[111]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[25] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i112.GSR = "ENABLED";
    FD1P3AX result_i_31___i113 (.D(result_i_ns_0__15__N_517[112]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i113.GSR = "ENABLED";
    FD1P3AX result_i_31___i114 (.D(result_i_ns_0__15__N_517[113]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i114.GSR = "ENABLED";
    FD1P3AX result_i_31___i115 (.D(result_i_ns_0__15__N_517[114]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i115.GSR = "ENABLED";
    FD1P3AX result_i_31___i116 (.D(result_i_ns_0__15__N_517[115]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i116.GSR = "ENABLED";
    FD1P3AX result_i_31___i117 (.D(result_i_ns_0__15__N_517[116]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i117.GSR = "ENABLED";
    FD1P3AX result_i_31___i118 (.D(result_i_ns_0__15__N_517[117]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i118.GSR = "ENABLED";
    FD1P3AX result_i_31___i119 (.D(result_i_ns_0__15__N_517[118]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i119.GSR = "ENABLED";
    FD1P3AX result_i_31___i120 (.D(result_i_ns_0__15__N_517[119]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i120.GSR = "ENABLED";
    FD1P3AX result_i_31___i121 (.D(result_i_ns_0__15__N_517[120]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i121.GSR = "ENABLED";
    FD1P3AX result_i_31___i122 (.D(result_i_ns_0__15__N_517[121]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i122.GSR = "ENABLED";
    FD1P3AX result_i_31___i123 (.D(result_i_ns_0__15__N_517[122]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i123.GSR = "ENABLED";
    FD1P3AX result_i_31___i124 (.D(result_i_ns_0__15__N_517[123]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i124.GSR = "ENABLED";
    FD1P3AX result_i_31___i125 (.D(result_i_ns_0__15__N_517[124]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i125.GSR = "ENABLED";
    FD1P3AX result_i_31___i126 (.D(result_i_ns_0__15__N_517[125]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i126.GSR = "ENABLED";
    FD1P3AX result_i_31___i127 (.D(result_i_ns_0__15__N_517[126]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i127.GSR = "ENABLED";
    FD1P3AX result_i_31___i128 (.D(result_i_ns_0__15__N_517[127]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[24] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i128.GSR = "ENABLED";
    FD1P3AX result_i_31___i129 (.D(result_i_ns_0__15__N_517[128]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i129.GSR = "ENABLED";
    FD1P3AX result_i_31___i130 (.D(result_i_ns_0__15__N_517[129]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i130.GSR = "ENABLED";
    FD1P3AX result_i_31___i131 (.D(result_i_ns_0__15__N_517[130]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i131.GSR = "ENABLED";
    FD1P3AX result_i_31___i132 (.D(result_i_ns_0__15__N_517[131]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i132.GSR = "ENABLED";
    FD1P3AX result_i_31___i133 (.D(result_i_ns_0__15__N_517[132]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i133.GSR = "ENABLED";
    FD1P3AX result_i_31___i134 (.D(result_i_ns_0__15__N_517[133]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i134.GSR = "ENABLED";
    FD1P3AX result_i_31___i135 (.D(result_i_ns_0__15__N_517[134]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i135.GSR = "ENABLED";
    FD1P3AX result_i_31___i136 (.D(result_i_ns_0__15__N_517[135]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i136.GSR = "ENABLED";
    FD1P3AX result_i_31___i137 (.D(result_i_ns_0__15__N_517[136]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i137.GSR = "ENABLED";
    FD1P3AX result_i_31___i138 (.D(result_i_ns_0__15__N_517[137]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i138.GSR = "ENABLED";
    FD1P3AX result_i_31___i139 (.D(result_i_ns_0__15__N_517[138]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i139.GSR = "ENABLED";
    FD1P3AX result_i_31___i140 (.D(result_i_ns_0__15__N_517[139]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i140.GSR = "ENABLED";
    FD1P3AX result_i_31___i141 (.D(result_i_ns_0__15__N_517[140]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i141.GSR = "ENABLED";
    FD1P3AX result_i_31___i142 (.D(result_i_ns_0__15__N_517[141]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i142.GSR = "ENABLED";
    FD1P3AX result_i_31___i143 (.D(result_i_ns_0__15__N_517[142]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i143.GSR = "ENABLED";
    FD1P3AX result_i_31___i144 (.D(result_i_ns_0__15__N_517[143]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[23] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i144.GSR = "ENABLED";
    FD1P3AX result_i_31___i145 (.D(result_i_ns_0__15__N_517[144]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i145.GSR = "ENABLED";
    FD1P3AX result_i_31___i146 (.D(result_i_ns_0__15__N_517[145]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i146.GSR = "ENABLED";
    FD1P3AX result_i_31___i147 (.D(result_i_ns_0__15__N_517[146]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i147.GSR = "ENABLED";
    FD1P3AX result_i_31___i148 (.D(result_i_ns_0__15__N_517[147]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i148.GSR = "ENABLED";
    FD1P3AX result_i_31___i149 (.D(result_i_ns_0__15__N_517[148]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i149.GSR = "ENABLED";
    FD1P3AX result_i_31___i150 (.D(result_i_ns_0__15__N_517[149]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i150.GSR = "ENABLED";
    FD1P3AX result_i_31___i151 (.D(result_i_ns_0__15__N_517[150]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i151.GSR = "ENABLED";
    FD1P3AX result_i_31___i152 (.D(result_i_ns_0__15__N_517[151]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i152.GSR = "ENABLED";
    FD1P3AX result_i_31___i153 (.D(result_i_ns_0__15__N_517[152]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i153.GSR = "ENABLED";
    FD1P3AX result_i_31___i154 (.D(result_i_ns_0__15__N_517[153]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i154.GSR = "ENABLED";
    FD1P3AX result_i_31___i155 (.D(result_i_ns_0__15__N_517[154]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i155.GSR = "ENABLED";
    FD1P3AX result_i_31___i156 (.D(result_i_ns_0__15__N_517[155]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i156.GSR = "ENABLED";
    FD1P3AX result_i_31___i157 (.D(result_i_ns_0__15__N_517[156]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i157.GSR = "ENABLED";
    FD1P3AX result_i_31___i158 (.D(result_i_ns_0__15__N_517[157]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i158.GSR = "ENABLED";
    FD1P3AX result_i_31___i159 (.D(result_i_ns_0__15__N_517[158]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i159.GSR = "ENABLED";
    FD1P3AX result_i_31___i160 (.D(result_i_ns_0__15__N_517[159]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[22] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i160.GSR = "ENABLED";
    FD1P3AX result_i_31___i161 (.D(result_i_ns_0__15__N_517[160]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i161.GSR = "ENABLED";
    FD1P3AX result_i_31___i162 (.D(result_i_ns_0__15__N_517[161]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i162.GSR = "ENABLED";
    FD1P3AX result_i_31___i163 (.D(result_i_ns_0__15__N_517[162]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i163.GSR = "ENABLED";
    FD1P3AX result_i_31___i164 (.D(result_i_ns_0__15__N_517[163]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i164.GSR = "ENABLED";
    FD1P3AX result_i_31___i165 (.D(result_i_ns_0__15__N_517[164]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i165.GSR = "ENABLED";
    FD1P3AX result_i_31___i166 (.D(result_i_ns_0__15__N_517[165]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i166.GSR = "ENABLED";
    FD1P3AX result_i_31___i167 (.D(result_i_ns_0__15__N_517[166]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i167.GSR = "ENABLED";
    FD1P3AX result_i_31___i168 (.D(result_i_ns_0__15__N_517[167]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i168.GSR = "ENABLED";
    FD1P3AX result_i_31___i169 (.D(result_i_ns_0__15__N_517[168]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i169.GSR = "ENABLED";
    FD1P3AX result_i_31___i170 (.D(result_i_ns_0__15__N_517[169]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i170.GSR = "ENABLED";
    FD1P3AX result_i_31___i171 (.D(result_i_ns_0__15__N_517[170]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i171.GSR = "ENABLED";
    FD1P3AX result_i_31___i172 (.D(result_i_ns_0__15__N_517[171]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i172.GSR = "ENABLED";
    FD1P3AX result_i_31___i173 (.D(result_i_ns_0__15__N_517[172]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i173.GSR = "ENABLED";
    FD1P3AX result_i_31___i174 (.D(result_i_ns_0__15__N_517[173]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i174.GSR = "ENABLED";
    FD1P3AX result_i_31___i175 (.D(result_i_ns_0__15__N_517[174]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i175.GSR = "ENABLED";
    FD1P3AX result_i_31___i176 (.D(result_i_ns_0__15__N_517[175]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[21] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i176.GSR = "ENABLED";
    FD1P3AX result_i_31___i177 (.D(result_i_ns_0__15__N_517[176]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i177.GSR = "ENABLED";
    FD1P3AX result_i_31___i178 (.D(result_i_ns_0__15__N_517[177]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i178.GSR = "ENABLED";
    FD1P3AX result_i_31___i179 (.D(result_i_ns_0__15__N_517[178]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i179.GSR = "ENABLED";
    FD1P3AX result_i_31___i180 (.D(result_i_ns_0__15__N_517[179]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i180.GSR = "ENABLED";
    FD1P3AX result_i_31___i181 (.D(result_i_ns_0__15__N_517[180]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i181.GSR = "ENABLED";
    FD1P3AX result_i_31___i182 (.D(result_i_ns_0__15__N_517[181]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i182.GSR = "ENABLED";
    FD1P3AX result_i_31___i183 (.D(result_i_ns_0__15__N_517[182]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i183.GSR = "ENABLED";
    FD1P3AX result_i_31___i184 (.D(result_i_ns_0__15__N_517[183]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i184.GSR = "ENABLED";
    FD1P3AX result_i_31___i185 (.D(result_i_ns_0__15__N_517[184]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i185.GSR = "ENABLED";
    FD1P3AX result_i_31___i186 (.D(result_i_ns_0__15__N_517[185]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i186.GSR = "ENABLED";
    FD1P3AX result_i_31___i187 (.D(result_i_ns_0__15__N_517[186]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i187.GSR = "ENABLED";
    FD1P3AX result_i_31___i188 (.D(result_i_ns_0__15__N_517[187]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i188.GSR = "ENABLED";
    FD1P3AX result_i_31___i189 (.D(result_i_ns_0__15__N_517[188]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i189.GSR = "ENABLED";
    FD1P3AX result_i_31___i190 (.D(result_i_ns_0__15__N_517[189]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i190.GSR = "ENABLED";
    FD1P3AX result_i_31___i191 (.D(result_i_ns_0__15__N_517[190]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i191.GSR = "ENABLED";
    FD1P3AX result_i_31___i192 (.D(result_i_ns_0__15__N_517[191]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[20] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i192.GSR = "ENABLED";
    FD1P3AX result_i_31___i193 (.D(result_i_ns_0__15__N_517[192]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i193.GSR = "ENABLED";
    FD1P3AX result_i_31___i194 (.D(result_i_ns_0__15__N_517[193]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i194.GSR = "ENABLED";
    FD1P3AX result_i_31___i195 (.D(result_i_ns_0__15__N_517[194]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i195.GSR = "ENABLED";
    FD1P3AX result_i_31___i196 (.D(result_i_ns_0__15__N_517[195]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i196.GSR = "ENABLED";
    FD1P3AX result_i_31___i197 (.D(result_i_ns_0__15__N_517[196]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i197.GSR = "ENABLED";
    FD1P3AX result_i_31___i198 (.D(result_i_ns_0__15__N_517[197]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i198.GSR = "ENABLED";
    FD1P3AX result_i_31___i199 (.D(result_i_ns_0__15__N_517[198]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i199.GSR = "ENABLED";
    FD1P3AX result_i_31___i200 (.D(result_i_ns_0__15__N_517[199]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i200.GSR = "ENABLED";
    FD1P3AX result_i_31___i201 (.D(result_i_ns_0__15__N_517[200]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i201.GSR = "ENABLED";
    FD1P3AX result_i_31___i202 (.D(result_i_ns_0__15__N_517[201]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i202.GSR = "ENABLED";
    FD1P3AX result_i_31___i203 (.D(result_i_ns_0__15__N_517[202]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i203.GSR = "ENABLED";
    FD1P3AX result_i_31___i204 (.D(result_i_ns_0__15__N_517[203]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i204.GSR = "ENABLED";
    FD1P3AX result_i_31___i205 (.D(result_i_ns_0__15__N_517[204]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i205.GSR = "ENABLED";
    FD1P3AX result_i_31___i206 (.D(result_i_ns_0__15__N_517[205]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i206.GSR = "ENABLED";
    FD1P3AX result_i_31___i207 (.D(result_i_ns_0__15__N_517[206]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i207.GSR = "ENABLED";
    FD1P3AX result_i_31___i208 (.D(result_i_ns_0__15__N_517[207]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[19] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i208.GSR = "ENABLED";
    FD1P3AX result_i_31___i209 (.D(result_i_ns_0__15__N_517[208]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i209.GSR = "ENABLED";
    FD1P3AX result_i_31___i210 (.D(result_i_ns_0__15__N_517[209]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i210.GSR = "ENABLED";
    FD1P3AX result_i_31___i211 (.D(result_i_ns_0__15__N_517[210]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i211.GSR = "ENABLED";
    FD1P3AX result_i_31___i212 (.D(result_i_ns_0__15__N_517[211]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i212.GSR = "ENABLED";
    FD1P3AX result_i_31___i213 (.D(result_i_ns_0__15__N_517[212]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i213.GSR = "ENABLED";
    FD1P3AX result_i_31___i214 (.D(result_i_ns_0__15__N_517[213]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i214.GSR = "ENABLED";
    FD1P3AX result_i_31___i215 (.D(result_i_ns_0__15__N_517[214]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i215.GSR = "ENABLED";
    FD1P3AX result_i_31___i216 (.D(result_i_ns_0__15__N_517[215]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i216.GSR = "ENABLED";
    FD1P3AX result_i_31___i217 (.D(result_i_ns_0__15__N_517[216]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i217.GSR = "ENABLED";
    FD1P3AX result_i_31___i218 (.D(result_i_ns_0__15__N_517[217]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i218.GSR = "ENABLED";
    FD1P3AX result_i_31___i219 (.D(result_i_ns_0__15__N_517[218]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i219.GSR = "ENABLED";
    FD1P3AX result_i_31___i220 (.D(result_i_ns_0__15__N_517[219]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i220.GSR = "ENABLED";
    FD1P3AX result_i_31___i221 (.D(result_i_ns_0__15__N_517[220]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i221.GSR = "ENABLED";
    FD1P3AX result_i_31___i222 (.D(result_i_ns_0__15__N_517[221]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i222.GSR = "ENABLED";
    FD1P3AX result_i_31___i223 (.D(result_i_ns_0__15__N_517[222]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i223.GSR = "ENABLED";
    FD1P3AX result_i_31___i224 (.D(result_i_ns_0__15__N_517[223]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[18] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i224.GSR = "ENABLED";
    FD1P3AX result_i_31___i225 (.D(result_i_ns_0__15__N_517[224]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i225.GSR = "ENABLED";
    FD1P3AX result_i_31___i226 (.D(result_i_ns_0__15__N_517[225]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i226.GSR = "ENABLED";
    FD1P3AX result_i_31___i227 (.D(result_i_ns_0__15__N_517[226]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i227.GSR = "ENABLED";
    FD1P3AX result_i_31___i228 (.D(result_i_ns_0__15__N_517[227]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i228.GSR = "ENABLED";
    FD1P3AX result_i_31___i229 (.D(result_i_ns_0__15__N_517[228]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i229.GSR = "ENABLED";
    FD1P3AX result_i_31___i230 (.D(result_i_ns_0__15__N_517[229]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i230.GSR = "ENABLED";
    FD1P3AX result_i_31___i231 (.D(result_i_ns_0__15__N_517[230]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i231.GSR = "ENABLED";
    FD1P3AX result_i_31___i232 (.D(result_i_ns_0__15__N_517[231]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i232.GSR = "ENABLED";
    FD1P3AX result_i_31___i233 (.D(result_i_ns_0__15__N_517[232]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i233.GSR = "ENABLED";
    FD1P3AX result_i_31___i234 (.D(result_i_ns_0__15__N_517[233]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i234.GSR = "ENABLED";
    FD1P3AX result_i_31___i235 (.D(result_i_ns_0__15__N_517[234]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i235.GSR = "ENABLED";
    FD1P3AX result_i_31___i236 (.D(result_i_ns_0__15__N_517[235]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i236.GSR = "ENABLED";
    FD1P3AX result_i_31___i237 (.D(result_i_ns_0__15__N_517[236]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i237.GSR = "ENABLED";
    FD1P3AX result_i_31___i238 (.D(result_i_ns_0__15__N_517[237]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i238.GSR = "ENABLED";
    FD1P3AX result_i_31___i239 (.D(result_i_ns_0__15__N_517[238]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i239.GSR = "ENABLED";
    FD1P3AX result_i_31___i240 (.D(result_i_ns_0__15__N_517[239]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[17] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i240.GSR = "ENABLED";
    FD1P3AX result_i_31___i241 (.D(result_i_ns_0__15__N_517[240]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i241.GSR = "ENABLED";
    FD1P3AX result_i_31___i242 (.D(result_i_ns_0__15__N_517[241]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i242.GSR = "ENABLED";
    FD1P3AX result_i_31___i243 (.D(result_i_ns_0__15__N_517[242]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i243.GSR = "ENABLED";
    FD1P3AX result_i_31___i244 (.D(result_i_ns_0__15__N_517[243]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i244.GSR = "ENABLED";
    FD1P3AX result_i_31___i245 (.D(result_i_ns_0__15__N_517[244]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i245.GSR = "ENABLED";
    FD1P3AX result_i_31___i246 (.D(result_i_ns_0__15__N_517[245]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i246.GSR = "ENABLED";
    FD1P3AX result_i_31___i247 (.D(result_i_ns_0__15__N_517[246]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i247.GSR = "ENABLED";
    FD1P3AX result_i_31___i248 (.D(result_i_ns_0__15__N_517[247]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i248.GSR = "ENABLED";
    FD1P3AX result_i_31___i249 (.D(result_i_ns_0__15__N_517[248]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i249.GSR = "ENABLED";
    FD1P3AX result_i_31___i250 (.D(result_i_ns_0__15__N_517[249]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i250.GSR = "ENABLED";
    FD1P3AX result_i_31___i251 (.D(result_i_ns_0__15__N_517[250]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i251.GSR = "ENABLED";
    FD1P3AX result_i_31___i252 (.D(result_i_ns_0__15__N_517[251]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i252.GSR = "ENABLED";
    FD1P3AX result_i_31___i253 (.D(result_i_ns_0__15__N_517[252]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i253.GSR = "ENABLED";
    FD1P3AX result_i_31___i254 (.D(result_i_ns_0__15__N_517[253]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i254.GSR = "ENABLED";
    FD1P3AX result_i_31___i255 (.D(result_i_ns_0__15__N_517[254]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i255.GSR = "ENABLED";
    FD1P3AX result_i_31___i256 (.D(result_i_ns_0__15__N_517[255]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[16] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i256.GSR = "ENABLED";
    FD1P3AX result_i_31___i257 (.D(result_i_ns_0__15__N_517[256]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i257.GSR = "ENABLED";
    FD1P3AX result_i_31___i258 (.D(result_i_ns_0__15__N_517[257]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i258.GSR = "ENABLED";
    FD1P3AX result_i_31___i259 (.D(result_i_ns_0__15__N_517[258]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i259.GSR = "ENABLED";
    FD1P3AX result_i_31___i260 (.D(result_i_ns_0__15__N_517[259]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i260.GSR = "ENABLED";
    FD1P3AX result_i_31___i261 (.D(result_i_ns_0__15__N_517[260]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i261.GSR = "ENABLED";
    FD1P3AX result_i_31___i262 (.D(result_i_ns_0__15__N_517[261]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i262.GSR = "ENABLED";
    FD1P3AX result_i_31___i263 (.D(result_i_ns_0__15__N_517[262]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i263.GSR = "ENABLED";
    FD1P3AX result_i_31___i264 (.D(result_i_ns_0__15__N_517[263]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i264.GSR = "ENABLED";
    FD1P3AX result_i_31___i265 (.D(result_i_ns_0__15__N_517[264]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i265.GSR = "ENABLED";
    FD1P3AX result_i_31___i266 (.D(result_i_ns_0__15__N_517[265]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i266.GSR = "ENABLED";
    FD1P3AX result_i_31___i267 (.D(result_i_ns_0__15__N_517[266]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i267.GSR = "ENABLED";
    FD1P3AX result_i_31___i268 (.D(result_i_ns_0__15__N_517[267]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i268.GSR = "ENABLED";
    FD1P3AX result_i_31___i269 (.D(result_i_ns_0__15__N_517[268]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i269.GSR = "ENABLED";
    FD1P3AX result_i_31___i270 (.D(result_i_ns_0__15__N_517[269]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i270.GSR = "ENABLED";
    FD1P3AX result_i_31___i271 (.D(result_i_ns_0__15__N_517[270]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i271.GSR = "ENABLED";
    FD1P3AX result_i_31___i272 (.D(result_i_ns_0__15__N_517[271]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[15] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i272.GSR = "ENABLED";
    FD1P3AX result_i_31___i273 (.D(result_i_ns_0__15__N_517[272]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i273.GSR = "ENABLED";
    FD1P3AX result_i_31___i274 (.D(result_i_ns_0__15__N_517[273]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i274.GSR = "ENABLED";
    FD1P3AX result_i_31___i275 (.D(result_i_ns_0__15__N_517[274]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i275.GSR = "ENABLED";
    FD1P3AX result_i_31___i276 (.D(result_i_ns_0__15__N_517[275]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i276.GSR = "ENABLED";
    FD1P3AX result_i_31___i277 (.D(result_i_ns_0__15__N_517[276]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i277.GSR = "ENABLED";
    FD1P3AX result_i_31___i278 (.D(result_i_ns_0__15__N_517[277]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i278.GSR = "ENABLED";
    FD1P3AX result_i_31___i279 (.D(result_i_ns_0__15__N_517[278]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i279.GSR = "ENABLED";
    FD1P3AX result_i_31___i280 (.D(result_i_ns_0__15__N_517[279]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i280.GSR = "ENABLED";
    FD1P3AX result_i_31___i281 (.D(result_i_ns_0__15__N_517[280]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i281.GSR = "ENABLED";
    FD1P3AX result_i_31___i282 (.D(result_i_ns_0__15__N_517[281]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i282.GSR = "ENABLED";
    FD1P3AX result_i_31___i283 (.D(result_i_ns_0__15__N_517[282]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i283.GSR = "ENABLED";
    FD1P3AX result_i_31___i284 (.D(result_i_ns_0__15__N_517[283]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i284.GSR = "ENABLED";
    FD1P3AX result_i_31___i285 (.D(result_i_ns_0__15__N_517[284]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i285.GSR = "ENABLED";
    FD1P3AX result_i_31___i286 (.D(result_i_ns_0__15__N_517[285]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i286.GSR = "ENABLED";
    FD1P3AX result_i_31___i287 (.D(result_i_ns_0__15__N_517[286]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i287.GSR = "ENABLED";
    FD1P3AX result_i_31___i288 (.D(result_i_ns_0__15__N_517[287]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[14] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i288.GSR = "ENABLED";
    FD1P3AX result_i_31___i289 (.D(result_i_ns_0__15__N_517[288]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i289.GSR = "ENABLED";
    FD1P3AX result_i_31___i290 (.D(result_i_ns_0__15__N_517[289]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i290.GSR = "ENABLED";
    FD1P3AX result_i_31___i291 (.D(result_i_ns_0__15__N_517[290]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i291.GSR = "ENABLED";
    FD1P3AX result_i_31___i292 (.D(result_i_ns_0__15__N_517[291]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i292.GSR = "ENABLED";
    FD1P3AX result_i_31___i293 (.D(result_i_ns_0__15__N_517[292]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i293.GSR = "ENABLED";
    FD1P3AX result_i_31___i294 (.D(result_i_ns_0__15__N_517[293]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i294.GSR = "ENABLED";
    FD1P3AX result_i_31___i295 (.D(result_i_ns_0__15__N_517[294]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i295.GSR = "ENABLED";
    FD1P3AX result_i_31___i296 (.D(result_i_ns_0__15__N_517[295]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i296.GSR = "ENABLED";
    FD1P3AX result_i_31___i297 (.D(result_i_ns_0__15__N_517[296]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i297.GSR = "ENABLED";
    FD1P3AX result_i_31___i298 (.D(result_i_ns_0__15__N_517[297]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i298.GSR = "ENABLED";
    FD1P3AX result_i_31___i299 (.D(result_i_ns_0__15__N_517[298]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i299.GSR = "ENABLED";
    FD1P3AX result_i_31___i300 (.D(result_i_ns_0__15__N_517[299]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i300.GSR = "ENABLED";
    FD1P3AX result_i_31___i301 (.D(result_i_ns_0__15__N_517[300]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i301.GSR = "ENABLED";
    FD1P3AX result_i_31___i302 (.D(result_i_ns_0__15__N_517[301]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i302.GSR = "ENABLED";
    FD1P3AX result_i_31___i303 (.D(result_i_ns_0__15__N_517[302]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i303.GSR = "ENABLED";
    FD1P3AX result_i_31___i304 (.D(result_i_ns_0__15__N_517[303]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[13] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i304.GSR = "ENABLED";
    FD1P3AX result_i_31___i305 (.D(result_i_ns_0__15__N_517[304]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i305.GSR = "ENABLED";
    FD1P3AX result_i_31___i306 (.D(result_i_ns_0__15__N_517[305]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i306.GSR = "ENABLED";
    FD1P3AX result_i_31___i307 (.D(result_i_ns_0__15__N_517[306]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i307.GSR = "ENABLED";
    FD1P3AX result_i_31___i308 (.D(result_i_ns_0__15__N_517[307]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i308.GSR = "ENABLED";
    FD1P3AX result_i_31___i309 (.D(result_i_ns_0__15__N_517[308]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i309.GSR = "ENABLED";
    FD1P3AX result_i_31___i310 (.D(result_i_ns_0__15__N_517[309]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i310.GSR = "ENABLED";
    FD1P3AX result_i_31___i311 (.D(result_i_ns_0__15__N_517[310]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i311.GSR = "ENABLED";
    FD1P3AX result_i_31___i312 (.D(result_i_ns_0__15__N_517[311]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i312.GSR = "ENABLED";
    FD1P3AX result_i_31___i313 (.D(result_i_ns_0__15__N_517[312]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i313.GSR = "ENABLED";
    FD1P3AX result_i_31___i314 (.D(result_i_ns_0__15__N_517[313]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i314.GSR = "ENABLED";
    FD1P3AX result_i_31___i315 (.D(result_i_ns_0__15__N_517[314]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i315.GSR = "ENABLED";
    FD1P3AX result_i_31___i316 (.D(result_i_ns_0__15__N_517[315]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i316.GSR = "ENABLED";
    FD1P3AX result_i_31___i317 (.D(result_i_ns_0__15__N_517[316]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i317.GSR = "ENABLED";
    FD1P3AX result_i_31___i318 (.D(result_i_ns_0__15__N_517[317]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i318.GSR = "ENABLED";
    FD1P3AX result_i_31___i319 (.D(result_i_ns_0__15__N_517[318]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i319.GSR = "ENABLED";
    FD1P3AX result_i_31___i320 (.D(result_i_ns_0__15__N_517[319]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[12] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i320.GSR = "ENABLED";
    FD1P3AX result_i_31___i321 (.D(result_i_ns_0__15__N_517[320]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i321.GSR = "ENABLED";
    FD1P3AX result_i_31___i322 (.D(result_i_ns_0__15__N_517[321]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i322.GSR = "ENABLED";
    FD1P3AX result_i_31___i323 (.D(result_i_ns_0__15__N_517[322]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i323.GSR = "ENABLED";
    FD1P3AX result_i_31___i324 (.D(result_i_ns_0__15__N_517[323]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i324.GSR = "ENABLED";
    FD1P3AX result_i_31___i325 (.D(result_i_ns_0__15__N_517[324]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i325.GSR = "ENABLED";
    FD1P3AX result_i_31___i326 (.D(result_i_ns_0__15__N_517[325]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i326.GSR = "ENABLED";
    FD1P3AX result_i_31___i327 (.D(result_i_ns_0__15__N_517[326]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i327.GSR = "ENABLED";
    FD1P3AX result_i_31___i328 (.D(result_i_ns_0__15__N_517[327]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i328.GSR = "ENABLED";
    FD1P3AX result_i_31___i329 (.D(result_i_ns_0__15__N_517[328]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i329.GSR = "ENABLED";
    FD1P3AX result_i_31___i330 (.D(result_i_ns_0__15__N_517[329]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i330.GSR = "ENABLED";
    FD1P3AX result_i_31___i331 (.D(result_i_ns_0__15__N_517[330]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i331.GSR = "ENABLED";
    FD1P3AX result_i_31___i332 (.D(result_i_ns_0__15__N_517[331]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i332.GSR = "ENABLED";
    FD1P3AX result_i_31___i333 (.D(result_i_ns_0__15__N_517[332]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i333.GSR = "ENABLED";
    FD1P3AX result_i_31___i334 (.D(result_i_ns_0__15__N_517[333]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i334.GSR = "ENABLED";
    FD1P3AX result_i_31___i335 (.D(result_i_ns_0__15__N_517[334]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i335.GSR = "ENABLED";
    FD1P3AX result_i_31___i336 (.D(result_i_ns_0__15__N_517[335]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[11] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i336.GSR = "ENABLED";
    FD1P3AX result_i_31___i337 (.D(result_i_ns_0__15__N_517[336]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i337.GSR = "ENABLED";
    FD1P3AX result_i_31___i338 (.D(result_i_ns_0__15__N_517[337]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i338.GSR = "ENABLED";
    FD1P3AX result_i_31___i339 (.D(result_i_ns_0__15__N_517[338]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i339.GSR = "ENABLED";
    FD1P3AX result_i_31___i340 (.D(result_i_ns_0__15__N_517[339]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i340.GSR = "ENABLED";
    FD1P3AX result_i_31___i341 (.D(result_i_ns_0__15__N_517[340]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i341.GSR = "ENABLED";
    FD1P3AX result_i_31___i342 (.D(result_i_ns_0__15__N_517[341]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i342.GSR = "ENABLED";
    FD1P3AX result_i_31___i343 (.D(result_i_ns_0__15__N_517[342]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i343.GSR = "ENABLED";
    FD1P3AX result_i_31___i344 (.D(result_i_ns_0__15__N_517[343]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i344.GSR = "ENABLED";
    FD1P3AX result_i_31___i345 (.D(result_i_ns_0__15__N_517[344]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i345.GSR = "ENABLED";
    FD1P3AX result_i_31___i346 (.D(result_i_ns_0__15__N_517[345]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i346.GSR = "ENABLED";
    FD1P3AX result_i_31___i347 (.D(result_i_ns_0__15__N_517[346]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i347.GSR = "ENABLED";
    FD1P3AX result_i_31___i348 (.D(result_i_ns_0__15__N_517[347]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i348.GSR = "ENABLED";
    FD1P3AX result_i_31___i349 (.D(result_i_ns_0__15__N_517[348]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i349.GSR = "ENABLED";
    FD1P3AX result_i_31___i350 (.D(result_i_ns_0__15__N_517[349]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i350.GSR = "ENABLED";
    FD1P3AX result_i_31___i351 (.D(result_i_ns_0__15__N_517[350]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i351.GSR = "ENABLED";
    FD1P3AX result_i_31___i352 (.D(result_i_ns_0__15__N_517[351]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[10] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i352.GSR = "ENABLED";
    FD1P3AX result_i_31___i353 (.D(result_i_ns_0__15__N_517[352]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i353.GSR = "ENABLED";
    FD1P3AX result_i_31___i354 (.D(result_i_ns_0__15__N_517[353]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i354.GSR = "ENABLED";
    FD1P3AX result_i_31___i355 (.D(result_i_ns_0__15__N_517[354]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i355.GSR = "ENABLED";
    FD1P3AX result_i_31___i356 (.D(result_i_ns_0__15__N_517[355]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i356.GSR = "ENABLED";
    FD1P3AX result_i_31___i357 (.D(result_i_ns_0__15__N_517[356]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i357.GSR = "ENABLED";
    FD1P3AX result_i_31___i358 (.D(result_i_ns_0__15__N_517[357]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i358.GSR = "ENABLED";
    FD1P3AX result_i_31___i359 (.D(result_i_ns_0__15__N_517[358]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i359.GSR = "ENABLED";
    FD1P3AX result_i_31___i360 (.D(result_i_ns_0__15__N_517[359]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i360.GSR = "ENABLED";
    FD1P3AX result_i_31___i361 (.D(result_i_ns_0__15__N_517[360]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i361.GSR = "ENABLED";
    FD1P3AX result_i_31___i362 (.D(result_i_ns_0__15__N_517[361]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i362.GSR = "ENABLED";
    FD1P3AX result_i_31___i363 (.D(result_i_ns_0__15__N_517[362]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i363.GSR = "ENABLED";
    FD1P3AX result_i_31___i364 (.D(result_i_ns_0__15__N_517[363]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i364.GSR = "ENABLED";
    FD1P3AX result_i_31___i365 (.D(result_i_ns_0__15__N_517[364]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i365.GSR = "ENABLED";
    FD1P3AX result_i_31___i366 (.D(result_i_ns_0__15__N_517[365]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i366.GSR = "ENABLED";
    FD1P3AX result_i_31___i367 (.D(result_i_ns_0__15__N_517[366]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i367.GSR = "ENABLED";
    FD1P3AX result_i_31___i368 (.D(result_i_ns_0__15__N_517[367]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[9] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i368.GSR = "ENABLED";
    FD1P3AX result_i_31___i369 (.D(result_i_ns_0__15__N_517[368]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i369.GSR = "ENABLED";
    FD1P3AX result_i_31___i370 (.D(result_i_ns_0__15__N_517[369]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i370.GSR = "ENABLED";
    FD1P3AX result_i_31___i371 (.D(result_i_ns_0__15__N_517[370]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i371.GSR = "ENABLED";
    FD1P3AX result_i_31___i372 (.D(result_i_ns_0__15__N_517[371]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i372.GSR = "ENABLED";
    FD1P3AX result_i_31___i373 (.D(result_i_ns_0__15__N_517[372]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i373.GSR = "ENABLED";
    FD1P3AX result_i_31___i374 (.D(result_i_ns_0__15__N_517[373]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i374.GSR = "ENABLED";
    FD1P3AX result_i_31___i375 (.D(result_i_ns_0__15__N_517[374]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i375.GSR = "ENABLED";
    FD1P3AX result_i_31___i376 (.D(result_i_ns_0__15__N_517[375]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i376.GSR = "ENABLED";
    FD1P3AX result_i_31___i377 (.D(result_i_ns_0__15__N_517[376]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i377.GSR = "ENABLED";
    FD1P3AX result_i_31___i378 (.D(result_i_ns_0__15__N_517[377]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i378.GSR = "ENABLED";
    FD1P3AX result_i_31___i379 (.D(result_i_ns_0__15__N_517[378]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i379.GSR = "ENABLED";
    FD1P3AX result_i_31___i380 (.D(result_i_ns_0__15__N_517[379]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i380.GSR = "ENABLED";
    FD1P3AX result_i_31___i381 (.D(result_i_ns_0__15__N_517[380]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i381.GSR = "ENABLED";
    FD1P3AX result_i_31___i382 (.D(result_i_ns_0__15__N_517[381]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i382.GSR = "ENABLED";
    FD1P3AX result_i_31___i383 (.D(result_i_ns_0__15__N_517[382]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i383.GSR = "ENABLED";
    FD1P3AX result_i_31___i384 (.D(result_i_ns_0__15__N_517[383]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[8] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i384.GSR = "ENABLED";
    FD1P3AX result_i_31___i385 (.D(result_i_ns_0__15__N_517[384]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i385.GSR = "ENABLED";
    FD1P3AX result_i_31___i386 (.D(result_i_ns_0__15__N_517[385]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i386.GSR = "ENABLED";
    FD1P3AX result_i_31___i387 (.D(result_i_ns_0__15__N_517[386]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i387.GSR = "ENABLED";
    FD1P3AX result_i_31___i388 (.D(result_i_ns_0__15__N_517[387]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i388.GSR = "ENABLED";
    FD1P3AX result_i_31___i389 (.D(result_i_ns_0__15__N_517[388]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i389.GSR = "ENABLED";
    FD1P3AX result_i_31___i390 (.D(result_i_ns_0__15__N_517[389]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i390.GSR = "ENABLED";
    FD1P3AX result_i_31___i391 (.D(result_i_ns_0__15__N_517[390]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i391.GSR = "ENABLED";
    FD1P3AX result_i_31___i392 (.D(result_i_ns_0__15__N_517[391]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i392.GSR = "ENABLED";
    FD1P3AX result_i_31___i393 (.D(result_i_ns_0__15__N_517[392]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i393.GSR = "ENABLED";
    FD1P3AX result_i_31___i394 (.D(result_i_ns_0__15__N_517[393]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i394.GSR = "ENABLED";
    FD1P3AX result_i_31___i395 (.D(result_i_ns_0__15__N_517[394]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i395.GSR = "ENABLED";
    FD1P3AX result_i_31___i396 (.D(result_i_ns_0__15__N_517[395]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i396.GSR = "ENABLED";
    FD1P3AX result_i_31___i397 (.D(result_i_ns_0__15__N_517[396]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i397.GSR = "ENABLED";
    FD1P3AX result_i_31___i398 (.D(result_i_ns_0__15__N_517[397]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i398.GSR = "ENABLED";
    FD1P3AX result_i_31___i399 (.D(result_i_ns_0__15__N_517[398]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i399.GSR = "ENABLED";
    FD1P3AX result_i_31___i400 (.D(result_i_ns_0__15__N_517[399]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[7] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i400.GSR = "ENABLED";
    FD1P3AX result_i_31___i401 (.D(result_i_ns_0__15__N_517[400]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i401.GSR = "ENABLED";
    FD1P3AX result_i_31___i402 (.D(result_i_ns_0__15__N_517[401]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i402.GSR = "ENABLED";
    FD1P3AX result_i_31___i403 (.D(result_i_ns_0__15__N_517[402]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i403.GSR = "ENABLED";
    FD1P3AX result_i_31___i404 (.D(result_i_ns_0__15__N_517[403]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i404.GSR = "ENABLED";
    FD1P3AX result_i_31___i405 (.D(result_i_ns_0__15__N_517[404]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i405.GSR = "ENABLED";
    FD1P3AX result_i_31___i406 (.D(result_i_ns_0__15__N_517[405]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i406.GSR = "ENABLED";
    FD1P3AX result_i_31___i407 (.D(result_i_ns_0__15__N_517[406]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i407.GSR = "ENABLED";
    FD1P3AX result_i_31___i408 (.D(result_i_ns_0__15__N_517[407]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i408.GSR = "ENABLED";
    FD1P3AX result_i_31___i409 (.D(result_i_ns_0__15__N_517[408]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i409.GSR = "ENABLED";
    FD1P3AX result_i_31___i410 (.D(result_i_ns_0__15__N_517[409]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i410.GSR = "ENABLED";
    FD1P3AX result_i_31___i411 (.D(result_i_ns_0__15__N_517[410]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i411.GSR = "ENABLED";
    FD1P3AX result_i_31___i412 (.D(result_i_ns_0__15__N_517[411]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i412.GSR = "ENABLED";
    FD1P3AX result_i_31___i413 (.D(result_i_ns_0__15__N_517[412]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i413.GSR = "ENABLED";
    FD1P3AX result_i_31___i414 (.D(result_i_ns_0__15__N_517[413]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i414.GSR = "ENABLED";
    FD1P3AX result_i_31___i415 (.D(result_i_ns_0__15__N_517[414]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i415.GSR = "ENABLED";
    FD1P3AX result_i_31___i416 (.D(result_i_ns_0__15__N_517[415]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[6] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i416.GSR = "ENABLED";
    FD1P3AX result_i_31___i417 (.D(result_i_ns_0__15__N_517[416]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i417.GSR = "ENABLED";
    FD1P3AX result_i_31___i418 (.D(result_i_ns_0__15__N_517[417]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i418.GSR = "ENABLED";
    FD1P3AX result_i_31___i419 (.D(result_i_ns_0__15__N_517[418]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i419.GSR = "ENABLED";
    FD1P3AX result_i_31___i420 (.D(result_i_ns_0__15__N_517[419]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i420.GSR = "ENABLED";
    FD1P3AX result_i_31___i421 (.D(result_i_ns_0__15__N_517[420]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i421.GSR = "ENABLED";
    FD1P3AX result_i_31___i422 (.D(result_i_ns_0__15__N_517[421]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i422.GSR = "ENABLED";
    FD1P3AX result_i_31___i423 (.D(result_i_ns_0__15__N_517[422]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i423.GSR = "ENABLED";
    FD1P3AX result_i_31___i424 (.D(result_i_ns_0__15__N_517[423]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i424.GSR = "ENABLED";
    FD1P3AX result_i_31___i425 (.D(result_i_ns_0__15__N_517[424]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i425.GSR = "ENABLED";
    FD1P3AX result_i_31___i426 (.D(result_i_ns_0__15__N_517[425]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i426.GSR = "ENABLED";
    FD1P3AX result_i_31___i427 (.D(result_i_ns_0__15__N_517[426]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i427.GSR = "ENABLED";
    FD1P3AX result_i_31___i428 (.D(result_i_ns_0__15__N_517[427]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i428.GSR = "ENABLED";
    FD1P3AX result_i_31___i429 (.D(result_i_ns_0__15__N_517[428]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i429.GSR = "ENABLED";
    FD1P3AX result_i_31___i430 (.D(result_i_ns_0__15__N_517[429]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i430.GSR = "ENABLED";
    FD1P3AX result_i_31___i431 (.D(result_i_ns_0__15__N_517[430]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i431.GSR = "ENABLED";
    FD1P3AX result_i_31___i432 (.D(result_i_ns_0__15__N_517[431]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[5] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i432.GSR = "ENABLED";
    FD1P3AX result_i_31___i433 (.D(result_i_ns_0__15__N_517[432]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i433.GSR = "ENABLED";
    FD1P3AX result_i_31___i434 (.D(result_i_ns_0__15__N_517[433]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i434.GSR = "ENABLED";
    FD1P3AX result_i_31___i435 (.D(result_i_ns_0__15__N_517[434]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i435.GSR = "ENABLED";
    FD1P3AX result_i_31___i436 (.D(result_i_ns_0__15__N_517[435]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i436.GSR = "ENABLED";
    FD1P3AX result_i_31___i437 (.D(result_i_ns_0__15__N_517[436]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i437.GSR = "ENABLED";
    FD1P3AX result_i_31___i438 (.D(result_i_ns_0__15__N_517[437]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i438.GSR = "ENABLED";
    FD1P3AX result_i_31___i439 (.D(result_i_ns_0__15__N_517[438]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i439.GSR = "ENABLED";
    FD1P3AX result_i_31___i440 (.D(result_i_ns_0__15__N_517[439]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i440.GSR = "ENABLED";
    FD1P3AX result_i_31___i441 (.D(result_i_ns_0__15__N_517[440]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i441.GSR = "ENABLED";
    FD1P3AX result_i_31___i442 (.D(result_i_ns_0__15__N_517[441]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i442.GSR = "ENABLED";
    FD1P3AX result_i_31___i443 (.D(result_i_ns_0__15__N_517[442]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i443.GSR = "ENABLED";
    FD1P3AX result_i_31___i444 (.D(result_i_ns_0__15__N_517[443]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i444.GSR = "ENABLED";
    FD1P3AX result_i_31___i445 (.D(result_i_ns_0__15__N_517[444]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i445.GSR = "ENABLED";
    FD1P3AX result_i_31___i446 (.D(result_i_ns_0__15__N_517[445]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i446.GSR = "ENABLED";
    FD1P3AX result_i_31___i447 (.D(result_i_ns_0__15__N_517[446]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i447.GSR = "ENABLED";
    FD1P3AX result_i_31___i448 (.D(result_i_ns_0__15__N_517[447]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[4] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i448.GSR = "ENABLED";
    FD1P3AX result_i_31___i449 (.D(result_i_ns_0__15__N_517[448]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i449.GSR = "ENABLED";
    FD1P3AX result_i_31___i450 (.D(result_i_ns_0__15__N_517[449]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i450.GSR = "ENABLED";
    FD1P3AX result_i_31___i451 (.D(result_i_ns_0__15__N_517[450]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i451.GSR = "ENABLED";
    FD1P3AX result_i_31___i452 (.D(result_i_ns_0__15__N_517[451]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i452.GSR = "ENABLED";
    FD1P3AX result_i_31___i453 (.D(result_i_ns_0__15__N_517[452]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i453.GSR = "ENABLED";
    FD1P3AX result_i_31___i454 (.D(result_i_ns_0__15__N_517[453]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i454.GSR = "ENABLED";
    FD1P3AX result_i_31___i455 (.D(result_i_ns_0__15__N_517[454]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i455.GSR = "ENABLED";
    FD1P3AX result_i_31___i456 (.D(result_i_ns_0__15__N_517[455]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i456.GSR = "ENABLED";
    FD1P3AX result_i_31___i457 (.D(result_i_ns_0__15__N_517[456]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i457.GSR = "ENABLED";
    FD1P3AX result_i_31___i458 (.D(result_i_ns_0__15__N_517[457]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i458.GSR = "ENABLED";
    FD1P3AX result_i_31___i459 (.D(result_i_ns_0__15__N_517[458]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i459.GSR = "ENABLED";
    FD1P3AX result_i_31___i460 (.D(result_i_ns_0__15__N_517[459]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i460.GSR = "ENABLED";
    FD1P3AX result_i_31___i461 (.D(result_i_ns_0__15__N_517[460]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i461.GSR = "ENABLED";
    FD1P3AX result_i_31___i462 (.D(result_i_ns_0__15__N_517[461]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i462.GSR = "ENABLED";
    FD1P3AX result_i_31___i463 (.D(result_i_ns_0__15__N_517[462]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i463.GSR = "ENABLED";
    FD1P3AX result_i_31___i464 (.D(result_i_ns_0__15__N_517[463]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[3] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i464.GSR = "ENABLED";
    FD1P3AX result_i_31___i465 (.D(result_i_ns_0__15__N_517[464]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i465.GSR = "ENABLED";
    FD1P3AX result_i_31___i466 (.D(result_i_ns_0__15__N_517[465]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i466.GSR = "ENABLED";
    FD1P3AX result_i_31___i467 (.D(result_i_ns_0__15__N_517[466]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i467.GSR = "ENABLED";
    FD1P3AX result_i_31___i468 (.D(result_i_ns_0__15__N_517[467]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i468.GSR = "ENABLED";
    FD1P3AX result_i_31___i469 (.D(result_i_ns_0__15__N_517[468]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i469.GSR = "ENABLED";
    FD1P3AX result_i_31___i470 (.D(result_i_ns_0__15__N_517[469]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i470.GSR = "ENABLED";
    FD1P3AX result_i_31___i471 (.D(result_i_ns_0__15__N_517[470]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i471.GSR = "ENABLED";
    FD1P3AX result_i_31___i472 (.D(result_i_ns_0__15__N_517[471]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i472.GSR = "ENABLED";
    FD1P3AX result_i_31___i473 (.D(result_i_ns_0__15__N_517[472]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i473.GSR = "ENABLED";
    FD1P3AX result_i_31___i474 (.D(result_i_ns_0__15__N_517[473]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i474.GSR = "ENABLED";
    FD1P3AX result_i_31___i475 (.D(result_i_ns_0__15__N_517[474]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i475.GSR = "ENABLED";
    FD1P3AX result_i_31___i476 (.D(result_i_ns_0__15__N_517[475]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i476.GSR = "ENABLED";
    FD1P3AX result_i_31___i477 (.D(result_i_ns_0__15__N_517[476]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i477.GSR = "ENABLED";
    FD1P3AX result_i_31___i478 (.D(result_i_ns_0__15__N_517[477]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i478.GSR = "ENABLED";
    FD1P3AX result_i_31___i479 (.D(result_i_ns_0__15__N_517[478]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i479.GSR = "ENABLED";
    FD1P3AX result_i_31___i480 (.D(result_i_ns_0__15__N_517[479]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[2] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i480.GSR = "ENABLED";
    FD1P3AX result_i_31___i481 (.D(result_i_ns_0__15__N_517[480]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i481.GSR = "ENABLED";
    FD1P3AX result_i_31___i482 (.D(result_i_ns_0__15__N_517[481]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i482.GSR = "ENABLED";
    FD1P3AX result_i_31___i483 (.D(result_i_ns_0__15__N_517[482]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i483.GSR = "ENABLED";
    FD1P3AX result_i_31___i484 (.D(result_i_ns_0__15__N_517[483]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i484.GSR = "ENABLED";
    FD1P3AX result_i_31___i485 (.D(result_i_ns_0__15__N_517[484]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i485.GSR = "ENABLED";
    FD1P3AX result_i_31___i486 (.D(result_i_ns_0__15__N_517[485]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i486.GSR = "ENABLED";
    FD1P3AX result_i_31___i487 (.D(result_i_ns_0__15__N_517[486]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i487.GSR = "ENABLED";
    FD1P3AX result_i_31___i488 (.D(result_i_ns_0__15__N_517[487]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i488.GSR = "ENABLED";
    FD1P3AX result_i_31___i489 (.D(result_i_ns_0__15__N_517[488]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i489.GSR = "ENABLED";
    FD1P3AX result_i_31___i490 (.D(result_i_ns_0__15__N_517[489]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i490.GSR = "ENABLED";
    FD1P3AX result_i_31___i491 (.D(result_i_ns_0__15__N_517[490]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i491.GSR = "ENABLED";
    FD1P3AX result_i_31___i492 (.D(result_i_ns_0__15__N_517[491]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i492.GSR = "ENABLED";
    FD1P3AX result_i_31___i493 (.D(result_i_ns_0__15__N_517[492]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i493.GSR = "ENABLED";
    FD1P3AX result_i_31___i494 (.D(result_i_ns_0__15__N_517[493]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i494.GSR = "ENABLED";
    FD1P3AX result_i_31___i495 (.D(result_i_ns_0__15__N_517[494]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i495.GSR = "ENABLED";
    FD1P3AX result_i_31___i496 (.D(result_i_ns_0__15__N_517[495]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[1] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i496.GSR = "ENABLED";
    FD1P3AX result_i_31___i497 (.D(result_i_ns_0__15__N_517[496]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i497.GSR = "ENABLED";
    FD1P3AX result_i_31___i498 (.D(result_i_ns_0__15__N_517[497]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i498.GSR = "ENABLED";
    FD1P3AX result_i_31___i499 (.D(result_i_ns_0__15__N_517[498]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i499.GSR = "ENABLED";
    FD1P3AX result_i_31___i500 (.D(result_i_ns_0__15__N_517[499]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i500.GSR = "ENABLED";
    FD1P3AX result_i_31___i501 (.D(result_i_ns_0__15__N_517[500]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i501.GSR = "ENABLED";
    FD1P3AX result_i_31___i502 (.D(result_i_ns_0__15__N_517[501]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i502.GSR = "ENABLED";
    FD1P3AX result_i_31___i503 (.D(result_i_ns_0__15__N_517[502]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i503.GSR = "ENABLED";
    FD1P3AX result_i_31___i504 (.D(result_i_ns_0__15__N_517[503]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i504.GSR = "ENABLED";
    FD1P3AX result_i_31___i505 (.D(result_i_ns_0__15__N_517[504]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i505.GSR = "ENABLED";
    FD1P3AX result_i_31___i506 (.D(result_i_ns_0__15__N_517[505]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i506.GSR = "ENABLED";
    FD1P3AX result_i_31___i507 (.D(result_i_ns_0__15__N_517[506]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i507.GSR = "ENABLED";
    FD1P3AX result_i_31___i508 (.D(result_i_ns_0__15__N_517[507]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i508.GSR = "ENABLED";
    FD1P3AX result_i_31___i509 (.D(result_i_ns_0__15__N_517[508]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i509.GSR = "ENABLED";
    FD1P3AX result_i_31___i510 (.D(result_i_ns_0__15__N_517[509]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i510.GSR = "ENABLED";
    FD1P3AX result_i_31___i511 (.D(result_i_ns_0__15__N_517[510]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i511.GSR = "ENABLED";
    FD1P3AX result_i_31___i512 (.D(result_i_ns_0__15__N_517[511]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_i[0] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_i_31___i512.GSR = "ENABLED";
    FD1S3AX y_1_delay_i1 (.D(n34812), .CK(clk_c), .Q(y_1_delay[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam y_1_delay_i1.GSR = "ENABLED";
    FD1S3AX y_1_delay_i2 (.D(n34739), .CK(clk_c), .Q(y_1_delay[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam y_1_delay_i2.GSR = "ENABLED";
    FD1S3AX y_1_delay_i3 (.D(n34741), .CK(clk_c), .Q(y_1_delay[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam y_1_delay_i3.GSR = "ENABLED";
    FD1S3AX y_1_delay_i4 (.D(n34811), .CK(clk_c), .Q(y_1_delay[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam y_1_delay_i4.GSR = "ENABLED";
    LUT4 i15844_3_lut (.A(\result_r[20] [1]), .B(\result_r[21] [1]), .C(y_1_delay[0]), 
         .Z(n34228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15844_3_lut.init = 16'hcaca;
    LUT4 i3449_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[391])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3449_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3441_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[392])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3441_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3433_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[393])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3433_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3425_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[394])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3425_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3417_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[395])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3417_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3409_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[396])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3409_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3401_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[397])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3401_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3393_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[398])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3393_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3385_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_i[7] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[399])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3385_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX din_r_reg_i2 (.D(din_r_c_1), .CK(clk_c), .Q(din_r_reg[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i2.GSR = "ENABLED";
    LUT4 i15415_3_lut (.A(\result_r[30] [15]), .B(\result_r[31] [15]), .C(y_1_delay[0]), 
         .Z(n33799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15415_3_lut.init = 16'hcaca;
    FD1S3AX din_r_reg_i3 (.D(din_r_c_2), .CK(clk_c), .Q(din_r_reg[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i3.GSR = "ENABLED";
    FD1S3AX din_r_reg_i4 (.D(din_r_c_3), .CK(clk_c), .Q(din_r_reg[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i4.GSR = "ENABLED";
    FD1S3AX din_r_reg_i5 (.D(din_r_c_4), .CK(clk_c), .Q(din_r_reg[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i5.GSR = "ENABLED";
    FD1S3AX din_r_reg_i6 (.D(din_r_c_5), .CK(clk_c), .Q(din_r_reg[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i6.GSR = "ENABLED";
    FD1S3AX din_r_reg_i7 (.D(din_r_c_6), .CK(clk_c), .Q(din_r_reg[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i7.GSR = "ENABLED";
    FD1S3AX din_r_reg_i8 (.D(din_r_c_7), .CK(clk_c), .Q(din_r_reg[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i8.GSR = "ENABLED";
    FD1S3AX din_r_reg_i9 (.D(din_r_c_8), .CK(clk_c), .Q(din_r_reg[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i9.GSR = "ENABLED";
    FD1S3AX din_r_reg_i10 (.D(din_r_c_9), .CK(clk_c), .Q(din_r_reg[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i10.GSR = "ENABLED";
    FD1S3AX din_r_reg_i11 (.D(din_r_c_10), .CK(clk_c), .Q(din_r_reg[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i11.GSR = "ENABLED";
    FD1S3AX din_r_reg_i12 (.D(din_r_c_11), .CK(clk_c), .Q(din_r_reg[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam din_r_reg_i12.GSR = "ENABLED";
    LUT4 i7593_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[384])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7593_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2631_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[493])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2631_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i7585_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[385])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7585_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15843_3_lut (.A(\result_r[18] [1]), .B(\result_r[19] [1]), .C(y_1_delay[0]), 
         .Z(n34227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15843_3_lut.init = 16'hcaca;
    LUT4 i7577_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[386])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7577_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7569_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[387])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7569_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7561_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[388])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7561_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7553_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[389])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7553_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7545_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[390])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7545_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1031_add_4_21 (.A0(n31484), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[18]), .A1(n31482), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[19]), .CIN(n31962), .COUT(n31963), .S0(op_i_23__N_1154_adj_7371[18]), 
          .S1(op_i_23__N_1154_adj_7371[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_21.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_21.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_19 (.A0(n31488), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[16]), .A1(n31486), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[17]), .CIN(n31961), .COUT(n31962), .S0(op_i_23__N_1154_adj_7371[16]), 
          .S1(op_i_23__N_1154_adj_7371[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_19.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_19.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_17 (.A0(n31492), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[14]), .A1(n31490), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[15]), .CIN(n31960), .COUT(n31961), .S0(op_i_23__N_1154_adj_7371[14]), 
          .S1(op_i_23__N_1154_adj_7371[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_17.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_17.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_15 (.A0(n31496), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[12]), .A1(n31494), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[13]), .CIN(n31959), .COUT(n31960), .S0(op_i_23__N_1154_adj_7371[12]), 
          .S1(op_i_23__N_1154_adj_7371[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_15.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_15.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_13 (.A0(n31500), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[10]), .A1(n31498), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[11]), .CIN(n31958), .COUT(n31959), .S0(op_i_23__N_1154_adj_7371[10]), 
          .S1(op_i_23__N_1154_adj_7371[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_13.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_13.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_11 (.A0(n31504), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[8]), .A1(n31502), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[9]), .CIN(n31957), .COUT(n31958), .S0(op_i_23__N_1154_adj_7371[8]), 
          .S1(op_i_23__N_1154_adj_7371[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_11.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_11.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_9 (.A0(n31508), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[6]), .A1(n31506), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[7]), .CIN(n31956), .COUT(n31957), .S0(op_i_23__N_1154_adj_7371[6]), 
          .S1(op_i_23__N_1154_adj_7371[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_9.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_9.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_7 (.A0(n31512), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[4]), .A1(n31510), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[5]), .CIN(n31955), .COUT(n31956), .S0(op_i_23__N_1154_adj_7371[4]), 
          .S1(op_i_23__N_1154_adj_7371[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_7.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_7.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_5 (.A0(n31516), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[2]), .A1(n31514), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[3]), .CIN(n31954), .COUT(n31955), .S0(op_i_23__N_1154_adj_7371[2]), 
          .S1(op_i_23__N_1154_adj_7371[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_5.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_5.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_3 (.A0(n31520), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_i[0]), .A1(n31518), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_i[1]), .CIN(n31953), .COUT(n31954), .S0(op_i_23__N_1154_adj_7371[0]), 
          .S1(op_i_23__N_1154_adj_7371[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_3.INIT0 = 16'h65aa;
    defparam _add_1_1031_add_4_3.INIT1 = 16'h65aa;
    defparam _add_1_1031_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1031_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(rom4_state[0]), .B1(n29826), .C1(n29827), 
          .D1(n29828), .COUT(n31953));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1031_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1031_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1031_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1031_add_4_1.INJECT1_1 = "NO";
    LUT4 i7537_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[391])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7537_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1023_add_4_26 (.A0(shift_4_dout_i[23]), .B0(shift_4_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31949), .S0(n319_adj_6714));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1023_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_24 (.A0(shift_4_dout_i[22]), .B0(shift_4_dout_r[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[23]), .B1(shift_4_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31948), .COUT(n31949), .S0(n10734), 
          .S1(n10735));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_22 (.A0(shift_4_dout_i[20]), .B0(shift_4_dout_r[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[21]), .B1(shift_4_dout_r[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31947), .COUT(n31948), .S0(n10732), 
          .S1(n10733));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_20 (.A0(shift_4_dout_i[18]), .B0(shift_4_dout_r[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[19]), .B1(shift_4_dout_r[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31946), .COUT(n31947), .S0(n10730), 
          .S1(n10731));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_18 (.A0(shift_4_dout_i[16]), .B0(shift_4_dout_r[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[17]), .B1(shift_4_dout_r[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31945), .COUT(n31946), .S0(n10728), 
          .S1(n10729));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_16 (.A0(shift_4_dout_i[14]), .B0(shift_4_dout_r[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[15]), .B1(shift_4_dout_r[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31944), .COUT(n31945), .S0(n10726), 
          .S1(n10727));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_14 (.A0(shift_4_dout_i[12]), .B0(shift_4_dout_r[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[13]), .B1(shift_4_dout_r[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31943), .COUT(n31944), .S0(n10724), 
          .S1(n10725));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_12 (.A0(shift_4_dout_i[10]), .B0(shift_4_dout_r[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[11]), .B1(shift_4_dout_r[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31942), .COUT(n31943), .S0(n10722), 
          .S1(n10723));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_10 (.A0(shift_4_dout_i[8]), .B0(shift_4_dout_r[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[9]), .B1(shift_4_dout_r[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31941), .COUT(n31942), .S0(n10720), 
          .S1(n10721));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_8 (.A0(shift_4_dout_i[6]), .B0(shift_4_dout_r[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[7]), .B1(shift_4_dout_r[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31940), .COUT(n31941), .S0(n10718), 
          .S1(n10719));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_6 (.A0(shift_4_dout_i[4]), .B0(shift_4_dout_r[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[5]), .B1(shift_4_dout_r[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31939), .COUT(n31940), .S0(n114_adj_7263), 
          .S1(n111_adj_7262));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_6.INJECT1_1 = "NO";
    LUT4 i15842_3_lut (.A(\result_r[16] [1]), .B(\result_r[17] [1]), .C(y_1_delay[0]), 
         .Z(n34226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15842_3_lut.init = 16'hcaca;
    LUT4 i14942_3_lut (.A(\result_i[14] [15]), .B(\result_i[15] [15]), .C(y_1_delay[0]), 
         .Z(n33326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14942_3_lut.init = 16'hcaca;
    LUT4 i7529_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[392])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7529_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15667 (.BLUT(n34038), .ALUT(n34039), .C0(y_1_delay[1]), .Z(n34051));
    LUT4 i870_4_lut_rep_441 (.A(count_y[4]), .B(n34771), .C(n34770), .D(count_y[3]), 
         .Z(n34811)) /* synthesis lut_function=(A ((C+(D))+!B)+!A !((C+(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i870_4_lut_rep_441.init = 16'haaa6;
    LUT4 i7521_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[393])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7521_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7513_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[394])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7513_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7505_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[395])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7505_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15841_3_lut (.A(\result_r[14] [1]), .B(\result_r[15] [1]), .C(y_1_delay[0]), 
         .Z(n34225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15841_3_lut.init = 16'hcaca;
    PFUMX i15483 (.BLUT(n33856), .ALUT(n33857), .C0(y_1_delay[1]), .Z(n33867));
    LUT4 i7497_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[396])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7497_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15840_3_lut (.A(\result_r[12] [1]), .B(\result_r[13] [1]), .C(y_1_delay[0]), 
         .Z(n34224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15840_3_lut.init = 16'hcaca;
    LUT4 i7489_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[397])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7489_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7481_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[398])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7481_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7473_3_lut_4_lut (.A(n34717), .B(n34704), .C(\result_r[7] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[399])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7473_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3633_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[368])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3633_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15839_3_lut (.A(\result_r[10] [1]), .B(\result_r[11] [1]), .C(y_1_delay[0]), 
         .Z(n34223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15839_3_lut.init = 16'hcaca;
    LUT4 i3625_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[369])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3625_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15761 (.BLUT(n34133), .ALUT(n34134), .C0(y_1_delay[1]), .Z(n34145));
    LUT4 i3617_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[370])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3617_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3609_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[371])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3609_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3601_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[372])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3601_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15838_3_lut (.A(\result_r[8] [1]), .B(\result_r[9] [1]), .C(y_1_delay[0]), 
         .Z(n34222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15838_3_lut.init = 16'hcaca;
    LUT4 i3593_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[373])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3593_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15668 (.BLUT(n34040), .ALUT(n34041), .C0(y_1_delay[1]), .Z(n34052));
    LUT4 i3585_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[374])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3585_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15484 (.BLUT(n33858), .ALUT(n33859), .C0(y_1_delay[1]), .Z(n33868));
    LUT4 i3577_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[375])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3577_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3569_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[376])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3569_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3561_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[377])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3561_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3553_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[378])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3553_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15837_3_lut (.A(\result_r[6] [1]), .B(\result_r[7] [1]), .C(y_1_delay[0]), 
         .Z(n34221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15837_3_lut.init = 16'hcaca;
    LUT4 i3545_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[379])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3545_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3537_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[380])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3537_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3529_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[381])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3529_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15485 (.BLUT(n33860), .ALUT(n33861), .C0(y_1_delay[1]), .Z(n33869));
    LUT4 i3521_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[382])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3521_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15836_3_lut (.A(\result_r[4] [1]), .B(\result_r[5] [1]), .C(y_1_delay[0]), 
         .Z(n34220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15836_3_lut.init = 16'hcaca;
    LUT4 i3513_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_i[8] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[383])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3513_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7721_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[368])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7721_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7713_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[369])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7713_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7705_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[370])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7705_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15762 (.BLUT(n34135), .ALUT(n34136), .C0(y_1_delay[1]), .Z(n34146));
    LUT4 i7697_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[371])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7697_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7689_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[372])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7689_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7681_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[373])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7681_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7673_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[374])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7673_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15835_3_lut (.A(\result_r[2] [1]), .B(\result_r[3] [1]), .C(y_1_delay[0]), 
         .Z(n34219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15835_3_lut.init = 16'hcaca;
    LUT4 i7665_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[375])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7665_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7657_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[376])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7657_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7649_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[377])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7649_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15669 (.BLUT(n34042), .ALUT(n34043), .C0(y_1_delay[1]), .Z(n34053));
    PFUMX i15175 (.BLUT(n33550), .ALUT(n33551), .C0(y_1_delay[1]), .Z(n33559));
    LUT4 i7641_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[378])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7641_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7633_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[379])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7633_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7625_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[380])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7625_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7617_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[381])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7617_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15834_3_lut (.A(\result_r[0] [1]), .B(\result_r[1] [1]), .C(y_1_delay[0]), 
         .Z(n34218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15834_3_lut.init = 16'hcaca;
    LUT4 i7609_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[382])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7609_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7601_3_lut_4_lut (.A(n34717), .B(n34705), .C(\result_r[8] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[383])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7601_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3761_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[352])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3761_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3753_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[353])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3753_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3745_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[354])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3745_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3737_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[355])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3737_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3729_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[356])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3729_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3721_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[357])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3721_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3713_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[358])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3713_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3705_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[359])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3705_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3697_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[360])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3697_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3689_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[361])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3689_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3681_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[362])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3681_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15763 (.BLUT(n34137), .ALUT(n34138), .C0(y_1_delay[1]), .Z(n34147));
    LUT4 i3673_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[363])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3673_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3665_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[364])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3665_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3657_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[365])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3657_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3649_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[366])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3649_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14069_2_lut (.A(shift_8_dout_i[0]), .B(shift_8_dout_r[0]), .Z(n11148)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14069_2_lut.init = 16'h6666;
    LUT4 i3641_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_i[9] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[367])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3641_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15198_3_lut (.A(\result_i[30] [7]), .B(\result_i[31] [7]), .C(y_1_delay[0]), 
         .Z(n33582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15198_3_lut.init = 16'hcaca;
    LUT4 i15197_3_lut (.A(\result_i[28] [7]), .B(\result_i[29] [7]), .C(y_1_delay[0]), 
         .Z(n33581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15197_3_lut.init = 16'hcaca;
    LUT4 i7849_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[352])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7849_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7841_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[353])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7841_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7833_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[354])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7833_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15539_3_lut (.A(\result_r[30] [11]), .B(\result_r[31] [11]), .C(y_1_delay[0]), 
         .Z(n33923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15539_3_lut.init = 16'hcaca;
    LUT4 i7825_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[355])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7825_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15538_3_lut (.A(\result_r[28] [11]), .B(\result_r[29] [11]), .C(y_1_delay[0]), 
         .Z(n33922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15538_3_lut.init = 16'hcaca;
    LUT4 i15287_3_lut (.A(\result_i[22] [4]), .B(\result_i[23] [4]), .C(y_1_delay[0]), 
         .Z(n33671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15287_3_lut.init = 16'hcaca;
    LUT4 i7817_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[356])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7817_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7809_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[357])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7809_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15196_3_lut (.A(\result_i[26] [7]), .B(\result_i[27] [7]), .C(y_1_delay[0]), 
         .Z(n33580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15196_3_lut.init = 16'hcaca;
    LUT4 i15195_3_lut (.A(\result_i[24] [7]), .B(\result_i[25] [7]), .C(y_1_delay[0]), 
         .Z(n33579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15195_3_lut.init = 16'hcaca;
    LUT4 i7801_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[358])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7801_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15286_3_lut (.A(\result_i[20] [4]), .B(\result_i[21] [4]), .C(y_1_delay[0]), 
         .Z(n33670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15286_3_lut.init = 16'hcaca;
    LUT4 i7793_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[359])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7793_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7785_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[360])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7785_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15194_3_lut (.A(\result_i[22] [7]), .B(\result_i[23] [7]), .C(y_1_delay[0]), 
         .Z(n33578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15194_3_lut.init = 16'hcaca;
    LUT4 i7777_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[361])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7777_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1023_add_4_4 (.A0(shift_4_dout_i[2]), .B0(shift_4_dout_r[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[3]), .B1(shift_4_dout_r[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31938), .COUT(n31939), .S0(n120_adj_7265), 
          .S1(n117_adj_7264));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_2 (.A0(shift_4_dout_i[0]), .B0(shift_4_dout_r[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[1]), .B1(shift_4_dout_r[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n31938), .S1(n123_adj_7266));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1023_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1023_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1023_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_26 (.A0(op_r_23__N_1106_adj_7370[23]), .B0(n34841), 
          .C0(shift_2_dout_r[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n31936), .S0(delay_r_23__N_1178_adj_7427[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_26.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1116_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_24 (.A0(op_r_23__N_1106_adj_7370[21]), .B0(n34841), 
          .C0(shift_2_dout_r[21]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[22]), 
          .B1(n34841), .C1(shift_2_dout_r[22]), .D1(VCC_net), .CIN(n31935), 
          .COUT(n31936), .S0(delay_r_23__N_1178_adj_7427[21]), .S1(delay_r_23__N_1178_adj_7427[22]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_24.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_24.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_22 (.A0(op_r_23__N_1106_adj_7370[19]), .B0(n34841), 
          .C0(shift_2_dout_r[19]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[20]), 
          .B1(n34841), .C1(shift_2_dout_r[20]), .D1(VCC_net), .CIN(n31934), 
          .COUT(n31935), .S0(delay_r_23__N_1178_adj_7427[19]), .S1(delay_r_23__N_1178_adj_7427[20]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_22.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_22.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_20 (.A0(op_r_23__N_1106_adj_7370[17]), .B0(n34841), 
          .C0(shift_2_dout_r[17]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[18]), 
          .B1(n34841), .C1(shift_2_dout_r[18]), .D1(VCC_net), .CIN(n31933), 
          .COUT(n31934), .S0(delay_r_23__N_1178_adj_7427[17]), .S1(delay_r_23__N_1178_adj_7427[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_20.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_20.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_18 (.A0(op_r_23__N_1106_adj_7370[15]), .B0(n34841), 
          .C0(shift_2_dout_r[15]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[16]), 
          .B1(n34841), .C1(shift_2_dout_r[16]), .D1(VCC_net), .CIN(n31932), 
          .COUT(n31933), .S0(delay_r_23__N_1178_adj_7427[15]), .S1(delay_r_23__N_1178_adj_7427[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_18.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_18.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_16 (.A0(op_r_23__N_1106_adj_7370[13]), .B0(n34841), 
          .C0(shift_2_dout_r[13]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[14]), 
          .B1(n34841), .C1(shift_2_dout_r[14]), .D1(VCC_net), .CIN(n31931), 
          .COUT(n31932), .S0(delay_r_23__N_1178_adj_7427[13]), .S1(delay_r_23__N_1178_adj_7427[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_16.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_16.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_14 (.A0(op_r_23__N_1106_adj_7370[11]), .B0(n34841), 
          .C0(shift_2_dout_r[11]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[12]), 
          .B1(n34841), .C1(shift_2_dout_r[12]), .D1(VCC_net), .CIN(n31930), 
          .COUT(n31931), .S0(delay_r_23__N_1178_adj_7427[11]), .S1(delay_r_23__N_1178_adj_7427[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_14.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_14.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_12 (.A0(op_r_23__N_1106_adj_7370[9]), .B0(n34841), 
          .C0(shift_2_dout_r[9]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[10]), 
          .B1(n34841), .C1(shift_2_dout_r[10]), .D1(VCC_net), .CIN(n31929), 
          .COUT(n31930), .S0(delay_r_23__N_1178_adj_7427[9]), .S1(delay_r_23__N_1178_adj_7427[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_12.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_12.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_10 (.A0(op_r_23__N_1106_adj_7370[7]), .B0(n34841), 
          .C0(shift_2_dout_r[7]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[8]), 
          .B1(n34841), .C1(shift_2_dout_r[8]), .D1(VCC_net), .CIN(n31928), 
          .COUT(n31929), .S0(delay_r_23__N_1178_adj_7427[7]), .S1(delay_r_23__N_1178_adj_7427[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_10.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_10.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_8 (.A0(op_r_23__N_1106_adj_7370[5]), .B0(n34841), 
          .C0(shift_2_dout_r[5]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[6]), 
          .B1(n34841), .C1(shift_2_dout_r[6]), .D1(VCC_net), .CIN(n31927), 
          .COUT(n31928), .S0(delay_r_23__N_1178_adj_7427[5]), .S1(delay_r_23__N_1178_adj_7427[6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_8.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_8.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_6 (.A0(op_r_23__N_1106_adj_7370[3]), .B0(n34841), 
          .C0(shift_2_dout_r[3]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[4]), 
          .B1(n34841), .C1(shift_2_dout_r[4]), .D1(VCC_net), .CIN(n31926), 
          .COUT(n31927), .S0(delay_r_23__N_1178_adj_7427[3]), .S1(delay_r_23__N_1178_adj_7427[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_6.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_6.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_4 (.A0(op_r_23__N_1106_adj_7370[1]), .B0(n34841), 
          .C0(shift_2_dout_r[1]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[2]), 
          .B1(n34841), .C1(shift_2_dout_r[2]), .D1(VCC_net), .CIN(n31925), 
          .COUT(n31926), .S0(delay_r_23__N_1178_adj_7427[1]), .S1(delay_r_23__N_1178_adj_7427[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_4.INIT0 = 16'h8787;
    defparam _add_1_1116_add_4_4.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1116_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(op_r_23__N_1106_adj_7370[0]), .B1(n34841), 
          .C1(shift_2_dout_r[0]), .D1(VCC_net), .COUT(n31925), .S1(delay_r_23__N_1178_adj_7427[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1116_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1116_add_4_2.INIT1 = 16'h8787;
    defparam _add_1_1116_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1116_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1143_add_4_12 (.A0(rom8_w_r[10]), .B0(n6_adj_7292), .C0(n5), 
          .D0(n34726), .A1(rom8_w_r[10]), .B1(n6_adj_7292), .C1(n5), 
          .D1(n34726), .CIN(n31923), .S0(n12453), .S1(n119));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1143_add_4_12.INIT0 = 16'h95aa;
    defparam _add_1_1143_add_4_12.INIT1 = 16'h95aa;
    defparam _add_1_1143_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1143_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1143_add_4_10 (.A0(n34761), .B0(n34760), .C0(s_count[3]), 
          .D0(n34752), .A1(n34754), .B1(n5), .C1(n6_adj_7292), .D1(n34726), 
          .CIN(n31922), .COUT(n31923), .S0(n12451), .S1(n12452));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1143_add_4_10.INIT0 = 16'h22d2;
    defparam _add_1_1143_add_4_10.INIT1 = 16'h6a55;
    defparam _add_1_1143_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1143_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1143_add_4_8 (.A0(s_count[1]), .B0(s_count[0]), .C0(s_count[2]), 
          .D0(s_count[3]), .A1(rom8_w_r[6]), .B1(n34788), .C1(n34787), 
          .D1(n29782), .CIN(n31921), .COUT(n31922), .S0(n12449), .S1(n12450));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1143_add_4_8.INIT0 = 16'hf1ff;
    defparam _add_1_1143_add_4_8.INIT1 = 16'h559a;
    defparam _add_1_1143_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1143_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1143_add_4_6 (.A0(rom8_w_r[3]), .B0(n34760), .C0(n34761), 
          .D0(n34762), .A1(n30191), .B1(n34742), .C1(s_count[3]), .D1(n34753), 
          .CIN(n31920), .COUT(n31921), .S0(n12447), .S1(n12448));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1143_add_4_6.INIT0 = 16'h9aaa;
    defparam _add_1_1143_add_4_6.INIT1 = 16'h8878;
    defparam _add_1_1143_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1143_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1143_add_4_4 (.A0(n30191), .B0(n34734), .C0(s_count[3]), 
          .D0(n34779), .A1(n34761), .B1(n34760), .C1(s_count[3]), .D1(n34752), 
          .CIN(n31919), .COUT(n31920), .S0(n12445), .S1(n12446));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1143_add_4_4.INIT0 = 16'h7888;
    defparam _add_1_1143_add_4_4.INIT1 = 16'h22d2;
    defparam _add_1_1143_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1143_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1143_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n30191), .B1(n34762), .C1(s_count[3]), .D1(n34778), 
          .COUT(n31919), .S1(n12444));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1143_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1143_add_4_2.INIT1 = 16'h7888;
    defparam _add_1_1143_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1143_add_4_2.INJECT1_1 = "NO";
    LUT4 i7769_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[362])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7769_3_lut_4_lut.init = 16'hf1e0;
    CCU2C _add_1_1026_add_4_25 (.A0(n31427), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[22]), .A1(n31425), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[23]), .CIN(n31917), .S0(op_r_23__N_1106_adj_7370[22]), 
          .S1(op_r_23__N_1106_adj_7370[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_25.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_25.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_23 (.A0(n31431), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[20]), .A1(n31429), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[21]), .CIN(n31916), .COUT(n31917), .S0(op_r_23__N_1106_adj_7370[20]), 
          .S1(op_r_23__N_1106_adj_7370[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_23.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_23.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_21 (.A0(n31435), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[18]), .A1(n31433), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[19]), .CIN(n31915), .COUT(n31916), .S0(op_r_23__N_1106_adj_7370[18]), 
          .S1(op_r_23__N_1106_adj_7370[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_21.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_21.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_19 (.A0(n31439), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[16]), .A1(n31437), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[17]), .CIN(n31914), .COUT(n31915), .S0(op_r_23__N_1106_adj_7370[16]), 
          .S1(op_r_23__N_1106_adj_7370[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_19.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_19.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_17 (.A0(n31443), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[14]), .A1(n31441), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[15]), .CIN(n31913), .COUT(n31914), .S0(op_r_23__N_1106_adj_7370[14]), 
          .S1(op_r_23__N_1106_adj_7370[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_17.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_17.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_15 (.A0(n31447), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[12]), .A1(n31445), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[13]), .CIN(n31912), .COUT(n31913), .S0(op_r_23__N_1106_adj_7370[12]), 
          .S1(op_r_23__N_1106_adj_7370[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_15.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_15.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_13 (.A0(n31451), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[10]), .A1(n31449), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[11]), .CIN(n31911), .COUT(n31912), .S0(op_r_23__N_1106_adj_7370[10]), 
          .S1(op_r_23__N_1106_adj_7370[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_13.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_13.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_11 (.A0(n31455), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[8]), .A1(n31453), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[9]), .CIN(n31910), .COUT(n31911), .S0(op_r_23__N_1106_adj_7370[8]), 
          .S1(op_r_23__N_1106_adj_7370[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_11.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_11.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_9 (.A0(n31459), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[6]), .A1(n31457), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[7]), .CIN(n31909), .COUT(n31910), .S0(op_r_23__N_1106_adj_7370[6]), 
          .S1(op_r_23__N_1106_adj_7370[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_9.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_9.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_7 (.A0(n31463), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[4]), .A1(n31461), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[5]), .CIN(n31908), .COUT(n31909), .S0(op_r_23__N_1106_adj_7370[4]), 
          .S1(op_r_23__N_1106_adj_7370[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_7.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_7.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_5 (.A0(n31467), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[2]), .A1(n31465), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[3]), .CIN(n31907), .COUT(n31908), .S0(op_r_23__N_1106_adj_7370[2]), 
          .S1(op_r_23__N_1106_adj_7370[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_5.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_5.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_3 (.A0(n31471), .B0(rom4_state[0]), .C0(n34799), 
          .D0(shift_4_dout_r[0]), .A1(n31469), .B1(rom4_state[0]), .C1(n34799), 
          .D1(shift_4_dout_r[1]), .CIN(n31906), .COUT(n31907), .S0(op_r_23__N_1106_adj_7370[0]), 
          .S1(op_r_23__N_1106_adj_7370[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_3.INIT0 = 16'h65aa;
    defparam _add_1_1026_add_4_3.INIT1 = 16'h65aa;
    defparam _add_1_1026_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1026_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n34520), .B1(n29819), .C1(n29820), .D1(n34799), 
          .COUT(n31906));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1026_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1026_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1026_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1026_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_26 (.A0(shift_4_dout_i[23]), .B0(shift_4_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[23]), .B1(shift_4_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31901), .S0(n12263), .S1(n12264));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_24 (.A0(shift_4_dout_i[21]), .B0(shift_4_dout_r[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[22]), .B1(shift_4_dout_r[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31900), .COUT(n31901), .S0(n12261), 
          .S1(n12262));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_22 (.A0(shift_4_dout_i[19]), .B0(shift_4_dout_r[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[20]), .B1(shift_4_dout_r[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31899), .COUT(n31900), .S0(n12259), 
          .S1(n12260));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_20 (.A0(shift_4_dout_i[17]), .B0(shift_4_dout_r[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[18]), .B1(shift_4_dout_r[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31898), .COUT(n31899), .S0(n12257), 
          .S1(n12258));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_18 (.A0(shift_4_dout_i[15]), .B0(shift_4_dout_r[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[16]), .B1(shift_4_dout_r[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31897), .COUT(n31898), .S0(n12255), 
          .S1(n12256));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_16 (.A0(shift_4_dout_i[13]), .B0(shift_4_dout_r[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[14]), .B1(shift_4_dout_r[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31896), .COUT(n31897), .S0(n12253), 
          .S1(n12254));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_14 (.A0(shift_4_dout_i[11]), .B0(shift_4_dout_r[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[12]), .B1(shift_4_dout_r[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31895), .COUT(n31896), .S0(n12251), 
          .S1(n12252));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_12 (.A0(shift_4_dout_i[9]), .B0(shift_4_dout_r[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[10]), .B1(shift_4_dout_r[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31894), .COUT(n31895), .S0(n12249), 
          .S1(n12250));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_10 (.A0(shift_4_dout_i[7]), .B0(shift_4_dout_r[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[8]), .B1(shift_4_dout_r[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31893), .COUT(n31894), .S0(n12247), 
          .S1(n12248));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_8 (.A0(shift_4_dout_i[5]), .B0(shift_4_dout_r[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[6]), .B1(shift_4_dout_r[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31892), .COUT(n31893), .S0(n12245), 
          .S1(n12246));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_6 (.A0(shift_4_dout_i[3]), .B0(shift_4_dout_r[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[4]), .B1(shift_4_dout_r[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31891), .COUT(n31892), .S0(n12243), 
          .S1(n12244));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_4 (.A0(shift_4_dout_i[1]), .B0(shift_4_dout_r[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_4_dout_i[2]), .B1(shift_4_dout_r[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31890), .COUT(n31891), .S0(n12241), 
          .S1(n12242));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1119_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1119_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(shift_4_dout_i[0]), .B1(shift_4_dout_r[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n31890), .S1(n12240));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1119_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1119_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1119_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1119_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_32 (.A0(op_r_23__N_1268_adj_7375[30]), .B0(op_i_23__N_1310_adj_7380[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[31]), 
          .B1(op_i_23__N_1310_adj_7380[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31888), .S0(op_i_23__N_1130_adj_7381[30]), .S1(op_i_23__N_1130_adj_7381[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_30 (.A0(op_r_23__N_1268_adj_7375[28]), .B0(op_i_23__N_1310_adj_7380[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[29]), 
          .B1(op_i_23__N_1310_adj_7380[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31887), .COUT(n31888), .S0(op_i_23__N_1130_adj_7381[28]), 
          .S1(op_i_23__N_1130_adj_7381[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_28 (.A0(op_r_23__N_1268_adj_7375[26]), .B0(op_i_23__N_1310_adj_7380[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[27]), 
          .B1(op_i_23__N_1310_adj_7380[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31886), .COUT(n31887), .S0(op_i_23__N_1130_adj_7381[26]), 
          .S1(op_i_23__N_1130_adj_7381[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_26 (.A0(op_r_23__N_1268_adj_7375[24]), .B0(op_i_23__N_1310_adj_7380[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[25]), 
          .B1(op_i_23__N_1310_adj_7380[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31885), .COUT(n31886), .S0(op_i_23__N_1130_adj_7381[24]), 
          .S1(op_i_23__N_1130_adj_7381[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_24 (.A0(op_r_23__N_1268_adj_7375[22]), .B0(op_i_23__N_1310_adj_7380[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[23]), 
          .B1(op_i_23__N_1310_adj_7380[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31884), .COUT(n31885), .S0(op_i_23__N_1130_adj_7381[22]), 
          .S1(op_i_23__N_1130_adj_7381[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_22 (.A0(op_r_23__N_1268_adj_7375[20]), .B0(op_i_23__N_1310_adj_7380[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[21]), 
          .B1(op_i_23__N_1310_adj_7380[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31883), .COUT(n31884), .S0(op_i_23__N_1130_adj_7381[20]), 
          .S1(op_i_23__N_1130_adj_7381[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_20 (.A0(op_r_23__N_1268_adj_7375[18]), .B0(op_i_23__N_1310_adj_7380[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[19]), 
          .B1(op_i_23__N_1310_adj_7380[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31882), .COUT(n31883), .S0(op_i_23__N_1130_adj_7381[18]), 
          .S1(op_i_23__N_1130_adj_7381[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_18 (.A0(op_r_23__N_1268_adj_7375[16]), .B0(op_i_23__N_1310_adj_7380[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[17]), 
          .B1(op_i_23__N_1310_adj_7380[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31881), .COUT(n31882), .S0(op_i_23__N_1130_adj_7381[16]), 
          .S1(op_i_23__N_1130_adj_7381[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_16 (.A0(op_r_23__N_1268_adj_7375[14]), .B0(op_i_23__N_1310_adj_7380[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[15]), 
          .B1(op_i_23__N_1310_adj_7380[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31880), .COUT(n31881), .S0(op_i_23__N_1130_adj_7381[14]), 
          .S1(op_i_23__N_1130_adj_7381[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_14 (.A0(op_r_23__N_1268_adj_7375[12]), .B0(op_i_23__N_1310_adj_7380[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[13]), 
          .B1(op_i_23__N_1310_adj_7380[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31879), .COUT(n31880), .S0(op_i_23__N_1130_adj_7381[12]), 
          .S1(op_i_23__N_1130_adj_7381[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_12 (.A0(op_r_23__N_1268_adj_7375[10]), .B0(op_i_23__N_1310_adj_7380[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[11]), 
          .B1(op_i_23__N_1310_adj_7380[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31878), .COUT(n31879), .S0(op_i_23__N_1130_adj_7381[10]), 
          .S1(op_i_23__N_1130_adj_7381[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_10 (.A0(op_r_23__N_1268_adj_7375[8]), .B0(op_i_23__N_1310_adj_7380[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[9]), 
          .B1(op_i_23__N_1310_adj_7380[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31877), .COUT(n31878), .S0(op_i_23__N_1130_adj_7381[8]), 
          .S1(op_i_23__N_1130_adj_7381[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_8 (.A0(op_r_23__N_1268_adj_7375[6]), .B0(op_i_23__N_1310_adj_7380[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[7]), 
          .B1(op_i_23__N_1310_adj_7380[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31876), .COUT(n31877));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_6 (.A0(op_r_23__N_1268_adj_7375[4]), .B0(op_i_23__N_1310_adj_7380[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[5]), 
          .B1(op_i_23__N_1310_adj_7380[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31875), .COUT(n31876));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_4 (.A0(op_r_23__N_1268_adj_7375[2]), .B0(op_i_23__N_1310_adj_7380[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[3]), 
          .B1(op_i_23__N_1310_adj_7380[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31874), .COUT(n31875));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1034_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_2 (.A0(op_r_23__N_1268_adj_7375[0]), .B0(op_i_23__N_1310_adj_7380[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[1]), 
          .B1(op_i_23__N_1310_adj_7380[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n31874));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1034_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1034_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1034_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_26 (.A0(shift_8_dout_i[23]), .B0(shift_8_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[23]), .B1(shift_8_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31872), .S0(n12293), .S1(n12294));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_24 (.A0(shift_8_dout_i[21]), .B0(shift_8_dout_r[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[22]), .B1(shift_8_dout_r[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31871), .COUT(n31872), .S0(n12291), 
          .S1(n12292));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_22 (.A0(shift_8_dout_i[19]), .B0(shift_8_dout_r[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[20]), .B1(shift_8_dout_r[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31870), .COUT(n31871), .S0(n12289), 
          .S1(n12290));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_20 (.A0(shift_8_dout_i[17]), .B0(shift_8_dout_r[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[18]), .B1(shift_8_dout_r[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31869), .COUT(n31870), .S0(n12287), 
          .S1(n12288));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_18 (.A0(shift_8_dout_i[15]), .B0(shift_8_dout_r[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[16]), .B1(shift_8_dout_r[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31868), .COUT(n31869), .S0(n12285), 
          .S1(n12286));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_16 (.A0(shift_8_dout_i[13]), .B0(shift_8_dout_r[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[14]), .B1(shift_8_dout_r[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31867), .COUT(n31868), .S0(n12283), 
          .S1(n12284));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_14 (.A0(shift_8_dout_i[11]), .B0(shift_8_dout_r[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[12]), .B1(shift_8_dout_r[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31866), .COUT(n31867), .S0(n12281), 
          .S1(n12282));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_12 (.A0(shift_8_dout_i[9]), .B0(shift_8_dout_r[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[10]), .B1(shift_8_dout_r[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31865), .COUT(n31866), .S0(n12279), 
          .S1(n12280));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_10 (.A0(shift_8_dout_i[7]), .B0(shift_8_dout_r[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[8]), .B1(shift_8_dout_r[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31864), .COUT(n31865), .S0(n12277), 
          .S1(n12278));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_8 (.A0(shift_8_dout_i[5]), .B0(shift_8_dout_r[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[6]), .B1(shift_8_dout_r[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31863), .COUT(n31864), .S0(n12275), 
          .S1(n12276));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_6 (.A0(shift_8_dout_i[3]), .B0(shift_8_dout_r[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[4]), .B1(shift_8_dout_r[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31862), .COUT(n31863), .S0(n12273), 
          .S1(n12274));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_4 (.A0(shift_8_dout_i[1]), .B0(shift_8_dout_r[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_8_dout_i[2]), .B1(shift_8_dout_r[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31861), .COUT(n31862), .S0(n12271), 
          .S1(n12272));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1122_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1122_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(shift_8_dout_i[0]), .B1(shift_8_dout_r[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n31861), .S1(n12270));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1122_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1122_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1122_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1122_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_25 (.A0(n31378), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[22]), .A1(n31376), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[23]), .CIN(n31859), .S0(op_i_23__N_1154_adj_7320[22]), 
          .S1(op_i_23__N_1154_adj_7320[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_25.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_25.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_23 (.A0(n31382), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[20]), .A1(n31380), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[21]), .CIN(n31858), .COUT(n31859), .S0(op_i_23__N_1154_adj_7320[20]), 
          .S1(op_i_23__N_1154_adj_7320[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_23.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_23.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_21 (.A0(n31386), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[18]), .A1(n31384), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[19]), .CIN(n31857), .COUT(n31858), .S0(op_i_23__N_1154_adj_7320[18]), 
          .S1(op_i_23__N_1154_adj_7320[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_21.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_21.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_19 (.A0(n31390), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[16]), .A1(n31388), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[17]), .CIN(n31856), .COUT(n31857), .S0(op_i_23__N_1154_adj_7320[16]), 
          .S1(op_i_23__N_1154_adj_7320[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_19.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_19.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_17 (.A0(n31394), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[14]), .A1(n31392), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[15]), .CIN(n31855), .COUT(n31856), .S0(op_i_23__N_1154_adj_7320[14]), 
          .S1(op_i_23__N_1154_adj_7320[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_17.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_17.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_15 (.A0(n31398), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[12]), .A1(n31396), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[13]), .CIN(n31854), .COUT(n31855), .S0(op_i_23__N_1154_adj_7320[12]), 
          .S1(op_i_23__N_1154_adj_7320[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_15.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_15.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_13 (.A0(n31402), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[10]), .A1(n31400), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[11]), .CIN(n31853), .COUT(n31854), .S0(op_i_23__N_1154_adj_7320[10]), 
          .S1(op_i_23__N_1154_adj_7320[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_13.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_13.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_11 (.A0(n31406), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[8]), .A1(n31404), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[9]), .CIN(n31852), .COUT(n31853), .S0(op_i_23__N_1154_adj_7320[8]), 
          .S1(op_i_23__N_1154_adj_7320[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_11.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_11.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_9 (.A0(n31410), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[6]), .A1(n31408), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[7]), .CIN(n31851), .COUT(n31852), .S0(op_i_23__N_1154_adj_7320[6]), 
          .S1(op_i_23__N_1154_adj_7320[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_9.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_9.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_7 (.A0(n31414), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[4]), .A1(n31412), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[5]), .CIN(n31850), .COUT(n31851), .S0(op_i_23__N_1154_adj_7320[4]), 
          .S1(op_i_23__N_1154_adj_7320[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_7.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_7.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_5 (.A0(n31418), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[2]), .A1(n31416), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[3]), .CIN(n31849), .COUT(n31850), .S0(op_i_23__N_1154_adj_7320[2]), 
          .S1(op_i_23__N_1154_adj_7320[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_5.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_5.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_3 (.A0(n31422), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_i[0]), .A1(n31420), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_i[1]), .CIN(n31848), .COUT(n31849), .S0(op_i_23__N_1154_adj_7320[0]), 
          .S1(op_i_23__N_1154_adj_7320[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_3.INIT0 = 16'h65aa;
    defparam _add_1_1009_add_4_3.INIT1 = 16'h65aa;
    defparam _add_1_1009_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1009_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n34532), .B1(n29815), .C1(n29816), .D1(n34794), 
          .COUT(n31848));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1009_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1009_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1009_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1009_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_32 (.A0(op_r_23__N_1268_adj_7375[30]), .B0(op_r_23__N_1226_adj_7377[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[31]), 
          .B1(op_r_23__N_1226_adj_7377[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31843), .S0(op_r_23__N_1082_adj_7378[30]), .S1(op_r_23__N_1082_adj_7378[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_30 (.A0(op_r_23__N_1268_adj_7375[28]), .B0(op_r_23__N_1226_adj_7377[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[29]), 
          .B1(op_r_23__N_1226_adj_7377[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31842), .COUT(n31843), .S0(op_r_23__N_1082_adj_7378[28]), 
          .S1(op_r_23__N_1082_adj_7378[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_28 (.A0(op_r_23__N_1268_adj_7375[26]), .B0(op_r_23__N_1226_adj_7377[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[27]), 
          .B1(op_r_23__N_1226_adj_7377[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31841), .COUT(n31842), .S0(op_r_23__N_1082_adj_7378[26]), 
          .S1(op_r_23__N_1082_adj_7378[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_26 (.A0(op_r_23__N_1268_adj_7375[24]), .B0(op_r_23__N_1226_adj_7377[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[25]), 
          .B1(op_r_23__N_1226_adj_7377[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31840), .COUT(n31841), .S0(op_r_23__N_1082_adj_7378[24]), 
          .S1(op_r_23__N_1082_adj_7378[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_24 (.A0(op_r_23__N_1268_adj_7375[22]), .B0(op_r_23__N_1226_adj_7377[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[23]), 
          .B1(op_r_23__N_1226_adj_7377[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31839), .COUT(n31840), .S0(op_r_23__N_1082_adj_7378[22]), 
          .S1(op_r_23__N_1082_adj_7378[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_22 (.A0(op_r_23__N_1268_adj_7375[20]), .B0(op_r_23__N_1226_adj_7377[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[21]), 
          .B1(op_r_23__N_1226_adj_7377[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31838), .COUT(n31839), .S0(op_r_23__N_1082_adj_7378[20]), 
          .S1(op_r_23__N_1082_adj_7378[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_20 (.A0(op_r_23__N_1268_adj_7375[18]), .B0(op_r_23__N_1226_adj_7377[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[19]), 
          .B1(op_r_23__N_1226_adj_7377[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31837), .COUT(n31838), .S0(op_r_23__N_1082_adj_7378[18]), 
          .S1(op_r_23__N_1082_adj_7378[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_18 (.A0(op_r_23__N_1268_adj_7375[16]), .B0(op_r_23__N_1226_adj_7377[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[17]), 
          .B1(op_r_23__N_1226_adj_7377[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31836), .COUT(n31837), .S0(op_r_23__N_1082_adj_7378[16]), 
          .S1(op_r_23__N_1082_adj_7378[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_16 (.A0(op_r_23__N_1268_adj_7375[14]), .B0(op_r_23__N_1226_adj_7377[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[15]), 
          .B1(op_r_23__N_1226_adj_7377[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31835), .COUT(n31836), .S0(op_r_23__N_1082_adj_7378[14]), 
          .S1(op_r_23__N_1082_adj_7378[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_14 (.A0(op_r_23__N_1268_adj_7375[12]), .B0(op_r_23__N_1226_adj_7377[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[13]), 
          .B1(op_r_23__N_1226_adj_7377[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31834), .COUT(n31835), .S0(op_r_23__N_1082_adj_7378[12]), 
          .S1(op_r_23__N_1082_adj_7378[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_12 (.A0(op_r_23__N_1268_adj_7375[10]), .B0(op_r_23__N_1226_adj_7377[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[11]), 
          .B1(op_r_23__N_1226_adj_7377[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31833), .COUT(n31834), .S0(op_r_23__N_1082_adj_7378[10]), 
          .S1(op_r_23__N_1082_adj_7378[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_10 (.A0(op_r_23__N_1268_adj_7375[8]), .B0(op_r_23__N_1226_adj_7377[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[9]), 
          .B1(op_r_23__N_1226_adj_7377[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31832), .COUT(n31833), .S0(op_r_23__N_1082_adj_7378[8]), 
          .S1(op_r_23__N_1082_adj_7378[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_8 (.A0(op_r_23__N_1268_adj_7375[6]), .B0(op_r_23__N_1226_adj_7377[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[7]), 
          .B1(op_r_23__N_1226_adj_7377[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31831), .COUT(n31832));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_6 (.A0(op_r_23__N_1268_adj_7375[4]), .B0(op_r_23__N_1226_adj_7377[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[5]), 
          .B1(op_r_23__N_1226_adj_7377[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31830), .COUT(n31831));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_4 (.A0(op_r_23__N_1268_adj_7375[2]), .B0(op_r_23__N_1226_adj_7377[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[3]), 
          .B1(op_r_23__N_1226_adj_7377[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31829), .COUT(n31830));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1042_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1042_add_4_2 (.A0(op_r_23__N_1268_adj_7375[0]), .B0(op_r_23__N_1226_adj_7377[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7375[1]), 
          .B1(op_r_23__N_1226_adj_7377[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n31829));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1042_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1042_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1042_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1042_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1125_add_4_12 (.A0(rom4_w_i[12]), .B0(s_count_adj_7402[0]), 
          .C0(s_count_adj_7402[2]), .D0(s_count_adj_7402[1]), .A1(rom4_w_i[12]), 
          .B1(s_count_adj_7402[0]), .C1(s_count_adj_7402[2]), .D1(s_count_adj_7402[1]), 
          .CIN(n31827), .S0(n12309), .S1(n119_adj_6625));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1125_add_4_12.INIT0 = 16'h9555;
    defparam _add_1_1125_add_4_12.INIT1 = 16'h9555;
    defparam _add_1_1125_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1125_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1125_add_4_10 (.A0(n34777), .B0(s_count_adj_7402[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(s_count_adj_7402[2]), .B1(n34776), .C1(rom4_w_i[12]), 
          .D1(VCC_net), .CIN(n31826), .COUT(n31827), .S0(n12307), .S1(n12308));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1125_add_4_10.INIT0 = 16'hddd2;
    defparam _add_1_1125_add_4_10.INIT1 = 16'h7877;
    defparam _add_1_1125_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1125_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1125_add_4_8 (.A0(n34777), .B0(s_count_adj_7402[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(n34777), .B1(s_count_adj_7402[0]), .C1(s_count_adj_7402[2]), 
          .D1(s_count_adj_7402[1]), .CIN(n31825), .COUT(n31826), .S0(n12305), 
          .S1(n12306));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1125_add_4_8.INIT0 = 16'hddd2;
    defparam _add_1_1125_add_4_8.INIT1 = 16'h9555;
    defparam _add_1_1125_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1125_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1125_add_4_6 (.A0(n34777), .B0(s_count_adj_7402[0]), .C0(s_count_adj_7402[2]), 
          .D0(s_count_adj_7402[1]), .A1(n34777), .B1(s_count_adj_7402[1]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31824), .COUT(n31825), .S0(n12303), 
          .S1(n12304));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1125_add_4_6.INIT0 = 16'h9555;
    defparam _add_1_1125_add_4_6.INIT1 = 16'hddd2;
    defparam _add_1_1125_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1125_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1125_add_4_4 (.A0(n34777), .B0(s_count_adj_7402[0]), .C0(s_count_adj_7402[2]), 
          .D0(s_count_adj_7402[1]), .A1(n34777), .B1(s_count_adj_7402[1]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n31823), .COUT(n31824), .S0(n12301), 
          .S1(n12302));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1125_add_4_4.INIT0 = 16'h9555;
    defparam _add_1_1125_add_4_4.INIT1 = 16'hddd2;
    defparam _add_1_1125_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1125_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1125_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(s_count_adj_7402[2]), .B1(s_count_adj_7402[0]), 
          .C1(n34777), .D1(VCC_net), .COUT(n31823), .S1(n12300));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1125_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1125_add_4_2.INIT1 = 16'h8788;
    defparam _add_1_1125_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1125_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_32 (.A0(op_r_23__N_1268_adj_7324[30]), .B0(op_i_23__N_1310_adj_7329[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[31]), 
          .B1(op_i_23__N_1310_adj_7329[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31821), .S0(op_i_23__N_1130_adj_7330[30]), .S1(op_i_23__N_1130_adj_7330[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_30 (.A0(op_r_23__N_1268_adj_7324[28]), .B0(op_i_23__N_1310_adj_7329[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[29]), 
          .B1(op_i_23__N_1310_adj_7329[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31820), .COUT(n31821), .S0(op_i_23__N_1130_adj_7330[28]), 
          .S1(op_i_23__N_1130_adj_7330[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_28 (.A0(op_r_23__N_1268_adj_7324[26]), .B0(op_i_23__N_1310_adj_7329[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[27]), 
          .B1(op_i_23__N_1310_adj_7329[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31819), .COUT(n31820), .S0(op_i_23__N_1130_adj_7330[26]), 
          .S1(op_i_23__N_1130_adj_7330[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_26 (.A0(op_r_23__N_1268_adj_7324[24]), .B0(op_i_23__N_1310_adj_7329[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[25]), 
          .B1(op_i_23__N_1310_adj_7329[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31818), .COUT(n31819), .S0(op_i_23__N_1130_adj_7330[24]), 
          .S1(op_i_23__N_1130_adj_7330[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_24 (.A0(op_r_23__N_1268_adj_7324[22]), .B0(op_i_23__N_1310_adj_7329[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[23]), 
          .B1(op_i_23__N_1310_adj_7329[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31817), .COUT(n31818), .S0(op_i_23__N_1130_adj_7330[22]), 
          .S1(op_i_23__N_1130_adj_7330[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_22 (.A0(op_r_23__N_1268_adj_7324[20]), .B0(op_i_23__N_1310_adj_7329[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[21]), 
          .B1(op_i_23__N_1310_adj_7329[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31816), .COUT(n31817), .S0(op_i_23__N_1130_adj_7330[20]), 
          .S1(op_i_23__N_1130_adj_7330[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_20 (.A0(op_r_23__N_1268_adj_7324[18]), .B0(op_i_23__N_1310_adj_7329[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[19]), 
          .B1(op_i_23__N_1310_adj_7329[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31815), .COUT(n31816), .S0(op_i_23__N_1130_adj_7330[18]), 
          .S1(op_i_23__N_1130_adj_7330[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_18 (.A0(op_r_23__N_1268_adj_7324[16]), .B0(op_i_23__N_1310_adj_7329[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[17]), 
          .B1(op_i_23__N_1310_adj_7329[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31814), .COUT(n31815), .S0(op_i_23__N_1130_adj_7330[16]), 
          .S1(op_i_23__N_1130_adj_7330[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_16 (.A0(op_r_23__N_1268_adj_7324[14]), .B0(op_i_23__N_1310_adj_7329[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[15]), 
          .B1(op_i_23__N_1310_adj_7329[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31813), .COUT(n31814), .S0(op_i_23__N_1130_adj_7330[14]), 
          .S1(op_i_23__N_1130_adj_7330[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_14 (.A0(op_r_23__N_1268_adj_7324[12]), .B0(op_i_23__N_1310_adj_7329[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[13]), 
          .B1(op_i_23__N_1310_adj_7329[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31812), .COUT(n31813), .S0(op_i_23__N_1130_adj_7330[12]), 
          .S1(op_i_23__N_1130_adj_7330[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_12 (.A0(op_r_23__N_1268_adj_7324[10]), .B0(op_i_23__N_1310_adj_7329[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[11]), 
          .B1(op_i_23__N_1310_adj_7329[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31811), .COUT(n31812), .S0(op_i_23__N_1130_adj_7330[10]), 
          .S1(op_i_23__N_1130_adj_7330[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_10 (.A0(op_r_23__N_1268_adj_7324[8]), .B0(op_i_23__N_1310_adj_7329[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[9]), 
          .B1(op_i_23__N_1310_adj_7329[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31810), .COUT(n31811), .S0(op_i_23__N_1130_adj_7330[8]), 
          .S1(op_i_23__N_1130_adj_7330[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_8 (.A0(op_r_23__N_1268_adj_7324[6]), .B0(op_i_23__N_1310_adj_7329[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[7]), 
          .B1(op_i_23__N_1310_adj_7329[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31809), .COUT(n31810));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_8.INJECT1_1 = "NO";
    PFUMX i15764 (.BLUT(n34139), .ALUT(n34140), .C0(y_1_delay[1]), .Z(n34148));
    CCU2C _add_1_1131_add_4_5 (.A0(n34735), .B0(n34730), .C0(count[5]), 
          .D0(n20095), .A1(n30197), .B1(n34729), .C1(count[5]), .D1(n20103), 
          .CIN(n31802), .COUT(n31803), .S0(n12347), .S1(n12348));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1131_add_4_5.INIT0 = 16'h8878;
    defparam _add_1_1131_add_4_5.INIT1 = 16'h8878;
    defparam _add_1_1131_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1131_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1012_add_4_4 (.A0(op_r_23__N_1268_adj_7324[2]), .B0(op_i_23__N_1310_adj_7329[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[3]), 
          .B1(op_i_23__N_1310_adj_7329[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31807), .COUT(n31808));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1131_add_4_11 (.A0(n34713), .B0(n34759), .C0(n34789), 
          .D0(count[5]), .A1(n34713), .B1(n34759), .C1(n34789), .D1(count[5]), 
          .CIN(n31805), .S0(n12353), .S1(n12368));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1131_add_4_11.INIT0 = 16'ha6aa;
    defparam _add_1_1131_add_4_11.INIT1 = 16'ha6aa;
    defparam _add_1_1131_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1131_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1131_add_4_7 (.A0(n30203), .B0(n34737), .C0(count[5]), 
          .D0(n28591), .A1(n34736), .B1(n33051), .C1(count[5]), .D1(n34733), 
          .CIN(n31803), .COUT(n31804), .S0(n12349), .S1(n12350));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1131_add_4_7.INIT0 = 16'h8878;
    defparam _add_1_1131_add_4_7.INIT1 = 16'h8878;
    defparam _add_1_1131_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1131_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1131_add_4_3 (.A0(n30499), .B0(n33030), .C0(count[5]), 
          .D0(n20089), .A1(n30207), .B1(n34730), .C1(count[5]), .D1(n28589), 
          .CIN(n31801), .COUT(n31802), .S0(n12345), .S1(n12346));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1131_add_4_3.INIT0 = 16'h8878;
    defparam _add_1_1131_add_4_3.INIT1 = 16'h8878;
    defparam _add_1_1131_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1131_add_4_3.INJECT1_1 = "NO";
    LUT4 i15193_3_lut (.A(\result_i[20] [7]), .B(\result_i[21] [7]), .C(y_1_delay[0]), 
         .Z(n33577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15193_3_lut.init = 16'hcaca;
    CCU2C _add_1_1012_add_4_6 (.A0(op_r_23__N_1268_adj_7324[4]), .B0(op_i_23__N_1310_adj_7329[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[5]), 
          .B1(op_i_23__N_1310_adj_7329[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31808), .COUT(n31809));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1012_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1012_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1012_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1012_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1131_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n34727), .B1(n34757), .C1(count[4]), .D1(count[5]), 
          .COUT(n31801), .S1(n12344));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[17:28])
    defparam _add_1_1131_add_4_1.INIT0 = 16'h000F;
    defparam _add_1_1131_add_4_1.INIT1 = 16'ha9aa;
    defparam _add_1_1131_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1131_add_4_1.INJECT1_1 = "NO";
    LUT4 i7761_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[363])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7761_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7753_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[364])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7753_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7745_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[365])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7745_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7737_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[366])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7737_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7729_3_lut_4_lut (.A(n34717), .B(n34706), .C(\result_r[9] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[367])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7729_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15537_3_lut (.A(\result_r[26] [11]), .B(\result_r[27] [11]), .C(y_1_delay[0]), 
         .Z(n33921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15537_3_lut.init = 16'hcaca;
    PFUMX i15509 (.BLUT(n33877), .ALUT(n33878), .C0(y_1_delay[1]), .Z(n33893));
    LUT4 i3889_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[336])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3889_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15536_3_lut (.A(\result_r[24] [11]), .B(\result_r[25] [11]), .C(y_1_delay[0]), 
         .Z(n33920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15536_3_lut.init = 16'hcaca;
    LUT4 i3881_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[337])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3881_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15285_3_lut (.A(\result_i[18] [4]), .B(\result_i[19] [4]), .C(y_1_delay[0]), 
         .Z(n33669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15285_3_lut.init = 16'hcaca;
    LUT4 i3873_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[338])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3873_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3865_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[339])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3865_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15192_3_lut (.A(\result_i[18] [7]), .B(\result_i[19] [7]), .C(y_1_delay[0]), 
         .Z(n33576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15192_3_lut.init = 16'hcaca;
    LUT4 i3857_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[340])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3857_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3849_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[341])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3849_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15510 (.BLUT(n33879), .ALUT(n33880), .C0(y_1_delay[1]), .Z(n33894));
    LUT4 i3841_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[342])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3841_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15191_3_lut (.A(\result_i[16] [7]), .B(\result_i[17] [7]), .C(y_1_delay[0]), 
         .Z(n33575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15191_3_lut.init = 16'hcaca;
    LUT4 i3833_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[343])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3833_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15511 (.BLUT(n33881), .ALUT(n33882), .C0(y_1_delay[1]), .Z(n33895));
    LUT4 i15284_3_lut (.A(\result_i[16] [4]), .B(\result_i[17] [4]), .C(y_1_delay[0]), 
         .Z(n33668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15284_3_lut.init = 16'hcaca;
    LUT4 i3825_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[344])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3825_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3817_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[345])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3817_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15535_3_lut (.A(\result_r[22] [11]), .B(\result_r[23] [11]), .C(y_1_delay[0]), 
         .Z(n33919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15535_3_lut.init = 16'hcaca;
    LUT4 i15716_3_lut (.A(\result_r[12] [5]), .B(\result_r[13] [5]), .C(y_1_delay[0]), 
         .Z(n34100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15716_3_lut.init = 16'hcaca;
    LUT4 i14940_3_lut (.A(\result_i[10] [15]), .B(\result_i[11] [15]), .C(y_1_delay[0]), 
         .Z(n33324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14940_3_lut.init = 16'hcaca;
    LUT4 i14939_3_lut (.A(\result_i[8] [15]), .B(\result_i[9] [15]), .C(y_1_delay[0]), 
         .Z(n33323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14939_3_lut.init = 16'hcaca;
    LUT4 i15715_3_lut (.A(\result_r[10] [5]), .B(\result_r[11] [5]), .C(y_1_delay[0]), 
         .Z(n34099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15715_3_lut.init = 16'hcaca;
    LUT4 i15714_3_lut (.A(\result_r[8] [5]), .B(\result_r[9] [5]), .C(y_1_delay[0]), 
         .Z(n34098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15714_3_lut.init = 16'hcaca;
    LUT4 i15713_3_lut (.A(\result_r[6] [5]), .B(\result_r[7] [5]), .C(y_1_delay[0]), 
         .Z(n34097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15713_3_lut.init = 16'hcaca;
    LUT4 i15712_3_lut (.A(\result_r[4] [5]), .B(\result_r[5] [5]), .C(y_1_delay[0]), 
         .Z(n34096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15712_3_lut.init = 16'hcaca;
    LUT4 i14919_3_lut (.A(\result_r[30] [0]), .B(\result_r[31] [0]), .C(y_1_delay[0]), 
         .Z(n33303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14919_3_lut.init = 16'hcaca;
    LUT4 i14918_3_lut (.A(\result_r[28] [0]), .B(\result_r[29] [0]), .C(y_1_delay[0]), 
         .Z(n33302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14918_3_lut.init = 16'hcaca;
    LUT4 i15711_3_lut (.A(\result_r[2] [5]), .B(\result_r[3] [5]), .C(y_1_delay[0]), 
         .Z(n34095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15711_3_lut.init = 16'hcaca;
    LUT4 i15710_3_lut (.A(\result_r[0] [5]), .B(\result_r[1] [5]), .C(y_1_delay[0]), 
         .Z(n34094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15710_3_lut.init = 16'hcaca;
    LUT4 i14917_3_lut (.A(\result_r[26] [0]), .B(\result_r[27] [0]), .C(y_1_delay[0]), 
         .Z(n33301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14917_3_lut.init = 16'hcaca;
    LUT4 i14916_3_lut (.A(\result_r[24] [0]), .B(\result_r[25] [0]), .C(y_1_delay[0]), 
         .Z(n33300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14916_3_lut.init = 16'hcaca;
    LUT4 i14915_3_lut (.A(\result_r[22] [0]), .B(\result_r[23] [0]), .C(y_1_delay[0]), 
         .Z(n33299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14915_3_lut.init = 16'hcaca;
    LUT4 i14914_3_lut (.A(\result_r[20] [0]), .B(\result_r[21] [0]), .C(y_1_delay[0]), 
         .Z(n33298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14914_3_lut.init = 16'hcaca;
    LUT4 i14981_3_lut (.A(\result_i[30] [14]), .B(\result_i[31] [14]), .C(y_1_delay[0]), 
         .Z(n33365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14981_3_lut.init = 16'hcaca;
    LUT4 i14980_3_lut (.A(\result_i[28] [14]), .B(\result_i[29] [14]), .C(y_1_delay[0]), 
         .Z(n33364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14980_3_lut.init = 16'hcaca;
    LUT4 i14979_3_lut (.A(\result_i[26] [14]), .B(\result_i[27] [14]), .C(y_1_delay[0]), 
         .Z(n33363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14979_3_lut.init = 16'hcaca;
    LUT4 i14978_3_lut (.A(\result_i[24] [14]), .B(\result_i[25] [14]), .C(y_1_delay[0]), 
         .Z(n33362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14978_3_lut.init = 16'hcaca;
    LUT4 i14913_3_lut (.A(\result_r[18] [0]), .B(\result_r[19] [0]), .C(y_1_delay[0]), 
         .Z(n33297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14913_3_lut.init = 16'hcaca;
    LUT4 i14912_3_lut (.A(\result_r[16] [0]), .B(\result_r[17] [0]), .C(y_1_delay[0]), 
         .Z(n33296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14912_3_lut.init = 16'hcaca;
    LUT4 i14977_3_lut (.A(\result_i[22] [14]), .B(\result_i[23] [14]), .C(y_1_delay[0]), 
         .Z(n33361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14977_3_lut.init = 16'hcaca;
    LUT4 i14976_3_lut (.A(\result_i[20] [14]), .B(\result_i[21] [14]), .C(y_1_delay[0]), 
         .Z(n33360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14976_3_lut.init = 16'hcaca;
    LUT4 i14911_3_lut (.A(\result_r[14] [0]), .B(\result_r[15] [0]), .C(y_1_delay[0]), 
         .Z(n33295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14911_3_lut.init = 16'hcaca;
    LUT4 i14910_3_lut (.A(\result_r[12] [0]), .B(\result_r[13] [0]), .C(y_1_delay[0]), 
         .Z(n33294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14910_3_lut.init = 16'hcaca;
    LUT4 i14909_3_lut (.A(\result_r[10] [0]), .B(\result_r[11] [0]), .C(y_1_delay[0]), 
         .Z(n33293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14909_3_lut.init = 16'hcaca;
    LUT4 i14908_3_lut (.A(\result_r[8] [0]), .B(\result_r[9] [0]), .C(y_1_delay[0]), 
         .Z(n33292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14908_3_lut.init = 16'hcaca;
    LUT4 i14907_3_lut (.A(\result_r[6] [0]), .B(\result_r[7] [0]), .C(y_1_delay[0]), 
         .Z(n33291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14907_3_lut.init = 16'hcaca;
    LUT4 i14906_3_lut (.A(\result_r[4] [0]), .B(\result_r[5] [0]), .C(y_1_delay[0]), 
         .Z(n33290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14906_3_lut.init = 16'hcaca;
    LUT4 i14975_3_lut (.A(\result_i[18] [14]), .B(\result_i[19] [14]), .C(y_1_delay[0]), 
         .Z(n33359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14975_3_lut.init = 16'hcaca;
    LUT4 i14974_3_lut (.A(\result_i[16] [14]), .B(\result_i[17] [14]), .C(y_1_delay[0]), 
         .Z(n33358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14974_3_lut.init = 16'hcaca;
    LUT4 i14905_3_lut (.A(\result_r[2] [0]), .B(\result_r[3] [0]), .C(y_1_delay[0]), 
         .Z(n33289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14905_3_lut.init = 16'hcaca;
    LUT4 i14904_3_lut (.A(\result_r[0] [0]), .B(\result_r[1] [0]), .C(y_1_delay[0]), 
         .Z(n33288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14904_3_lut.init = 16'hcaca;
    LUT4 i14973_3_lut (.A(\result_i[14] [14]), .B(\result_i[15] [14]), .C(y_1_delay[0]), 
         .Z(n33357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14973_3_lut.init = 16'hcaca;
    LUT4 i14972_3_lut (.A(\result_i[12] [14]), .B(\result_i[13] [14]), .C(y_1_delay[0]), 
         .Z(n33356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14972_3_lut.init = 16'hcaca;
    LUT4 i14971_3_lut (.A(\result_i[10] [14]), .B(\result_i[11] [14]), .C(y_1_delay[0]), 
         .Z(n33355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14971_3_lut.init = 16'hcaca;
    LUT4 i14970_3_lut (.A(\result_i[8] [14]), .B(\result_i[9] [14]), .C(y_1_delay[0]), 
         .Z(n33354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14970_3_lut.init = 16'hcaca;
    LUT4 i14969_3_lut (.A(\result_i[6] [14]), .B(\result_i[7] [14]), .C(y_1_delay[0]), 
         .Z(n33353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14969_3_lut.init = 16'hcaca;
    LUT4 i14968_3_lut (.A(\result_i[4] [14]), .B(\result_i[5] [14]), .C(y_1_delay[0]), 
         .Z(n33352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14968_3_lut.init = 16'hcaca;
    LUT4 i14967_3_lut (.A(\result_i[2] [14]), .B(\result_i[3] [14]), .C(y_1_delay[0]), 
         .Z(n33351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14967_3_lut.init = 16'hcaca;
    LUT4 i14966_3_lut (.A(\result_i[0] [14]), .B(\result_i[1] [14]), .C(y_1_delay[0]), 
         .Z(n33350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14966_3_lut.init = 16'hcaca;
    LUT4 i14938_3_lut (.A(\result_i[6] [15]), .B(\result_i[7] [15]), .C(y_1_delay[0]), 
         .Z(n33322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14938_3_lut.init = 16'hcaca;
    LUT4 i14937_3_lut (.A(\result_i[4] [15]), .B(\result_i[5] [15]), .C(y_1_delay[0]), 
         .Z(n33321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14937_3_lut.init = 16'hcaca;
    LUT4 i15384_3_lut (.A(\result_i[30] [1]), .B(\result_i[31] [1]), .C(y_1_delay[0]), 
         .Z(n33768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15384_3_lut.init = 16'hcaca;
    LUT4 i15383_3_lut (.A(\result_i[28] [1]), .B(\result_i[29] [1]), .C(y_1_delay[0]), 
         .Z(n33767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15383_3_lut.init = 16'hcaca;
    LUT4 i15382_3_lut (.A(\result_i[26] [1]), .B(\result_i[27] [1]), .C(y_1_delay[0]), 
         .Z(n33766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15382_3_lut.init = 16'hcaca;
    LUT4 i15381_3_lut (.A(\result_i[24] [1]), .B(\result_i[25] [1]), .C(y_1_delay[0]), 
         .Z(n33765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15381_3_lut.init = 16'hcaca;
    LUT4 i15380_3_lut (.A(\result_i[22] [1]), .B(\result_i[23] [1]), .C(y_1_delay[0]), 
         .Z(n33764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15380_3_lut.init = 16'hcaca;
    LUT4 i15379_3_lut (.A(\result_i[20] [1]), .B(\result_i[21] [1]), .C(y_1_delay[0]), 
         .Z(n33763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15379_3_lut.init = 16'hcaca;
    LUT4 i15378_3_lut (.A(\result_i[18] [1]), .B(\result_i[19] [1]), .C(y_1_delay[0]), 
         .Z(n33762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15378_3_lut.init = 16'hcaca;
    LUT4 i15377_3_lut (.A(\result_i[16] [1]), .B(\result_i[17] [1]), .C(y_1_delay[0]), 
         .Z(n33761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15377_3_lut.init = 16'hcaca;
    LUT4 i15376_3_lut (.A(\result_i[14] [1]), .B(\result_i[15] [1]), .C(y_1_delay[0]), 
         .Z(n33760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15376_3_lut.init = 16'hcaca;
    LUT4 i15375_3_lut (.A(\result_i[12] [1]), .B(\result_i[13] [1]), .C(y_1_delay[0]), 
         .Z(n33759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15375_3_lut.init = 16'hcaca;
    LUT4 i15374_3_lut (.A(\result_i[10] [1]), .B(\result_i[11] [1]), .C(y_1_delay[0]), 
         .Z(n33758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15374_3_lut.init = 16'hcaca;
    LUT4 i15373_3_lut (.A(\result_i[8] [1]), .B(\result_i[9] [1]), .C(y_1_delay[0]), 
         .Z(n33757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15373_3_lut.init = 16'hcaca;
    LUT4 i15372_3_lut (.A(\result_i[6] [1]), .B(\result_i[7] [1]), .C(y_1_delay[0]), 
         .Z(n33756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15372_3_lut.init = 16'hcaca;
    LUT4 i15371_3_lut (.A(\result_i[4] [1]), .B(\result_i[5] [1]), .C(y_1_delay[0]), 
         .Z(n33755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15371_3_lut.init = 16'hcaca;
    LUT4 i15370_3_lut (.A(\result_i[2] [1]), .B(\result_i[3] [1]), .C(y_1_delay[0]), 
         .Z(n33754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15370_3_lut.init = 16'hcaca;
    LUT4 i15369_3_lut (.A(\result_i[0] [1]), .B(\result_i[1] [1]), .C(y_1_delay[0]), 
         .Z(n33753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15369_3_lut.init = 16'hcaca;
    LUT4 i14888_3_lut (.A(\result_i[30] [0]), .B(\result_i[31] [0]), .C(y_1_delay[0]), 
         .Z(n33272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14888_3_lut.init = 16'hcaca;
    LUT4 i14887_3_lut (.A(\result_i[28] [0]), .B(\result_i[29] [0]), .C(y_1_delay[0]), 
         .Z(n33271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14887_3_lut.init = 16'hcaca;
    LUT4 i14886_3_lut (.A(\result_i[26] [0]), .B(\result_i[27] [0]), .C(y_1_delay[0]), 
         .Z(n33270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14886_3_lut.init = 16'hcaca;
    LUT4 i14885_3_lut (.A(\result_i[24] [0]), .B(\result_i[25] [0]), .C(y_1_delay[0]), 
         .Z(n33269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14885_3_lut.init = 16'hcaca;
    LUT4 i14884_3_lut (.A(\result_i[22] [0]), .B(\result_i[23] [0]), .C(y_1_delay[0]), 
         .Z(n33268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14884_3_lut.init = 16'hcaca;
    LUT4 i14883_3_lut (.A(\result_i[20] [0]), .B(\result_i[21] [0]), .C(y_1_delay[0]), 
         .Z(n33267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14883_3_lut.init = 16'hcaca;
    LUT4 i14882_3_lut (.A(\result_i[18] [0]), .B(\result_i[19] [0]), .C(y_1_delay[0]), 
         .Z(n33266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14882_3_lut.init = 16'hcaca;
    LUT4 i14881_3_lut (.A(\result_i[16] [0]), .B(\result_i[17] [0]), .C(y_1_delay[0]), 
         .Z(n33265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14881_3_lut.init = 16'hcaca;
    LUT4 i14880_3_lut (.A(\result_i[14] [0]), .B(\result_i[15] [0]), .C(y_1_delay[0]), 
         .Z(n33264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14880_3_lut.init = 16'hcaca;
    LUT4 i14879_3_lut (.A(\result_i[12] [0]), .B(\result_i[13] [0]), .C(y_1_delay[0]), 
         .Z(n33263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14879_3_lut.init = 16'hcaca;
    LUT4 i14878_3_lut (.A(\result_i[10] [0]), .B(\result_i[11] [0]), .C(y_1_delay[0]), 
         .Z(n33262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14878_3_lut.init = 16'hcaca;
    LUT4 i14877_3_lut (.A(\result_i[8] [0]), .B(\result_i[9] [0]), .C(y_1_delay[0]), 
         .Z(n33261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14877_3_lut.init = 16'hcaca;
    LUT4 i14876_3_lut (.A(\result_i[6] [0]), .B(\result_i[7] [0]), .C(y_1_delay[0]), 
         .Z(n33260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14876_3_lut.init = 16'hcaca;
    LUT4 i14875_3_lut (.A(\result_i[4] [0]), .B(\result_i[5] [0]), .C(y_1_delay[0]), 
         .Z(n33259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14875_3_lut.init = 16'hcaca;
    LUT4 i14874_3_lut (.A(\result_i[2] [0]), .B(\result_i[3] [0]), .C(y_1_delay[0]), 
         .Z(n33258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14874_3_lut.init = 16'hcaca;
    LUT4 i14873_3_lut (.A(\result_i[0] [0]), .B(\result_i[1] [0]), .C(y_1_delay[0]), 
         .Z(n33257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14873_3_lut.init = 16'hcaca;
    LUT4 i15694_3_lut (.A(\result_r[30] [6]), .B(\result_r[31] [6]), .C(y_1_delay[0]), 
         .Z(n34078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15694_3_lut.init = 16'hcaca;
    LUT4 i15693_3_lut (.A(\result_r[28] [6]), .B(\result_r[29] [6]), .C(y_1_delay[0]), 
         .Z(n34077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15693_3_lut.init = 16'hcaca;
    LUT4 i15692_3_lut (.A(\result_r[26] [6]), .B(\result_r[27] [6]), .C(y_1_delay[0]), 
         .Z(n34076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15692_3_lut.init = 16'hcaca;
    LUT4 i15691_3_lut (.A(\result_r[24] [6]), .B(\result_r[25] [6]), .C(y_1_delay[0]), 
         .Z(n34075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15691_3_lut.init = 16'hcaca;
    LUT4 i15690_3_lut (.A(\result_r[22] [6]), .B(\result_r[23] [6]), .C(y_1_delay[0]), 
         .Z(n34074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15690_3_lut.init = 16'hcaca;
    LUT4 i15689_3_lut (.A(\result_r[20] [6]), .B(\result_r[21] [6]), .C(y_1_delay[0]), 
         .Z(n34073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15689_3_lut.init = 16'hcaca;
    LUT4 i15353_3_lut (.A(\result_i[30] [2]), .B(\result_i[31] [2]), .C(y_1_delay[0]), 
         .Z(n33737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15353_3_lut.init = 16'hcaca;
    LUT4 i15352_3_lut (.A(\result_i[28] [2]), .B(\result_i[29] [2]), .C(y_1_delay[0]), 
         .Z(n33736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15352_3_lut.init = 16'hcaca;
    LUT4 i15351_3_lut (.A(\result_i[26] [2]), .B(\result_i[27] [2]), .C(y_1_delay[0]), 
         .Z(n33735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15351_3_lut.init = 16'hcaca;
    LUT4 i15350_3_lut (.A(\result_i[24] [2]), .B(\result_i[25] [2]), .C(y_1_delay[0]), 
         .Z(n33734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15350_3_lut.init = 16'hcaca;
    LUT4 i15349_3_lut (.A(\result_i[22] [2]), .B(\result_i[23] [2]), .C(y_1_delay[0]), 
         .Z(n33733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15349_3_lut.init = 16'hcaca;
    LUT4 i15348_3_lut (.A(\result_i[20] [2]), .B(\result_i[21] [2]), .C(y_1_delay[0]), 
         .Z(n33732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15348_3_lut.init = 16'hcaca;
    LUT4 i15347_3_lut (.A(\result_i[18] [2]), .B(\result_i[19] [2]), .C(y_1_delay[0]), 
         .Z(n33731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15347_3_lut.init = 16'hcaca;
    LUT4 i15346_3_lut (.A(\result_i[16] [2]), .B(\result_i[17] [2]), .C(y_1_delay[0]), 
         .Z(n33730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15346_3_lut.init = 16'hcaca;
    LUT4 i15345_3_lut (.A(\result_i[14] [2]), .B(\result_i[15] [2]), .C(y_1_delay[0]), 
         .Z(n33729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15345_3_lut.init = 16'hcaca;
    LUT4 i15344_3_lut (.A(\result_i[12] [2]), .B(\result_i[13] [2]), .C(y_1_delay[0]), 
         .Z(n33728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15344_3_lut.init = 16'hcaca;
    LUT4 i15343_3_lut (.A(\result_i[10] [2]), .B(\result_i[11] [2]), .C(y_1_delay[0]), 
         .Z(n33727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15343_3_lut.init = 16'hcaca;
    LUT4 i15342_3_lut (.A(\result_i[8] [2]), .B(\result_i[9] [2]), .C(y_1_delay[0]), 
         .Z(n33726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15342_3_lut.init = 16'hcaca;
    LUT4 i15341_3_lut (.A(\result_i[6] [2]), .B(\result_i[7] [2]), .C(y_1_delay[0]), 
         .Z(n33725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15341_3_lut.init = 16'hcaca;
    LUT4 i15340_3_lut (.A(\result_i[4] [2]), .B(\result_i[5] [2]), .C(y_1_delay[0]), 
         .Z(n33724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15340_3_lut.init = 16'hcaca;
    LUT4 i15339_3_lut (.A(\result_i[2] [2]), .B(\result_i[3] [2]), .C(y_1_delay[0]), 
         .Z(n33723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15339_3_lut.init = 16'hcaca;
    LUT4 i15338_3_lut (.A(\result_i[0] [2]), .B(\result_i[1] [2]), .C(y_1_delay[0]), 
         .Z(n33722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15338_3_lut.init = 16'hcaca;
    LUT4 i15322_3_lut (.A(\result_i[30] [3]), .B(\result_i[31] [3]), .C(y_1_delay[0]), 
         .Z(n33706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15322_3_lut.init = 16'hcaca;
    LUT4 i15321_3_lut (.A(\result_i[28] [3]), .B(\result_i[29] [3]), .C(y_1_delay[0]), 
         .Z(n33705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15321_3_lut.init = 16'hcaca;
    LUT4 i15320_3_lut (.A(\result_i[26] [3]), .B(\result_i[27] [3]), .C(y_1_delay[0]), 
         .Z(n33704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15320_3_lut.init = 16'hcaca;
    LUT4 i15319_3_lut (.A(\result_i[24] [3]), .B(\result_i[25] [3]), .C(y_1_delay[0]), 
         .Z(n33703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15319_3_lut.init = 16'hcaca;
    LUT4 i15318_3_lut (.A(\result_i[22] [3]), .B(\result_i[23] [3]), .C(y_1_delay[0]), 
         .Z(n33702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15318_3_lut.init = 16'hcaca;
    LUT4 i15317_3_lut (.A(\result_i[20] [3]), .B(\result_i[21] [3]), .C(y_1_delay[0]), 
         .Z(n33701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15317_3_lut.init = 16'hcaca;
    LUT4 i15316_3_lut (.A(\result_i[18] [3]), .B(\result_i[19] [3]), .C(y_1_delay[0]), 
         .Z(n33700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15316_3_lut.init = 16'hcaca;
    LUT4 i15315_3_lut (.A(\result_i[16] [3]), .B(\result_i[17] [3]), .C(y_1_delay[0]), 
         .Z(n33699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15315_3_lut.init = 16'hcaca;
    LUT4 i15314_3_lut (.A(\result_i[14] [3]), .B(\result_i[15] [3]), .C(y_1_delay[0]), 
         .Z(n33698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15314_3_lut.init = 16'hcaca;
    LUT4 i15313_3_lut (.A(\result_i[12] [3]), .B(\result_i[13] [3]), .C(y_1_delay[0]), 
         .Z(n33697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15313_3_lut.init = 16'hcaca;
    LUT4 i15688_3_lut (.A(\result_r[18] [6]), .B(\result_r[19] [6]), .C(y_1_delay[0]), 
         .Z(n34072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15688_3_lut.init = 16'hcaca;
    LUT4 i15687_3_lut (.A(\result_r[16] [6]), .B(\result_r[17] [6]), .C(y_1_delay[0]), 
         .Z(n34071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15687_3_lut.init = 16'hcaca;
    LUT4 i15074_3_lut (.A(\result_i[30] [11]), .B(\result_i[31] [11]), .C(y_1_delay[0]), 
         .Z(n33458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15074_3_lut.init = 16'hcaca;
    LUT4 i15073_3_lut (.A(\result_i[28] [11]), .B(\result_i[29] [11]), .C(y_1_delay[0]), 
         .Z(n33457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15073_3_lut.init = 16'hcaca;
    LUT4 i15312_3_lut (.A(\result_i[10] [3]), .B(\result_i[11] [3]), .C(y_1_delay[0]), 
         .Z(n33696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15312_3_lut.init = 16'hcaca;
    LUT4 i15311_3_lut (.A(\result_i[8] [3]), .B(\result_i[9] [3]), .C(y_1_delay[0]), 
         .Z(n33695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15311_3_lut.init = 16'hcaca;
    LUT4 i15072_3_lut (.A(\result_i[26] [11]), .B(\result_i[27] [11]), .C(y_1_delay[0]), 
         .Z(n33456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15072_3_lut.init = 16'hcaca;
    LUT4 i15071_3_lut (.A(\result_i[24] [11]), .B(\result_i[25] [11]), .C(y_1_delay[0]), 
         .Z(n33455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15071_3_lut.init = 16'hcaca;
    LUT4 i15310_3_lut (.A(\result_i[6] [3]), .B(\result_i[7] [3]), .C(y_1_delay[0]), 
         .Z(n33694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15310_3_lut.init = 16'hcaca;
    LUT4 i15093_3_lut (.A(\result_i[6] [10]), .B(\result_i[7] [10]), .C(y_1_delay[0]), 
         .Z(n33477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15093_3_lut.init = 16'hcaca;
    LUT4 i14947_3_lut (.A(\result_i[24] [15]), .B(\result_i[25] [15]), .C(y_1_delay[0]), 
         .Z(n33331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14947_3_lut.init = 16'hcaca;
    LUT4 i15309_3_lut (.A(\result_i[4] [3]), .B(\result_i[5] [3]), .C(y_1_delay[0]), 
         .Z(n33693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15309_3_lut.init = 16'hcaca;
    LUT4 i15070_3_lut (.A(\result_i[22] [11]), .B(\result_i[23] [11]), .C(y_1_delay[0]), 
         .Z(n33454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15070_3_lut.init = 16'hcaca;
    LUT4 i15069_3_lut (.A(\result_i[20] [11]), .B(\result_i[21] [11]), .C(y_1_delay[0]), 
         .Z(n33453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15069_3_lut.init = 16'hcaca;
    LUT4 i15686_3_lut (.A(\result_r[14] [6]), .B(\result_r[15] [6]), .C(y_1_delay[0]), 
         .Z(n34070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15686_3_lut.init = 16'hcaca;
    LUT4 i15685_3_lut (.A(\result_r[12] [6]), .B(\result_r[13] [6]), .C(y_1_delay[0]), 
         .Z(n34069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15685_3_lut.init = 16'hcaca;
    LUT4 i15068_3_lut (.A(\result_i[18] [11]), .B(\result_i[19] [11]), .C(y_1_delay[0]), 
         .Z(n33452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15068_3_lut.init = 16'hcaca;
    LUT4 i15067_3_lut (.A(\result_i[16] [11]), .B(\result_i[17] [11]), .C(y_1_delay[0]), 
         .Z(n33451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15067_3_lut.init = 16'hcaca;
    LUT4 i15684_3_lut (.A(\result_r[10] [6]), .B(\result_r[11] [6]), .C(y_1_delay[0]), 
         .Z(n34068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15684_3_lut.init = 16'hcaca;
    LUT4 i15683_3_lut (.A(\result_r[8] [6]), .B(\result_r[9] [6]), .C(y_1_delay[0]), 
         .Z(n34067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15683_3_lut.init = 16'hcaca;
    LUT4 i15308_3_lut (.A(\result_i[2] [3]), .B(\result_i[3] [3]), .C(y_1_delay[0]), 
         .Z(n33692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15308_3_lut.init = 16'hcaca;
    LUT4 i15092_3_lut (.A(\result_i[4] [10]), .B(\result_i[5] [10]), .C(y_1_delay[0]), 
         .Z(n33476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15092_3_lut.init = 16'hcaca;
    LUT4 i15307_3_lut (.A(\result_i[0] [3]), .B(\result_i[1] [3]), .C(y_1_delay[0]), 
         .Z(n33691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15307_3_lut.init = 16'hcaca;
    LUT4 i15066_3_lut (.A(\result_i[14] [11]), .B(\result_i[15] [11]), .C(y_1_delay[0]), 
         .Z(n33450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15066_3_lut.init = 16'hcaca;
    LUT4 i15065_3_lut (.A(\result_i[12] [11]), .B(\result_i[13] [11]), .C(y_1_delay[0]), 
         .Z(n33449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15065_3_lut.init = 16'hcaca;
    LUT4 i15064_3_lut (.A(\result_i[10] [11]), .B(\result_i[11] [11]), .C(y_1_delay[0]), 
         .Z(n33448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15064_3_lut.init = 16'hcaca;
    LUT4 i15063_3_lut (.A(\result_i[8] [11]), .B(\result_i[9] [11]), .C(y_1_delay[0]), 
         .Z(n33447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15063_3_lut.init = 16'hcaca;
    LUT4 i15682_3_lut (.A(\result_r[6] [6]), .B(\result_r[7] [6]), .C(y_1_delay[0]), 
         .Z(n34066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15682_3_lut.init = 16'hcaca;
    LUT4 i15681_3_lut (.A(\result_r[4] [6]), .B(\result_r[5] [6]), .C(y_1_delay[0]), 
         .Z(n34065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15681_3_lut.init = 16'hcaca;
    LUT4 i15680_3_lut (.A(\result_r[2] [6]), .B(\result_r[3] [6]), .C(y_1_delay[0]), 
         .Z(n34064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15680_3_lut.init = 16'hcaca;
    LUT4 i15679_3_lut (.A(\result_r[0] [6]), .B(\result_r[1] [6]), .C(y_1_delay[0]), 
         .Z(n34063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15679_3_lut.init = 16'hcaca;
    LUT4 i14936_3_lut (.A(\result_i[2] [15]), .B(\result_i[3] [15]), .C(y_1_delay[0]), 
         .Z(n33320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14936_3_lut.init = 16'hcaca;
    LUT4 i14935_3_lut (.A(\result_i[0] [15]), .B(\result_i[1] [15]), .C(y_1_delay[0]), 
         .Z(n33319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14935_3_lut.init = 16'hcaca;
    LUT4 i15062_3_lut (.A(\result_i[6] [11]), .B(\result_i[7] [11]), .C(y_1_delay[0]), 
         .Z(n33446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15062_3_lut.init = 16'hcaca;
    LUT4 i15061_3_lut (.A(\result_i[4] [11]), .B(\result_i[5] [11]), .C(y_1_delay[0]), 
         .Z(n33445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15061_3_lut.init = 16'hcaca;
    LUT4 i15060_3_lut (.A(\result_i[2] [11]), .B(\result_i[3] [11]), .C(y_1_delay[0]), 
         .Z(n33444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15060_3_lut.init = 16'hcaca;
    LUT4 i15059_3_lut (.A(\result_i[0] [11]), .B(\result_i[1] [11]), .C(y_1_delay[0]), 
         .Z(n33443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15059_3_lut.init = 16'hcaca;
    LUT4 i14943_3_lut (.A(\result_i[16] [15]), .B(\result_i[17] [15]), .C(y_1_delay[0]), 
         .Z(n33327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14943_3_lut.init = 16'hcaca;
    LUT4 i14944_3_lut (.A(\result_i[18] [15]), .B(\result_i[19] [15]), .C(y_1_delay[0]), 
         .Z(n33328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14944_3_lut.init = 16'hcaca;
    LUT4 i6745_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[490])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6745_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_2_lut_4_lut_4_lut_4_lut (.A(count_y[4]), .B(n34771), .C(n34770), 
         .D(count_y[3]), .Z(n32944)) /* synthesis lut_function=(A (C (D))+!A !((C+(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_4_lut_4_lut_4_lut.init = 16'ha004;
    LUT4 i3809_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[346])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3809_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3801_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[347])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3801_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3793_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[348])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3793_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3785_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[349])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3785_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3777_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[350])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3777_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3769_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_i[10] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[351])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3769_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7977_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[336])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7977_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7969_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[337])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7969_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7961_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[338])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7961_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7953_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[339])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7953_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7945_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[340])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7945_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7937_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[341])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7937_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7929_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[342])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7929_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7921_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[343])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7921_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7913_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[344])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7913_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2623_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[494])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2623_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i7905_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[345])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7905_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7897_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[346])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7897_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7889_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[347])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7889_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7881_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[348])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7881_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7873_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[349])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7873_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7865_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[350])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7865_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7857_3_lut_4_lut (.A(n34717), .B(n34707), .C(\result_r[10] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[351])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7857_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14946_3_lut (.A(\result_i[22] [15]), .B(\result_i[23] [15]), .C(y_1_delay[0]), 
         .Z(n33330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14946_3_lut.init = 16'hcaca;
    LUT4 i4017_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[320])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4017_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4009_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[321])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4009_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2615_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[495])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2615_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i14076_2_lut (.A(n8849), .B(n89_adj_7291), .Z(op_i_23__N_1310_adj_7380[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14076_2_lut.init = 16'h6666;
    LUT4 i849_4_lut_rep_442 (.A(count_y[1]), .B(count_y[3]), .C(count_y[0]), 
         .D(n32925), .Z(n34812)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i849_4_lut_rep_442.init = 16'ha5a6;
    LUT4 i1_2_lut_rep_369_3_lut_4_lut_4_lut_4_lut (.A(count_y[1]), .B(count_y[3]), 
         .C(count_y[0]), .D(n32925), .Z(n34731)) /* synthesis lut_function=(!(A+(B (C)+!B (C+!(D))))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_369_3_lut_4_lut_4_lut_4_lut.init = 16'h0504;
    LUT4 i14079_2_lut (.A(n8721), .B(n89), .Z(op_i_23__N_1310_adj_7329[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14079_2_lut.init = 16'h6666;
    LUT4 i14080_2_lut (.A(n9105), .B(n89_adj_6552), .Z(op_i_23__N_1310_adj_7491[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14080_2_lut.init = 16'h6666;
    LUT4 i14078_2_lut (.A(n8977), .B(n89_adj_7261), .Z(op_i_23__N_1310_adj_7435[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14078_2_lut.init = 16'h6666;
    LUT4 i15399_3_lut (.A(n33781), .B(n33782), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15399_3_lut.init = 16'hcaca;
    LUT4 i15368_3_lut (.A(n33750), .B(n33751), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15368_3_lut.init = 16'hcaca;
    LUT4 i15337_3_lut (.A(n33719), .B(n33720), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15337_3_lut.init = 16'hcaca;
    LUT4 i15306_3_lut (.A(n33688), .B(n33689), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15306_3_lut.init = 16'hcaca;
    LUT4 i15275_3_lut (.A(n33657), .B(n33658), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15275_3_lut.init = 16'hcaca;
    LUT4 i15244_3_lut (.A(n33626), .B(n33627), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15244_3_lut.init = 16'hcaca;
    LUT4 i15213_3_lut (.A(n33595), .B(n33596), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15213_3_lut.init = 16'hcaca;
    LUT4 i15182_3_lut (.A(n33564), .B(n33565), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15182_3_lut.init = 16'hcaca;
    LUT4 i15151_3_lut (.A(n33533), .B(n33534), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15151_3_lut.init = 16'hcaca;
    LUT4 i15120_3_lut (.A(n33502), .B(n33503), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15120_3_lut.init = 16'hcaca;
    LUT4 i15089_3_lut (.A(n33471), .B(n33472), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15089_3_lut.init = 16'hcaca;
    LUT4 i15058_3_lut (.A(n33440), .B(n33441), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15058_3_lut.init = 16'hcaca;
    LUT4 i15027_3_lut (.A(n33409), .B(n33410), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15027_3_lut.init = 16'hcaca;
    LUT4 i14996_3_lut (.A(n33378), .B(n33379), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14996_3_lut.init = 16'hcaca;
    LUT4 i14965_3_lut (.A(n33347), .B(n33348), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14965_3_lut.init = 16'hcaca;
    LUT4 i15864_3_lut (.A(n34246), .B(n34247), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15864_3_lut.init = 16'hcaca;
    LUT4 i14092_2_lut (.A(s_count_adj_7402[0]), .B(state_1__N_5502), .Z(n30041)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(33[24:35])
    defparam i14092_2_lut.init = 16'h6666;
    LUT4 i12330_4_lut (.A(s_count[3]), .B(s_count[2]), .C(clk_c_enable_2285), 
         .D(n34785), .Z(n30040)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam i12330_4_lut.init = 16'h6aaa;
    LUT4 i15833_3_lut (.A(n34215), .B(n34216), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15833_3_lut.init = 16'hcaca;
    LUT4 i15802_3_lut (.A(n34184), .B(n34185), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15802_3_lut.init = 16'hcaca;
    LUT4 i15771_3_lut (.A(n34153), .B(n34154), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15771_3_lut.init = 16'hcaca;
    LUT4 i15740_3_lut (.A(n34122), .B(n34123), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15740_3_lut.init = 16'hcaca;
    LUT4 i15709_3_lut (.A(n34091), .B(n34092), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15709_3_lut.init = 16'hcaca;
    LUT4 i15678_3_lut (.A(n34060), .B(n34061), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15678_3_lut.init = 16'hcaca;
    LUT4 i15647_3_lut (.A(n34029), .B(n34030), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15647_3_lut.init = 16'hcaca;
    LUT4 i15616_3_lut (.A(n33998), .B(n33999), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15616_3_lut.init = 16'hcaca;
    LUT4 i15585_3_lut (.A(n33967), .B(n33968), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15585_3_lut.init = 16'hcaca;
    LUT4 i15554_3_lut (.A(n33936), .B(n33937), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15554_3_lut.init = 16'hcaca;
    LUT4 i15523_3_lut (.A(n33905), .B(n33906), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15523_3_lut.init = 16'hcaca;
    LUT4 i15492_3_lut (.A(n33874), .B(n33875), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15492_3_lut.init = 16'hcaca;
    LUT4 i15461_3_lut (.A(n33843), .B(n33844), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15461_3_lut.init = 16'hcaca;
    LUT4 i15430_3_lut (.A(n33812), .B(n33813), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15430_3_lut.init = 16'hcaca;
    LUT4 i2344_2_lut (.A(s5_count), .B(r4_valid), .Z(n19995)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam i2344_2_lut.init = 16'h6666;
    LUT4 i14903_3_lut (.A(n33285), .B(n33286), .C(y_1_delay[4]), .Z(next_dout_i_15__N_1045[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14903_3_lut.init = 16'hcaca;
    LUT4 i4001_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[322])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4001_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3993_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[323])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3993_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15534_3_lut (.A(\result_r[20] [11]), .B(\result_r[21] [11]), .C(y_1_delay[0]), 
         .Z(n33918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15534_3_lut.init = 16'hcaca;
    LUT4 i3985_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[324])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3985_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3977_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[325])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3977_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15190_3_lut (.A(\result_i[14] [7]), .B(\result_i[15] [7]), .C(y_1_delay[0]), 
         .Z(n33574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15190_3_lut.init = 16'hcaca;
    LUT4 i3969_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[326])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3969_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3961_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[327])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3961_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3953_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[328])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3953_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3945_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[329])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3945_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3937_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[330])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3937_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3929_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[331])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3929_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3921_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[332])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3921_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15189_3_lut (.A(\result_i[12] [7]), .B(\result_i[13] [7]), .C(y_1_delay[0]), 
         .Z(n33573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15189_3_lut.init = 16'hcaca;
    LUT4 i3913_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[333])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3913_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3905_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[334])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3905_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3897_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_i[11] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[335])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i3897_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8105_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[320])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8105_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8097_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[321])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8097_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8089_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[322])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8089_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8081_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[323])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8081_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8073_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[324])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8073_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i14934_3_lut (.A(n33316), .B(n33317), .C(y_1_delay[4]), .Z(next_dout_r_15__N_1029[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14934_3_lut.init = 16'hcaca;
    LUT4 i8065_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[325])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8065_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15188_3_lut (.A(\result_i[10] [7]), .B(\result_i[11] [7]), .C(y_1_delay[0]), 
         .Z(n33572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15188_3_lut.init = 16'hcaca;
    LUT4 i8057_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[326])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8057_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8049_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[327])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8049_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15187_3_lut (.A(\result_i[8] [7]), .B(\result_i[9] [7]), .C(y_1_delay[0]), 
         .Z(n33571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15187_3_lut.init = 16'hcaca;
    LUT4 i8041_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[328])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8041_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8033_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[329])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8033_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8025_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[330])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8025_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8017_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[331])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8017_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8009_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[332])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8009_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15283_3_lut (.A(\result_i[14] [4]), .B(\result_i[15] [4]), .C(y_1_delay[0]), 
         .Z(n33667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15283_3_lut.init = 16'hcaca;
    LUT4 i8001_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[333])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8001_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i7993_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[334])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7993_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i7985_3_lut_4_lut (.A(n30503), .B(n34704), .C(\result_r[11] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[335])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i7985_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4145_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[304])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4145_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4137_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[305])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4137_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4129_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[306])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4129_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15533_3_lut (.A(\result_r[18] [11]), .B(\result_r[19] [11]), .C(y_1_delay[0]), 
         .Z(n33917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15533_3_lut.init = 16'hcaca;
    LUT4 i4121_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[307])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4121_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4113_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[308])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4113_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4105_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[309])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4105_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15532_3_lut (.A(\result_r[16] [11]), .B(\result_r[17] [11]), .C(y_1_delay[0]), 
         .Z(n33916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15532_3_lut.init = 16'hcaca;
    LUT4 i4097_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[310])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4097_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4089_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[311])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4089_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4081_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[312])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4081_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15186_3_lut (.A(\result_i[6] [7]), .B(\result_i[7] [7]), .C(y_1_delay[0]), 
         .Z(n33570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15186_3_lut.init = 16'hcaca;
    LUT4 i4073_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[313])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4073_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4065_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[314])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4065_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15185_3_lut (.A(\result_i[4] [7]), .B(\result_i[5] [7]), .C(y_1_delay[0]), 
         .Z(n33569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15185_3_lut.init = 16'hcaca;
    LUT4 i4057_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[315])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4057_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4049_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[316])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4049_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15282_3_lut (.A(\result_i[12] [4]), .B(\result_i[13] [4]), .C(y_1_delay[0]), 
         .Z(n33666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15282_3_lut.init = 16'hcaca;
    LUT4 i4041_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[317])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4041_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4033_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[318])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4033_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4025_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_i[12] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[319])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4025_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8233_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[304])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8233_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8225_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[305])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8225_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8217_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[306])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8217_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8209_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[307])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8209_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8201_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[308])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8201_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8193_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[309])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8193_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8185_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[310])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8185_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8177_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[311])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8177_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8169_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[312])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8169_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15184_3_lut (.A(\result_i[2] [7]), .B(\result_i[3] [7]), .C(y_1_delay[0]), 
         .Z(n33568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15184_3_lut.init = 16'hcaca;
    LUT4 i15183_3_lut (.A(\result_i[0] [7]), .B(\result_i[1] [7]), .C(y_1_delay[0]), 
         .Z(n33567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15183_3_lut.init = 16'hcaca;
    LUT4 i8161_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[313])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8161_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8153_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[314])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8153_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8145_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[315])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8145_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8137_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[316])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8137_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15512 (.BLUT(n33883), .ALUT(n33884), .C0(y_1_delay[1]), .Z(n33896));
    LUT4 i8129_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[317])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8129_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15513 (.BLUT(n33885), .ALUT(n33886), .C0(y_1_delay[1]), .Z(n33897));
    LUT4 i8121_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[318])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8121_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8113_3_lut_4_lut (.A(n30503), .B(n34705), .C(\result_r[12] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[319])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8113_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4273_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[288])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4273_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4265_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[289])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4265_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15531_3_lut (.A(\result_r[14] [11]), .B(\result_r[15] [11]), .C(y_1_delay[0]), 
         .Z(n33915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15531_3_lut.init = 16'hcaca;
    LUT4 i15530_3_lut (.A(\result_r[12] [11]), .B(\result_r[13] [11]), .C(y_1_delay[0]), 
         .Z(n33914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15530_3_lut.init = 16'hcaca;
    LUT4 i15818_3_lut (.A(\result_r[30] [2]), .B(\result_r[31] [2]), .C(y_1_delay[0]), 
         .Z(n34202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15818_3_lut.init = 16'hcaca;
    LUT4 i4257_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[290])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4257_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4249_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[291])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4249_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4241_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[292])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4241_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4233_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[293])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4233_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4225_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[294])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4225_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4217_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[295])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4217_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4209_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[296])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4209_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15817_3_lut (.A(\result_r[28] [2]), .B(\result_r[29] [2]), .C(y_1_delay[0]), 
         .Z(n34201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15817_3_lut.init = 16'hcaca;
    LUT4 i4201_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[297])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4201_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15281_3_lut (.A(\result_i[10] [4]), .B(\result_i[11] [4]), .C(y_1_delay[0]), 
         .Z(n33665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15281_3_lut.init = 16'hcaca;
    LUT4 i4193_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[298])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4193_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15816_3_lut (.A(\result_r[26] [2]), .B(\result_r[27] [2]), .C(y_1_delay[0]), 
         .Z(n34200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15816_3_lut.init = 16'hcaca;
    LUT4 i15815_3_lut (.A(\result_r[24] [2]), .B(\result_r[25] [2]), .C(y_1_delay[0]), 
         .Z(n34199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15815_3_lut.init = 16'hcaca;
    PFUMX i15514 (.BLUT(n33887), .ALUT(n33888), .C0(y_1_delay[1]), .Z(n33898));
    LUT4 i14065_2_lut (.A(shift_2_dout_i[0]), .B(shift_2_dout_r[0]), .Z(n126)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14065_2_lut.init = 16'h6666;
    LUT4 i4185_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[299])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4185_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15280_3_lut (.A(\result_i[8] [4]), .B(\result_i[9] [4]), .C(y_1_delay[0]), 
         .Z(n33664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15280_3_lut.init = 16'hcaca;
    LUT4 i4177_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[300])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4177_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4169_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[301])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4169_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15814_3_lut (.A(\result_r[22] [2]), .B(\result_r[23] [2]), .C(y_1_delay[0]), 
         .Z(n34198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15814_3_lut.init = 16'hcaca;
    LUT4 i15813_3_lut (.A(\result_r[20] [2]), .B(\result_r[21] [2]), .C(y_1_delay[0]), 
         .Z(n34197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15813_3_lut.init = 16'hcaca;
    LUT4 i15812_3_lut (.A(\result_r[18] [2]), .B(\result_r[19] [2]), .C(y_1_delay[0]), 
         .Z(n34196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15812_3_lut.init = 16'hcaca;
    LUT4 i4161_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[302])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4161_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15515 (.BLUT(n33889), .ALUT(n33890), .C0(y_1_delay[1]), .Z(n33899));
    LUT4 i4153_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_i[13] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[303])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4153_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8361_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[288])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8361_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15811_3_lut (.A(\result_r[16] [2]), .B(\result_r[17] [2]), .C(y_1_delay[0]), 
         .Z(n34195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15811_3_lut.init = 16'hcaca;
    LUT4 i8353_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[289])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8353_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8345_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[290])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8345_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15292 (.BLUT(n33660), .ALUT(n33661), .C0(y_1_delay[1]), .Z(n33676));
    LUT4 i15810_3_lut (.A(\result_r[14] [2]), .B(\result_r[15] [2]), .C(y_1_delay[0]), 
         .Z(n34194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15810_3_lut.init = 16'hcaca;
    PFUMX i15516 (.BLUT(n33891), .ALUT(n33892), .C0(y_1_delay[1]), .Z(n33900));
    LUT4 i8337_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[291])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8337_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8329_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[292])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8329_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15663_3_lut (.A(\result_r[30] [7]), .B(\result_r[31] [7]), .C(y_1_delay[0]), 
         .Z(n34047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15663_3_lut.init = 16'hcaca;
    LUT4 i8321_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[293])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8321_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8313_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[294])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8313_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15809_3_lut (.A(\result_r[12] [2]), .B(\result_r[13] [2]), .C(y_1_delay[0]), 
         .Z(n34193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15809_3_lut.init = 16'hcaca;
    LUT4 i8305_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[295])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8305_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8297_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[296])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8297_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15788 (.BLUT(n34156), .ALUT(n34157), .C0(y_1_delay[1]), .Z(n34172));
    LUT4 i8289_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[297])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8289_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8281_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[298])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8281_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i14060_2_lut (.A(shift_4_dout_i[0]), .B(shift_4_dout_r[0]), .Z(n126_adj_7267)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14060_2_lut.init = 16'h6666;
    LUT4 i8273_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[299])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8273_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8265_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[300])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8265_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8257_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[301])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8257_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15808_3_lut (.A(\result_r[10] [2]), .B(\result_r[11] [2]), .C(y_1_delay[0]), 
         .Z(n34192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15808_3_lut.init = 16'hcaca;
    LUT4 i8249_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[302])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8249_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8241_3_lut_4_lut (.A(n30503), .B(n34706), .C(\result_r[13] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[303])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8241_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4401_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[272])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4401_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15807_3_lut (.A(\result_r[8] [2]), .B(\result_r[9] [2]), .C(y_1_delay[0]), 
         .Z(n34191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15807_3_lut.init = 16'hcaca;
    PFUMX i15789 (.BLUT(n34158), .ALUT(n34159), .C0(y_1_delay[1]), .Z(n34173));
    LUT4 i15662_3_lut (.A(\result_r[28] [7]), .B(\result_r[29] [7]), .C(y_1_delay[0]), 
         .Z(n34046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15662_3_lut.init = 16'hcaca;
    LUT4 i4393_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[273])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4393_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4385_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[274])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4385_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4377_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[275])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4377_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4369_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[276])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4369_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4361_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[277])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4361_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4353_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[278])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4353_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4345_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[279])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4345_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4337_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[280])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4337_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4329_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[281])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4329_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i14077_2_lut (.A(n8593), .B(n89_adj_7164), .Z(op_i_23__N_1310[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i14077_2_lut.init = 16'h6666;
    LUT4 i4321_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[282])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4321_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4313_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[283])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4313_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4305_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[284])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4305_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15806_3_lut (.A(\result_r[6] [2]), .B(\result_r[7] [2]), .C(y_1_delay[0]), 
         .Z(n34190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15806_3_lut.init = 16'hcaca;
    LUT4 i4297_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[285])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4297_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4289_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[286])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4289_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15805_3_lut (.A(\result_r[4] [2]), .B(\result_r[5] [2]), .C(y_1_delay[0]), 
         .Z(n34189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15805_3_lut.init = 16'hcaca;
    LUT4 i4281_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_i[14] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[287])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4281_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_990_add_4_6 (.A0(op_i_23__N_1154[4]), .B0(op_r_23__N_1106[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[5]), .B1(op_r_23__N_1106[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32057), .COUT(n32058), .S0(n9987), 
          .S1(n9988));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_16 (.A0(n9091), .B0(n75_adj_6566), .C0(GND_net), 
          .D0(VCC_net), .A1(n9090), .B1(n74_adj_6567), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32355), .COUT(n32356), .S0(op_i_23__N_1310_adj_7491[20]), 
          .S1(op_i_23__N_1310_adj_7491[21]));
    defparam _add_1_1086_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_4 (.A0(op_i_23__N_1154[2]), .B0(op_r_23__N_1106[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[3]), .B1(op_r_23__N_1106[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32056), .COUT(n32057), .S0(n9985), 
          .S1(n9986));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_2 (.A0(op_i_23__N_1154[0]), .B0(op_r_23__N_1106[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[1]), .B1(op_r_23__N_1106[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32056), .S1(n9984));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_990_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_990_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_14 (.A0(n9093), .B0(n77_adj_6564), .C0(GND_net), 
          .D0(VCC_net), .A1(n9092), .B1(n76_adj_6565), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32354), .COUT(n32355), .S0(op_i_23__N_1310_adj_7491[18]), 
          .S1(op_i_23__N_1310_adj_7491[19]));
    defparam _add_1_1086_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_14.INJECT1_1 = "NO";
    LUT4 i8489_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[272])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8489_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1001_add_4_32 (.A0(op_r_23__N_1268[30]), .B0(op_r_23__N_1226[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[31]), .B1(op_r_23__N_1226[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32053), .S0(op_r_23__N_1082[30]), 
          .S1(op_r_23__N_1082[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_12 (.A0(n9095), .B0(n79_adj_6562), .C0(GND_net), 
          .D0(VCC_net), .A1(n9094), .B1(n78_adj_6563), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32353), .COUT(n32354), .S0(op_i_23__N_1310_adj_7491[16]), 
          .S1(op_i_23__N_1310_adj_7491[17]));
    defparam _add_1_1086_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_30 (.A0(op_r_23__N_1268[28]), .B0(op_r_23__N_1226[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[29]), .B1(op_r_23__N_1226[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32052), .COUT(n32053), .S0(op_r_23__N_1082[28]), 
          .S1(op_r_23__N_1082[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_28 (.A0(op_r_23__N_1268[26]), .B0(op_r_23__N_1226[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[27]), .B1(op_r_23__N_1226[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32051), .COUT(n32052), .S0(op_r_23__N_1082[26]), 
          .S1(op_r_23__N_1082[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_10 (.A0(n9097), .B0(n81_adj_6560), .C0(GND_net), 
          .D0(VCC_net), .A1(n9096), .B1(n80_adj_6561), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32352), .COUT(n32353), .S0(op_i_23__N_1310_adj_7491[14]), 
          .S1(op_i_23__N_1310_adj_7491[15]));
    defparam _add_1_1086_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_10.INJECT1_1 = "NO";
    PFUMX i15790 (.BLUT(n34160), .ALUT(n34161), .C0(y_1_delay[1]), .Z(n34174));
    CCU2C _add_1_1001_add_4_26 (.A0(op_r_23__N_1268[24]), .B0(op_r_23__N_1226[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[25]), .B1(op_r_23__N_1226[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32050), .COUT(n32051), .S0(op_r_23__N_1082[24]), 
          .S1(op_r_23__N_1082[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_24 (.A0(op_r_23__N_1268[22]), .B0(op_r_23__N_1226[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[23]), .B1(op_r_23__N_1226[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32049), .COUT(n32050), .S0(op_r_23__N_1082[22]), 
          .S1(op_r_23__N_1082[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_8 (.A0(n9099), .B0(n83_adj_6558), .C0(GND_net), 
          .D0(VCC_net), .A1(n9098), .B1(n82_adj_6559), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32351), .COUT(n32352), .S0(op_i_23__N_1310_adj_7491[12]), 
          .S1(op_i_23__N_1310_adj_7491[13]));
    defparam _add_1_1086_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_22 (.A0(op_r_23__N_1268[20]), .B0(op_r_23__N_1226[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[21]), .B1(op_r_23__N_1226[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32048), .COUT(n32049), .S0(op_r_23__N_1082[20]), 
          .S1(op_r_23__N_1082[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_20 (.A0(op_r_23__N_1268[18]), .B0(op_r_23__N_1226[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[19]), .B1(op_r_23__N_1226[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32047), .COUT(n32048), .S0(op_r_23__N_1082[18]), 
          .S1(op_r_23__N_1082[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_6 (.A0(n9101), .B0(n85_adj_6556), .C0(GND_net), 
          .D0(VCC_net), .A1(n9100), .B1(n84_adj_6557), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32350), .COUT(n32351), .S0(op_i_23__N_1310_adj_7491[10]), 
          .S1(op_i_23__N_1310_adj_7491[11]));
    defparam _add_1_1086_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_6.INJECT1_1 = "NO";
    LUT4 i8481_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[273])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8481_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1001_add_4_18 (.A0(op_r_23__N_1268[16]), .B0(op_r_23__N_1226[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[17]), .B1(op_r_23__N_1226[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32046), .COUT(n32047), .S0(op_r_23__N_1082[16]), 
          .S1(op_r_23__N_1082[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_16 (.A0(op_r_23__N_1268[14]), .B0(op_r_23__N_1226[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[15]), .B1(op_r_23__N_1226[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32045), .COUT(n32046), .S0(op_r_23__N_1082[14]), 
          .S1(op_r_23__N_1082[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_4 (.A0(n9103), .B0(n87_adj_6554), .C0(GND_net), 
          .D0(VCC_net), .A1(n9102), .B1(n86_adj_6555), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32349), .COUT(n32350), .S0(op_i_23__N_1310_adj_7491[8]), 
          .S1(op_i_23__N_1310_adj_7491[9]));
    defparam _add_1_1086_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1086_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_14 (.A0(op_r_23__N_1268[12]), .B0(op_r_23__N_1226[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[13]), .B1(op_r_23__N_1226[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32044), .COUT(n32045), .S0(op_r_23__N_1082[12]), 
          .S1(op_r_23__N_1082[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_12 (.A0(op_r_23__N_1268[10]), .B0(op_r_23__N_1226[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[11]), .B1(op_r_23__N_1226[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32043), .COUT(n32044), .S0(op_r_23__N_1082[10]), 
          .S1(op_r_23__N_1082[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1086_add_4_2 (.A0(n9105), .B0(n89_adj_6552), .C0(GND_net), 
          .D0(VCC_net), .A1(n9104), .B1(n88_adj_6553), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32349), .S1(op_i_23__N_1310_adj_7491[7]));
    defparam _add_1_1086_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1086_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1086_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1086_add_4_2.INJECT1_1 = "NO";
    LUT4 i8473_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[274])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8473_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8465_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[275])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8465_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1001_add_4_10 (.A0(op_r_23__N_1268[8]), .B0(op_r_23__N_1226[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[9]), .B1(op_r_23__N_1226[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32042), .COUT(n32043), .S0(op_r_23__N_1082[8]), 
          .S1(op_r_23__N_1082[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_8 (.A0(op_r_23__N_1268[6]), .B0(op_r_23__N_1226[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[7]), .B1(op_r_23__N_1226[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32041), .COUT(n32042));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_6 (.A0(op_r_23__N_1268[4]), .B0(op_r_23__N_1226[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[5]), .B1(op_r_23__N_1226[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32040), .COUT(n32041));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_18 (.A0(din_i_reg[23]), .B0(shift_16_dout_i[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n32347), .S0(delay_i_23__N_1202[23]));
    defparam _add_1_1134_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_18.INIT1 = 16'h0000;
    defparam _add_1_1134_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_18.INJECT1_1 = "NO";
    LUT4 i8457_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[276])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8457_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1001_add_4_4 (.A0(op_r_23__N_1268[2]), .B0(op_r_23__N_1226[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[3]), .B1(op_r_23__N_1226[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32039), .COUT(n32040));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1001_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1001_add_4_2 (.A0(op_r_23__N_1268[0]), .B0(op_r_23__N_1226[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268[1]), .B1(op_r_23__N_1226[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32039));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1001_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1001_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1001_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1001_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_16 (.A0(din_i_reg[23]), .B0(shift_16_dout_i[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[23]), .B1(shift_16_dout_i[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32346), .COUT(n32347), .S0(delay_i_23__N_1202[21]), 
          .S1(delay_i_23__N_1202[22]));
    defparam _add_1_1134_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_25 (.A0(n31574), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[22]), .A1(n31572), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[23]), .CIN(n32037), .S0(op_r_23__N_1106_adj_7319[22]), 
          .S1(op_r_23__N_1106_adj_7319[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_25.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_25.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_14 (.A0(din_i_reg[23]), .B0(shift_16_dout_i[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[23]), .B1(shift_16_dout_i[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32345), .COUT(n32346), .S0(delay_i_23__N_1202[19]), 
          .S1(delay_i_23__N_1202[20]));
    defparam _add_1_1134_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_23 (.A0(n31578), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[20]), .A1(n31576), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[21]), .CIN(n32036), .COUT(n32037), .S0(op_r_23__N_1106_adj_7319[20]), 
          .S1(op_r_23__N_1106_adj_7319[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_23.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_23.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_21 (.A0(n31582), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[18]), .A1(n31580), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[19]), .CIN(n32035), .COUT(n32036), .S0(op_r_23__N_1106_adj_7319[18]), 
          .S1(op_r_23__N_1106_adj_7319[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_21.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_21.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_12 (.A0(din_i_reg[17]), .B0(shift_16_dout_i[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[18]), .B1(shift_16_dout_i[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32344), .COUT(n32345), .S0(delay_i_23__N_1202[17]), 
          .S1(delay_i_23__N_1202[18]));
    defparam _add_1_1134_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_19 (.A0(n31586), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[16]), .A1(n31584), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[17]), .CIN(n32034), .COUT(n32035), .S0(op_r_23__N_1106_adj_7319[16]), 
          .S1(op_r_23__N_1106_adj_7319[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_19.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_19.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_17 (.A0(n31590), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[14]), .A1(n31588), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[15]), .CIN(n32033), .COUT(n32034), .S0(op_r_23__N_1106_adj_7319[14]), 
          .S1(op_r_23__N_1106_adj_7319[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_17.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_17.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_10 (.A0(din_i_reg[15]), .B0(shift_16_dout_i[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[16]), .B1(shift_16_dout_i[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32343), .COUT(n32344), .S0(delay_i_23__N_1202[15]), 
          .S1(delay_i_23__N_1202[16]));
    defparam _add_1_1134_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_10.INJECT1_1 = "NO";
    LUT4 i8449_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[277])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8449_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1004_add_4_15 (.A0(n31594), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[12]), .A1(n31592), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[13]), .CIN(n32032), .COUT(n32033), .S0(op_r_23__N_1106_adj_7319[12]), 
          .S1(op_r_23__N_1106_adj_7319[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_15.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_15.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_13 (.A0(n31598), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[10]), .A1(n31596), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[11]), .CIN(n32031), .COUT(n32032), .S0(op_r_23__N_1106_adj_7319[10]), 
          .S1(op_r_23__N_1106_adj_7319[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_13.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_13.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_8 (.A0(din_i_reg[13]), .B0(shift_16_dout_i[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[14]), .B1(shift_16_dout_i[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32342), .COUT(n32343), .S0(delay_i_23__N_1202[13]), 
          .S1(delay_i_23__N_1202[14]));
    defparam _add_1_1134_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_11 (.A0(n31602), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[8]), .A1(n31600), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[9]), .CIN(n32030), .COUT(n32031), .S0(op_r_23__N_1106_adj_7319[8]), 
          .S1(op_r_23__N_1106_adj_7319[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_11.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_11.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_9 (.A0(n31606), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[6]), .A1(n31604), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[7]), .CIN(n32029), .COUT(n32030), .S0(op_r_23__N_1106_adj_7319[6]), 
          .S1(op_r_23__N_1106_adj_7319[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_9.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_9.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_6 (.A0(din_i_reg[11]), .B0(shift_16_dout_i[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[12]), .B1(shift_16_dout_i[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32341), .COUT(n32342), .S0(delay_i_23__N_1202[11]), 
          .S1(delay_i_23__N_1202[12]));
    defparam _add_1_1134_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_6.INJECT1_1 = "NO";
    PFUMX i15791 (.BLUT(n34162), .ALUT(n34163), .C0(y_1_delay[1]), .Z(n34175));
    LUT4 i15804_3_lut (.A(\result_r[2] [2]), .B(\result_r[3] [2]), .C(y_1_delay[0]), 
         .Z(n34188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15804_3_lut.init = 16'hcaca;
    CCU2C _add_1_1004_add_4_7 (.A0(n31610), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[4]), .A1(n31608), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[5]), .CIN(n32028), .COUT(n32029), .S0(op_r_23__N_1106_adj_7319[4]), 
          .S1(op_r_23__N_1106_adj_7319[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_7.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_7.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_4 (.A0(din_i_reg[9]), .B0(shift_16_dout_i[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_i_reg[10]), .B1(shift_16_dout_i[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32340), .COUT(n32341), .S0(delay_i_23__N_1202[9]), 
          .S1(delay_i_23__N_1202[10]));
    defparam _add_1_1134_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1134_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_5 (.A0(n31614), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[2]), .A1(n31612), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[3]), .CIN(n32027), .COUT(n32028), .S0(op_r_23__N_1106_adj_7319[2]), 
          .S1(op_r_23__N_1106_adj_7319[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_5.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_5.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1004_add_4_3 (.A0(n31618), .B0(rom8_state[0]), .C0(n34794), 
          .D0(shift_8_dout_r[0]), .A1(n31616), .B1(rom8_state[0]), .C1(n34794), 
          .D1(shift_8_dout_r[1]), .CIN(n32026), .COUT(n32027), .S0(op_r_23__N_1106_adj_7319[0]), 
          .S1(op_r_23__N_1106_adj_7319[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_3.INIT0 = 16'h65aa;
    defparam _add_1_1004_add_4_3.INIT1 = 16'h65aa;
    defparam _add_1_1004_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1134_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(din_i_reg[8]), .B1(shift_16_dout_i[8]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32340), .S1(delay_i_23__N_1202[8]));
    defparam _add_1_1134_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1134_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1134_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1134_add_4_2.INJECT1_1 = "NO";
    LUT4 i15803_3_lut (.A(\result_r[0] [2]), .B(\result_r[1] [2]), .C(y_1_delay[0]), 
         .Z(n34187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15803_3_lut.init = 16'hcaca;
    CCU2C _add_1_1004_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(rom8_state[0]), .B1(n29822), .C1(n29823), 
          .D1(n29824), .COUT(n32026));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1004_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1004_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1004_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1004_add_4_1.INJECT1_1 = "NO";
    LUT4 i15529_3_lut (.A(\result_r[10] [11]), .B(\result_r[11] [11]), .C(y_1_delay[0]), 
         .Z(n33913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15529_3_lut.init = 16'hcaca;
    CCU2C _add_1_1081_add_4_32 (.A0(op_r_23__N_1268_adj_7486[30]), .B0(op_i_23__N_1310_adj_7491[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[31]), 
          .B1(op_i_23__N_1310_adj_7491[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32338), .S0(op_i_23__N_1130_adj_7492[30]), .S1(op_i_23__N_1130_adj_7492[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_26 (.A0(shift_2_dout_i[23]), .B0(shift_2_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n32022), .S0(n319_adj_6944));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1045_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_24 (.A0(shift_2_dout_i[22]), .B0(shift_2_dout_r[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[23]), .B1(shift_2_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32021), .COUT(n32022), .S0(n11142), 
          .S1(n11143));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_30 (.A0(op_r_23__N_1268_adj_7486[28]), .B0(op_i_23__N_1310_adj_7491[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[29]), 
          .B1(op_i_23__N_1310_adj_7491[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32337), .COUT(n32338), .S0(op_i_23__N_1130_adj_7492[28]), 
          .S1(op_i_23__N_1130_adj_7492[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_22 (.A0(shift_2_dout_i[20]), .B0(shift_2_dout_r[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[21]), .B1(shift_2_dout_r[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32020), .COUT(n32021), .S0(n11140), 
          .S1(n11141));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_20 (.A0(shift_2_dout_i[18]), .B0(shift_2_dout_r[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[19]), .B1(shift_2_dout_r[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32019), .COUT(n32020), .S0(n11138), 
          .S1(n11139));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_28 (.A0(op_r_23__N_1268_adj_7486[26]), .B0(op_i_23__N_1310_adj_7491[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[27]), 
          .B1(op_i_23__N_1310_adj_7491[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32336), .COUT(n32337), .S0(op_i_23__N_1130_adj_7492[26]), 
          .S1(op_i_23__N_1130_adj_7492[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_18 (.A0(shift_2_dout_i[16]), .B0(shift_2_dout_r[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[17]), .B1(shift_2_dout_r[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32018), .COUT(n32019), .S0(n11136), 
          .S1(n11137));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_16 (.A0(shift_2_dout_i[14]), .B0(shift_2_dout_r[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[15]), .B1(shift_2_dout_r[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32017), .COUT(n32018), .S0(n11134), 
          .S1(n11135));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_26 (.A0(op_r_23__N_1268_adj_7486[24]), .B0(op_i_23__N_1310_adj_7491[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[25]), 
          .B1(op_i_23__N_1310_adj_7491[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32335), .COUT(n32336), .S0(op_i_23__N_1130_adj_7492[24]), 
          .S1(op_i_23__N_1130_adj_7492[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_26.INJECT1_1 = "NO";
    LUT4 i8441_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[278])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8441_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1045_add_4_14 (.A0(shift_2_dout_i[12]), .B0(shift_2_dout_r[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[13]), .B1(shift_2_dout_r[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32016), .COUT(n32017), .S0(n11132), 
          .S1(n11133));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_12 (.A0(shift_2_dout_i[10]), .B0(shift_2_dout_r[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[11]), .B1(shift_2_dout_r[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32015), .COUT(n32016), .S0(n11130), 
          .S1(n11131));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_24 (.A0(op_r_23__N_1268_adj_7486[22]), .B0(op_i_23__N_1310_adj_7491[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[23]), 
          .B1(op_i_23__N_1310_adj_7491[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32334), .COUT(n32335), .S0(op_i_23__N_1130_adj_7492[22]), 
          .S1(op_i_23__N_1130_adj_7492[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_10 (.A0(shift_2_dout_i[8]), .B0(shift_2_dout_r[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[9]), .B1(shift_2_dout_r[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32014), .COUT(n32015), .S0(n11128), 
          .S1(n11129));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_8 (.A0(shift_2_dout_i[6]), .B0(shift_2_dout_r[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[7]), .B1(shift_2_dout_r[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32013), .COUT(n32014), .S0(n11126), 
          .S1(n11127));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_22 (.A0(op_r_23__N_1268_adj_7486[20]), .B0(op_i_23__N_1310_adj_7491[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[21]), 
          .B1(op_i_23__N_1310_adj_7491[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32333), .COUT(n32334), .S0(op_i_23__N_1130_adj_7492[20]), 
          .S1(op_i_23__N_1130_adj_7492[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_22.INJECT1_1 = "NO";
    LUT4 i15661_3_lut (.A(\result_r[26] [7]), .B(\result_r[27] [7]), .C(y_1_delay[0]), 
         .Z(n34045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15661_3_lut.init = 16'hcaca;
    LUT4 i8433_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[279])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8433_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1045_add_4_6 (.A0(shift_2_dout_i[4]), .B0(shift_2_dout_r[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[5]), .B1(shift_2_dout_r[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32012), .COUT(n32013), .S0(n114), 
          .S1(n111));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_20 (.A0(op_r_23__N_1268_adj_7486[18]), .B0(op_i_23__N_1310_adj_7491[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[19]), 
          .B1(op_i_23__N_1310_adj_7491[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32332), .COUT(n32333), .S0(op_i_23__N_1130_adj_7492[18]), 
          .S1(op_i_23__N_1130_adj_7492[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_4 (.A0(shift_2_dout_i[2]), .B0(shift_2_dout_r[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[3]), .B1(shift_2_dout_r[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32011), .COUT(n32012), .S0(n120), 
          .S1(n117));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1045_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1045_add_4_2 (.A0(shift_2_dout_i[0]), .B0(shift_2_dout_r[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[1]), .B1(shift_2_dout_r[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32011), .S1(n123));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1045_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1045_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1045_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1045_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_18 (.A0(op_r_23__N_1268_adj_7486[16]), .B0(op_i_23__N_1310_adj_7491[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[17]), 
          .B1(op_i_23__N_1310_adj_7491[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32331), .COUT(n32332), .S0(op_i_23__N_1130_adj_7492[16]), 
          .S1(op_i_23__N_1130_adj_7492[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_18.INJECT1_1 = "NO";
    LUT4 i8425_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[280])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8425_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15528_3_lut (.A(\result_r[8] [11]), .B(\result_r[9] [11]), .C(y_1_delay[0]), 
         .Z(n33912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15528_3_lut.init = 16'hcaca;
    CCU2C _add_1_1081_add_4_16 (.A0(op_r_23__N_1268_adj_7486[14]), .B0(op_i_23__N_1310_adj_7491[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[15]), 
          .B1(op_i_23__N_1310_adj_7491[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32330), .COUT(n32331));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_25 (.A0(shift_2_dout_i[22]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[30]), .D0(n34576), .A1(shift_2_dout_i[23]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[31]), .D1(n34575), 
          .CIN(n32008), .S0(op_i_23__N_1154_adj_7426[22]), .S1(op_i_23__N_1154_adj_7426[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_23 (.A0(shift_2_dout_i[20]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[28]), .D0(n34580), .A1(shift_2_dout_i[21]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[29]), .D1(n34579), 
          .CIN(n32007), .COUT(n32008), .S0(op_i_23__N_1154_adj_7426[20]), 
          .S1(op_i_23__N_1154_adj_7426[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_14 (.A0(op_r_23__N_1268_adj_7486[12]), .B0(op_i_23__N_1310_adj_7491[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[13]), 
          .B1(op_i_23__N_1310_adj_7491[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32329), .COUT(n32330));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_14.INJECT1_1 = "NO";
    LUT4 i15527_3_lut (.A(\result_r[6] [11]), .B(\result_r[7] [11]), .C(y_1_delay[0]), 
         .Z(n33911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15527_3_lut.init = 16'hcaca;
    CCU2C _add_1_1056_add_4_21 (.A0(shift_2_dout_i[18]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[26]), .D0(n34584), .A1(shift_2_dout_i[19]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[27]), .D1(n34583), 
          .CIN(n32006), .COUT(n32007), .S0(op_i_23__N_1154_adj_7426[18]), 
          .S1(op_i_23__N_1154_adj_7426[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_19 (.A0(shift_2_dout_i[16]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[24]), .D0(n34588), .A1(shift_2_dout_i[17]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[25]), .D1(n34587), 
          .CIN(n32005), .COUT(n32006), .S0(op_i_23__N_1154_adj_7426[16]), 
          .S1(op_i_23__N_1154_adj_7426[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_12 (.A0(op_r_23__N_1268_adj_7486[10]), .B0(op_i_23__N_1310_adj_7491[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[11]), 
          .B1(op_i_23__N_1310_adj_7491[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32328), .COUT(n32329));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_17 (.A0(shift_2_dout_i[14]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[22]), .D0(n34596), .A1(shift_2_dout_i[15]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[23]), .D1(n34595), 
          .CIN(n32004), .COUT(n32005), .S0(op_i_23__N_1154_adj_7426[14]), 
          .S1(op_i_23__N_1154_adj_7426[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_15 (.A0(shift_2_dout_i[12]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[20]), .D0(n34604), .A1(shift_2_dout_i[13]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[21]), .D1(n34603), 
          .CIN(n32003), .COUT(n32004), .S0(op_i_23__N_1154_adj_7426[12]), 
          .S1(op_i_23__N_1154_adj_7426[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_10 (.A0(op_r_23__N_1268_adj_7486[8]), .B0(op_i_23__N_1310_adj_7491[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[9]), 
          .B1(op_i_23__N_1310_adj_7491[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32327), .COUT(n32328));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_10.INJECT1_1 = "NO";
    LUT4 i15526_3_lut (.A(\result_r[4] [11]), .B(\result_r[5] [11]), .C(y_1_delay[0]), 
         .Z(n33910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15526_3_lut.init = 16'hcaca;
    CCU2C _add_1_1056_add_4_13 (.A0(shift_2_dout_i[10]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[18]), .D0(n34612), .A1(shift_2_dout_i[11]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[19]), .D1(n34611), 
          .CIN(n32002), .COUT(n32003), .S0(op_i_23__N_1154_adj_7426[10]), 
          .S1(op_i_23__N_1154_adj_7426[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_11 (.A0(shift_2_dout_i[8]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[16]), .D0(n34624), .A1(shift_2_dout_i[9]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[17]), .D1(n34623), 
          .CIN(n32001), .COUT(n32002), .S0(op_i_23__N_1154_adj_7426[8]), 
          .S1(op_i_23__N_1154_adj_7426[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_8 (.A0(op_r_23__N_1268_adj_7486[6]), .B0(op_i_23__N_1310_adj_7491[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[7]), 
          .B1(op_i_23__N_1310_adj_7491[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32326), .COUT(n32327));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_9 (.A0(shift_2_dout_i[6]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[14]), .D0(n34636), .A1(shift_2_dout_i[7]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[15]), .D1(n34635), 
          .CIN(n32000), .COUT(n32001), .S0(op_i_23__N_1154_adj_7426[6]), 
          .S1(op_i_23__N_1154_adj_7426[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_7 (.A0(shift_2_dout_i[4]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[12]), .D0(n34646), .A1(shift_2_dout_i[5]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[13]), .D1(n34645), 
          .CIN(n31999), .COUT(n32000), .S0(op_i_23__N_1154_adj_7426[4]), 
          .S1(op_i_23__N_1154_adj_7426[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_6 (.A0(op_r_23__N_1268_adj_7486[4]), .B0(op_i_23__N_1310_adj_7491[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[5]), 
          .B1(op_i_23__N_1310_adj_7491[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32325), .COUT(n32326));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_6.INJECT1_1 = "NO";
    LUT4 i8417_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[281])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8417_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1056_add_4_5 (.A0(shift_2_dout_i[2]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[10]), .D0(n34656), .A1(shift_2_dout_i[3]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[11]), .D1(n34655), 
          .CIN(n31998), .COUT(n31999), .S0(op_i_23__N_1154_adj_7426[2]), 
          .S1(op_i_23__N_1154_adj_7426[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_4 (.A0(op_r_23__N_1268_adj_7486[2]), .B0(op_i_23__N_1310_adj_7491[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[3]), 
          .B1(op_i_23__N_1310_adj_7491[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32324), .COUT(n32325));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1081_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_3 (.A0(shift_2_dout_i[0]), .B0(state_1__N_5843[1]), 
          .C0(op_i_23__N_1130_adj_7436[8]), .D0(n34668), .A1(shift_2_dout_i[1]), 
          .B1(state_1__N_5843[1]), .C1(op_i_23__N_1130_adj_7436[9]), .D1(n34667), 
          .CIN(n31997), .COUT(n31998), .S0(op_i_23__N_1154_adj_7426[0]), 
          .S1(op_i_23__N_1154_adj_7426[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1056_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1056_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1056_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n34800), .B1(n34801), .C1(count_adj_7456[1]), 
          .D1(s_count_adj_7458[1]), .COUT(n31997));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1056_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1056_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1056_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1056_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1081_add_4_2 (.A0(op_r_23__N_1268_adj_7486[0]), .B0(op_i_23__N_1310_adj_7491[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[1]), 
          .B1(op_i_23__N_1310_adj_7491[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32324));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1081_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1081_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1081_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1081_add_4_2.INJECT1_1 = "NO";
    LUT4 i15660_3_lut (.A(\result_r[24] [7]), .B(\result_r[25] [7]), .C(y_1_delay[0]), 
         .Z(n34044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15660_3_lut.init = 16'hcaca;
    PFUMX i15792 (.BLUT(n34164), .ALUT(n34165), .C0(y_1_delay[1]), .Z(n34176));
    CCU2C _add_1_1067_add_4_32 (.A0(op_r_23__N_1268_adj_7430[30]), .B0(op_r_23__N_1226_adj_7432[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[31]), 
          .B1(op_r_23__N_1226_adj_7432[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31992), .S0(op_r_23__N_1082_adj_7433[30]), .S1(op_r_23__N_1082_adj_7433[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_26 (.A0(n8697), .B0(n65_adj_6358), .C0(GND_net), 
          .D0(VCC_net), .A1(n8696), .B1(n65_adj_6358), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32322), .S0(op_i_23__N_1310_adj_7329[30]), 
          .S1(op_i_23__N_1310_adj_7329[31]));
    defparam _add_1_1017_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_30 (.A0(op_r_23__N_1268_adj_7430[28]), .B0(op_r_23__N_1226_adj_7432[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[29]), 
          .B1(op_r_23__N_1226_adj_7432[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31991), .COUT(n31992), .S0(op_r_23__N_1082_adj_7433[28]), 
          .S1(op_r_23__N_1082_adj_7433[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_28 (.A0(op_r_23__N_1268_adj_7430[26]), .B0(op_r_23__N_1226_adj_7432[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[27]), 
          .B1(op_r_23__N_1226_adj_7432[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31990), .COUT(n31991), .S0(op_r_23__N_1082_adj_7433[26]), 
          .S1(op_r_23__N_1082_adj_7433[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_24 (.A0(n8699), .B0(n67), .C0(GND_net), .D0(VCC_net), 
          .A1(n8698), .B1(n66), .C1(GND_net), .D1(VCC_net), .CIN(n32321), 
          .COUT(n32322), .S0(op_i_23__N_1310_adj_7329[28]), .S1(op_i_23__N_1310_adj_7329[29]));
    defparam _add_1_1017_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_24.INJECT1_1 = "NO";
    LUT4 i8409_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[282])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8409_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1067_add_4_26 (.A0(op_r_23__N_1268_adj_7430[24]), .B0(op_r_23__N_1226_adj_7432[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[25]), 
          .B1(op_r_23__N_1226_adj_7432[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31989), .COUT(n31990), .S0(op_r_23__N_1082_adj_7433[24]), 
          .S1(op_r_23__N_1082_adj_7433[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_24 (.A0(op_r_23__N_1268_adj_7430[22]), .B0(op_r_23__N_1226_adj_7432[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[23]), 
          .B1(op_r_23__N_1226_adj_7432[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31988), .COUT(n31989), .S0(op_r_23__N_1082_adj_7433[22]), 
          .S1(op_r_23__N_1082_adj_7433[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_22 (.A0(n8701), .B0(n69), .C0(GND_net), .D0(VCC_net), 
          .A1(n8700), .B1(n68), .C1(GND_net), .D1(VCC_net), .CIN(n32320), 
          .COUT(n32321), .S0(op_i_23__N_1310_adj_7329[26]), .S1(op_i_23__N_1310_adj_7329[27]));
    defparam _add_1_1017_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_22 (.A0(op_r_23__N_1268_adj_7430[20]), .B0(op_r_23__N_1226_adj_7432[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[21]), 
          .B1(op_r_23__N_1226_adj_7432[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31987), .COUT(n31988), .S0(op_r_23__N_1082_adj_7433[20]), 
          .S1(op_r_23__N_1082_adj_7433[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_20 (.A0(op_r_23__N_1268_adj_7430[18]), .B0(op_r_23__N_1226_adj_7432[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[19]), 
          .B1(op_r_23__N_1226_adj_7432[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31986), .COUT(n31987), .S0(op_r_23__N_1082_adj_7433[18]), 
          .S1(op_r_23__N_1082_adj_7433[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_20 (.A0(n8703), .B0(n71), .C0(GND_net), .D0(VCC_net), 
          .A1(n8702), .B1(n70), .C1(GND_net), .D1(VCC_net), .CIN(n32319), 
          .COUT(n32320), .S0(op_i_23__N_1310_adj_7329[24]), .S1(op_i_23__N_1310_adj_7329[25]));
    defparam _add_1_1017_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_18 (.A0(op_r_23__N_1268_adj_7430[16]), .B0(op_r_23__N_1226_adj_7432[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[17]), 
          .B1(op_r_23__N_1226_adj_7432[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31985), .COUT(n31986), .S0(op_r_23__N_1082_adj_7433[16]), 
          .S1(op_r_23__N_1082_adj_7433[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_16 (.A0(op_r_23__N_1268_adj_7430[14]), .B0(op_r_23__N_1226_adj_7432[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[15]), 
          .B1(op_r_23__N_1226_adj_7432[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31984), .COUT(n31985), .S0(op_r_23__N_1082_adj_7433[14]), 
          .S1(op_r_23__N_1082_adj_7433[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_18 (.A0(n8705), .B0(n73), .C0(GND_net), .D0(VCC_net), 
          .A1(n8704), .B1(n72), .C1(GND_net), .D1(VCC_net), .CIN(n32318), 
          .COUT(n32319), .S0(op_i_23__N_1310_adj_7329[22]), .S1(op_i_23__N_1310_adj_7329[23]));
    defparam _add_1_1017_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_14 (.A0(op_r_23__N_1268_adj_7430[12]), .B0(op_r_23__N_1226_adj_7432[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[13]), 
          .B1(op_r_23__N_1226_adj_7432[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31983), .COUT(n31984), .S0(op_r_23__N_1082_adj_7433[12]), 
          .S1(op_r_23__N_1082_adj_7433[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_12 (.A0(op_r_23__N_1268_adj_7430[10]), .B0(op_r_23__N_1226_adj_7432[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[11]), 
          .B1(op_r_23__N_1226_adj_7432[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31982), .COUT(n31983), .S0(op_r_23__N_1082_adj_7433[10]), 
          .S1(op_r_23__N_1082_adj_7433[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_16 (.A0(n8707), .B0(n75), .C0(GND_net), .D0(VCC_net), 
          .A1(n8706), .B1(n74), .C1(GND_net), .D1(VCC_net), .CIN(n32317), 
          .COUT(n32318), .S0(op_i_23__N_1310_adj_7329[20]), .S1(op_i_23__N_1310_adj_7329[21]));
    defparam _add_1_1017_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_16.INJECT1_1 = "NO";
    LUT4 i8401_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[283])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8401_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8393_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[284])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8393_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1067_add_4_10 (.A0(op_r_23__N_1268_adj_7430[8]), .B0(op_r_23__N_1226_adj_7432[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[9]), 
          .B1(op_r_23__N_1226_adj_7432[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31981), .COUT(n31982), .S0(op_r_23__N_1082_adj_7433[8]), 
          .S1(op_r_23__N_1082_adj_7433[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_14 (.A0(n8709), .B0(n77), .C0(GND_net), .D0(VCC_net), 
          .A1(n8708), .B1(n76), .C1(GND_net), .D1(VCC_net), .CIN(n32316), 
          .COUT(n32317), .S0(op_i_23__N_1310_adj_7329[18]), .S1(op_i_23__N_1310_adj_7329[19]));
    defparam _add_1_1017_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_8 (.A0(op_r_23__N_1268_adj_7430[6]), .B0(op_r_23__N_1226_adj_7432[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[7]), 
          .B1(op_r_23__N_1226_adj_7432[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31980), .COUT(n31981));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_6 (.A0(op_r_23__N_1268_adj_7430[4]), .B0(op_r_23__N_1226_adj_7432[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[5]), 
          .B1(op_r_23__N_1226_adj_7432[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31979), .COUT(n31980));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_12 (.A0(n8711), .B0(n79), .C0(GND_net), .D0(VCC_net), 
          .A1(n8710), .B1(n78), .C1(GND_net), .D1(VCC_net), .CIN(n32315), 
          .COUT(n32316), .S0(op_i_23__N_1310_adj_7329[16]), .S1(op_i_23__N_1310_adj_7329[17]));
    defparam _add_1_1017_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_12.INJECT1_1 = "NO";
    LUT4 i8385_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[285])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8385_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1067_add_4_4 (.A0(op_r_23__N_1268_adj_7430[2]), .B0(op_r_23__N_1226_adj_7432[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[3]), 
          .B1(op_r_23__N_1226_adj_7432[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31978), .COUT(n31979));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1067_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_2 (.A0(op_r_23__N_1268_adj_7430[0]), .B0(op_r_23__N_1226_adj_7432[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[1]), 
          .B1(op_r_23__N_1226_adj_7432[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n31978));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1067_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1067_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1067_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_10 (.A0(n8713), .B0(n81), .C0(GND_net), .D0(VCC_net), 
          .A1(n8712), .B1(n80), .C1(GND_net), .D1(VCC_net), .CIN(n32314), 
          .COUT(n32315), .S0(op_i_23__N_1310_adj_7329[14]), .S1(op_i_23__N_1310_adj_7329[15]));
    defparam _add_1_1017_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1078_add_4_25 (.A0(shift_1_dout_i[23]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[23]), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n31977), .S0(op_i_23__N_1154_adj_7482[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_25.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_25.INIT1 = 16'h0000;
    defparam _add_1_1078_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1078_add_4_23 (.A0(shift_1_dout_i[21]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[21]), .A1(shift_1_dout_i[22]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[22]), .CIN(n31976), 
          .COUT(n31977), .S0(op_i_23__N_1154_adj_7482[21]), .S1(op_i_23__N_1154_adj_7482[22]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_23.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_23.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_8 (.A0(n8715), .B0(n83), .C0(GND_net), .D0(VCC_net), 
          .A1(n8714), .B1(n82), .C1(GND_net), .D1(VCC_net), .CIN(n32313), 
          .COUT(n32314), .S0(op_i_23__N_1310_adj_7329[12]), .S1(op_i_23__N_1310_adj_7329[13]));
    defparam _add_1_1017_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_8.INJECT1_1 = "NO";
    LUT4 i15787_3_lut (.A(\result_r[30] [3]), .B(\result_r[31] [3]), .C(y_1_delay[0]), 
         .Z(n34171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15787_3_lut.init = 16'hcaca;
    CCU2C _add_1_1078_add_4_21 (.A0(shift_1_dout_i[19]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[19]), .A1(shift_1_dout_i[20]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[20]), .CIN(n31975), 
          .COUT(n31976), .S0(op_i_23__N_1154_adj_7482[19]), .S1(op_i_23__N_1154_adj_7482[20]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_21.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_21.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1078_add_4_19 (.A0(shift_1_dout_i[17]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[17]), .A1(shift_1_dout_i[18]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[18]), .CIN(n31974), 
          .COUT(n31975), .S0(op_i_23__N_1154_adj_7482[17]), .S1(op_i_23__N_1154_adj_7482[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_19.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_19.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_6 (.A0(n8717), .B0(n85), .C0(GND_net), .D0(VCC_net), 
          .A1(n8716), .B1(n84), .C1(GND_net), .D1(VCC_net), .CIN(n32312), 
          .COUT(n32313), .S0(op_i_23__N_1310_adj_7329[10]), .S1(op_i_23__N_1310_adj_7329[11]));
    defparam _add_1_1017_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1078_add_4_17 (.A0(shift_1_dout_i[15]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[15]), .A1(shift_1_dout_i[16]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[16]), .CIN(n31973), 
          .COUT(n31974), .S0(op_i_23__N_1154_adj_7482[15]), .S1(op_i_23__N_1154_adj_7482[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_17.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_17.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1078_add_4_15 (.A0(shift_1_dout_i[13]), .B0(n34769), .C0(n34839), 
          .D0(op_i_23__N_1154_adj_7426[13]), .A1(shift_1_dout_i[14]), .B1(n34769), 
          .C1(n34839), .D1(op_i_23__N_1154_adj_7426[14]), .CIN(n31972), 
          .COUT(n31973), .S0(op_i_23__N_1154_adj_7482[13]), .S1(op_i_23__N_1154_adj_7482[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_1078_add_4_15.INIT0 = 16'h56aa;
    defparam _add_1_1078_add_4_15.INIT1 = 16'h56aa;
    defparam _add_1_1078_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1078_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_4 (.A0(n8719), .B0(n87), .C0(GND_net), .D0(VCC_net), 
          .A1(n8718), .B1(n86), .C1(GND_net), .D1(VCC_net), .CIN(n32311), 
          .COUT(n32312), .S0(op_i_23__N_1310_adj_7329[8]), .S1(op_i_23__N_1310_adj_7329[9]));
    defparam _add_1_1017_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1017_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_4.INJECT1_1 = "NO";
    PFUMX i15293 (.BLUT(n33662), .ALUT(n33663), .C0(y_1_delay[1]), .Z(n33677));
    CCU2C _add_1_1017_add_4_2 (.A0(n8721), .B0(n89), .C0(GND_net), .D0(VCC_net), 
          .A1(n8720), .B1(n88), .C1(GND_net), .D1(VCC_net), .COUT(n32311), 
          .S1(op_i_23__N_1310_adj_7329[7]));
    defparam _add_1_1017_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1017_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1017_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_2.INJECT1_1 = "NO";
    LUT4 i15786_3_lut (.A(\result_r[28] [3]), .B(\result_r[29] [3]), .C(y_1_delay[0]), 
         .Z(n34170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15786_3_lut.init = 16'hcaca;
    PFUMX i15793 (.BLUT(n34166), .ALUT(n34167), .C0(y_1_delay[1]), .Z(n34177));
    CCU2C _add_1_1064_add_4_26 (.A0(n8953), .B0(n65), .C0(GND_net), .D0(VCC_net), 
          .A1(n8952), .B1(n65), .C1(GND_net), .D1(VCC_net), .CIN(n32308), 
          .S0(op_i_23__N_1310_adj_7435[30]), .S1(op_i_23__N_1310_adj_7435[31]));
    defparam _add_1_1064_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_24 (.A0(n8955), .B0(n67_adj_7239), .C0(GND_net), 
          .D0(VCC_net), .A1(n8954), .B1(n66_adj_7238), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32307), .COUT(n32308), .S0(op_i_23__N_1310_adj_7435[28]), 
          .S1(op_i_23__N_1310_adj_7435[29]));
    defparam _add_1_1064_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_24.INJECT1_1 = "NO";
    LUT4 i8377_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[286])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8377_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_1064_add_4_22 (.A0(n8957), .B0(n69_adj_7241), .C0(GND_net), 
          .D0(VCC_net), .A1(n8956), .B1(n68_adj_7240), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32306), .COUT(n32307), .S0(op_i_23__N_1310_adj_7435[26]), 
          .S1(op_i_23__N_1310_adj_7435[27]));
    defparam _add_1_1064_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_20 (.A0(n8959), .B0(n71_adj_7243), .C0(GND_net), 
          .D0(VCC_net), .A1(n8958), .B1(n70_adj_7242), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32305), .COUT(n32306), .S0(op_i_23__N_1310_adj_7435[24]), 
          .S1(op_i_23__N_1310_adj_7435[25]));
    defparam _add_1_1064_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_20.INJECT1_1 = "NO";
    CCU2C add_13626_25 (.A0(n7433), .B0(n34799), .C0(n34591), .D0(rom4_state[0]), 
          .A1(n7432), .B1(n34799), .C1(n34592), .D1(rom4_state[0]), 
          .CIN(n32464), .S0(dout_r_23__N_5203[22]), .S1(dout_r_23__N_5203[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_25.INIT0 = 16'ha9aa;
    defparam add_13626_25.INIT1 = 16'ha9aa;
    defparam add_13626_25.INJECT1_0 = "NO";
    defparam add_13626_25.INJECT1_1 = "NO";
    LUT4 i8369_3_lut_4_lut (.A(n30503), .B(n34707), .C(\result_r[14] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[287])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8369_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i4529_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[8]), .D(\result_i[15] [0]), 
         .Z(result_i_ns_0__15__N_517[256])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4529_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1064_add_4_18 (.A0(n8961), .B0(n73_adj_7245), .C0(GND_net), 
          .D0(VCC_net), .A1(n8960), .B1(n72_adj_7244), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32304), .COUT(n32305), .S0(op_i_23__N_1310_adj_7435[22]), 
          .S1(op_i_23__N_1310_adj_7435[23]));
    defparam _add_1_1064_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_18.INJECT1_1 = "NO";
    LUT4 i4521_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[9]), .D(\result_i[15] [1]), 
         .Z(result_i_ns_0__15__N_517[257])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4521_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1064_add_4_16 (.A0(n8963), .B0(n75_adj_7247), .C0(GND_net), 
          .D0(VCC_net), .A1(n8962), .B1(n74_adj_7246), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32303), .COUT(n32304), .S0(op_i_23__N_1310_adj_7435[20]), 
          .S1(op_i_23__N_1310_adj_7435[21]));
    defparam _add_1_1064_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_16.INJECT1_1 = "NO";
    CCU2C add_13626_23 (.A0(n7435), .B0(n34799), .C0(n34599), .D0(rom4_state[0]), 
          .A1(n7434), .B1(n34799), .C1(n34600), .D1(rom4_state[0]), 
          .CIN(n32463), .COUT(n32464), .S0(dout_r_23__N_5203[20]), .S1(dout_r_23__N_5203[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_23.INIT0 = 16'ha9aa;
    defparam add_13626_23.INIT1 = 16'ha9aa;
    defparam add_13626_23.INJECT1_0 = "NO";
    defparam add_13626_23.INJECT1_1 = "NO";
    LUT4 i4513_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[10]), .D(\result_i[15] [2]), 
         .Z(result_i_ns_0__15__N_517[258])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4513_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1064_add_4_14 (.A0(n8965), .B0(n77_adj_7249), .C0(GND_net), 
          .D0(VCC_net), .A1(n8964), .B1(n76_adj_7248), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32302), .COUT(n32303), .S0(op_i_23__N_1310_adj_7435[18]), 
          .S1(op_i_23__N_1310_adj_7435[19]));
    defparam _add_1_1064_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_12 (.A0(n8967), .B0(n79_adj_7251), .C0(GND_net), 
          .D0(VCC_net), .A1(n8966), .B1(n78_adj_7250), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32301), .COUT(n32302), .S0(op_i_23__N_1310_adj_7435[16]), 
          .S1(op_i_23__N_1310_adj_7435[17]));
    defparam _add_1_1064_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_12.INJECT1_1 = "NO";
    CCU2C add_13626_21 (.A0(n7437), .B0(n34799), .C0(n34607), .D0(rom4_state[0]), 
          .A1(n7436), .B1(n34799), .C1(n34608), .D1(rom4_state[0]), 
          .CIN(n32462), .COUT(n32463), .S0(dout_r_23__N_5203[18]), .S1(dout_r_23__N_5203[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_21.INIT0 = 16'ha9aa;
    defparam add_13626_21.INIT1 = 16'ha9aa;
    defparam add_13626_21.INJECT1_0 = "NO";
    defparam add_13626_21.INJECT1_1 = "NO";
    LUT4 i15785_3_lut (.A(\result_r[26] [3]), .B(\result_r[27] [3]), .C(y_1_delay[0]), 
         .Z(n34169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15785_3_lut.init = 16'hcaca;
    LUT4 i4505_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[11]), .D(\result_i[15] [3]), 
         .Z(result_i_ns_0__15__N_517[259])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4505_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1064_add_4_10 (.A0(n8969), .B0(n81_adj_7253), .C0(GND_net), 
          .D0(VCC_net), .A1(n8968), .B1(n80_adj_7252), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32300), .COUT(n32301), .S0(op_i_23__N_1310_adj_7435[14]), 
          .S1(op_i_23__N_1310_adj_7435[15]));
    defparam _add_1_1064_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_10.INJECT1_1 = "NO";
    LUT4 i4497_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[12]), .D(\result_i[15] [4]), 
         .Z(result_i_ns_0__15__N_517[260])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4497_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1064_add_4_8 (.A0(n8971), .B0(n83_adj_7255), .C0(GND_net), 
          .D0(VCC_net), .A1(n8970), .B1(n82_adj_7254), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32299), .COUT(n32300), .S0(op_i_23__N_1310_adj_7435[12]), 
          .S1(op_i_23__N_1310_adj_7435[13]));
    defparam _add_1_1064_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_8.INJECT1_1 = "NO";
    CCU2C add_13626_19 (.A0(n7439), .B0(n34799), .C0(n34619), .D0(rom4_state[0]), 
          .A1(n7438), .B1(n34799), .C1(n34620), .D1(rom4_state[0]), 
          .CIN(n32461), .COUT(n32462), .S0(dout_r_23__N_5203[16]), .S1(dout_r_23__N_5203[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_19.INIT0 = 16'ha9aa;
    defparam add_13626_19.INIT1 = 16'ha9aa;
    defparam add_13626_19.INJECT1_0 = "NO";
    defparam add_13626_19.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_6 (.A0(n8973), .B0(n85_adj_7257), .C0(GND_net), 
          .D0(VCC_net), .A1(n8972), .B1(n84_adj_7256), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32298), .COUT(n32299), .S0(op_i_23__N_1310_adj_7435[10]), 
          .S1(op_i_23__N_1310_adj_7435[11]));
    defparam _add_1_1064_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_4 (.A0(n8975), .B0(n87_adj_7259), .C0(GND_net), 
          .D0(VCC_net), .A1(n8974), .B1(n86_adj_7258), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32297), .COUT(n32298), .S0(op_i_23__N_1310_adj_7435[8]), 
          .S1(op_i_23__N_1310_adj_7435[9]));
    defparam _add_1_1064_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1064_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_4.INJECT1_1 = "NO";
    CCU2C add_13626_17 (.A0(n7441), .B0(n34799), .C0(n34631), .D0(rom4_state[0]), 
          .A1(n7440), .B1(n34799), .C1(n34632), .D1(rom4_state[0]), 
          .CIN(n32460), .COUT(n32461), .S0(dout_r_23__N_5203[14]), .S1(dout_r_23__N_5203[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_17.INIT0 = 16'ha9aa;
    defparam add_13626_17.INIT1 = 16'ha9aa;
    defparam add_13626_17.INJECT1_0 = "NO";
    defparam add_13626_17.INJECT1_1 = "NO";
    LUT4 i4489_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[13]), .D(\result_i[15] [5]), 
         .Z(result_i_ns_0__15__N_517[261])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4489_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1064_add_4_2 (.A0(n8977), .B0(n89_adj_7261), .C0(GND_net), 
          .D0(VCC_net), .A1(n8976), .B1(n88_adj_7260), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32297), .S1(op_i_23__N_1310_adj_7435[7]));
    defparam _add_1_1064_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1064_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1064_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_2.INJECT1_1 = "NO";
    CCU2C add_13626_15 (.A0(n7443), .B0(n34799), .C0(n34643), .D0(rom4_state[0]), 
          .A1(n7442), .B1(n34799), .C1(n34644), .D1(rom4_state[0]), 
          .CIN(n32459), .COUT(n32460), .S0(dout_r_23__N_5203[12]), .S1(dout_r_23__N_5203[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_15.INIT0 = 16'ha9aa;
    defparam add_13626_15.INIT1 = 16'ha9aa;
    defparam add_13626_15.INJECT1_0 = "NO";
    defparam add_13626_15.INJECT1_1 = "NO";
    LUT4 i6777_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[486])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6777_3_lut_4_lut.init = 16'hf2d0;
    CCU2C _add_1_998_add_4_26 (.A0(n8569), .B0(n65_adj_7237), .C0(GND_net), 
          .D0(VCC_net), .A1(n8568), .B1(n65_adj_7237), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32294), .S0(op_i_23__N_1310[30]), .S1(op_i_23__N_1310[31]));
    defparam _add_1_998_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_26.INJECT1_1 = "NO";
    PFUMX i15540 (.BLUT(n33908), .ALUT(n33909), .C0(y_1_delay[1]), .Z(n33924));
    LUT4 i15784_3_lut (.A(\result_r[24] [3]), .B(\result_r[25] [3]), .C(y_1_delay[0]), 
         .Z(n34168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15784_3_lut.init = 16'hcaca;
    CCU2C _add_1_998_add_4_24 (.A0(n8571), .B0(n67_adj_7235), .C0(GND_net), 
          .D0(VCC_net), .A1(n8570), .B1(n66_adj_7236), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32293), .COUT(n32294), .S0(op_i_23__N_1310[28]), 
          .S1(op_i_23__N_1310[29]));
    defparam _add_1_998_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_24.INJECT1_1 = "NO";
    CCU2C add_13626_13 (.A0(n7445), .B0(n34799), .C0(n34653), .D0(rom4_state[0]), 
          .A1(n7444), .B1(n34799), .C1(n34654), .D1(rom4_state[0]), 
          .CIN(n32458), .COUT(n32459), .S0(dout_r_23__N_5203[10]), .S1(dout_r_23__N_5203[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_13.INIT0 = 16'ha9aa;
    defparam add_13626_13.INIT1 = 16'ha9aa;
    defparam add_13626_13.INJECT1_0 = "NO";
    defparam add_13626_13.INJECT1_1 = "NO";
    LUT4 i4481_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[14]), .D(\result_i[15] [6]), 
         .Z(result_i_ns_0__15__N_517[262])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4481_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_998_add_4_22 (.A0(n8573), .B0(n69_adj_7233), .C0(GND_net), 
          .D0(VCC_net), .A1(n8572), .B1(n68_adj_7234), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32292), .COUT(n32293), .S0(op_i_23__N_1310[26]), 
          .S1(op_i_23__N_1310[27]));
    defparam _add_1_998_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_998_add_4_20 (.A0(n8575), .B0(n71_adj_7231), .C0(GND_net), 
          .D0(VCC_net), .A1(n8574), .B1(n70_adj_7232), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32291), .COUT(n32292), .S0(op_i_23__N_1310[24]), 
          .S1(op_i_23__N_1310[25]));
    defparam _add_1_998_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_20.INJECT1_1 = "NO";
    CCU2C add_13626_11 (.A0(n7447), .B0(n34799), .C0(n34663), .D0(rom4_state[0]), 
          .A1(n7446), .B1(n34799), .C1(n34664), .D1(rom4_state[0]), 
          .CIN(n32457), .COUT(n32458), .S0(dout_r_23__N_5203[8]), .S1(dout_r_23__N_5203[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_11.INIT0 = 16'ha9aa;
    defparam add_13626_11.INIT1 = 16'ha9aa;
    defparam add_13626_11.INJECT1_0 = "NO";
    defparam add_13626_11.INJECT1_1 = "NO";
    LUT4 i4473_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[15]), .D(\result_i[15] [7]), 
         .Z(result_i_ns_0__15__N_517[263])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4473_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_998_add_4_18 (.A0(n8577), .B0(n73_adj_7229), .C0(GND_net), 
          .D0(VCC_net), .A1(n8576), .B1(n72_adj_7230), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32290), .COUT(n32291), .S0(op_i_23__N_1310[22]), 
          .S1(op_i_23__N_1310[23]));
    defparam _add_1_998_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_18.INJECT1_1 = "NO";
    LUT4 i4465_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[16]), .D(\result_i[15] [8]), 
         .Z(result_i_ns_0__15__N_517[264])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4465_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_998_add_4_16 (.A0(n8579), .B0(n75_adj_7227), .C0(GND_net), 
          .D0(VCC_net), .A1(n8578), .B1(n74_adj_7228), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32289), .COUT(n32290), .S0(op_i_23__N_1310[20]), 
          .S1(op_i_23__N_1310[21]));
    defparam _add_1_998_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_16.INJECT1_1 = "NO";
    CCU2C add_13626_9 (.A0(n7449), .B0(n34799), .C0(n34687), .D0(rom4_state[0]), 
          .A1(n7448), .B1(n34799), .C1(n34688), .D1(rom4_state[0]), 
          .CIN(n32456), .COUT(n32457), .S0(dout_r_23__N_5203[6]), .S1(dout_r_23__N_5203[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_9.INIT0 = 16'ha9aa;
    defparam add_13626_9.INIT1 = 16'ha9aa;
    defparam add_13626_9.INJECT1_0 = "NO";
    defparam add_13626_9.INJECT1_1 = "NO";
    LUT4 i4457_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[17]), .D(\result_i[15] [9]), 
         .Z(result_i_ns_0__15__N_517[265])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4457_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15279_3_lut (.A(\result_i[6] [4]), .B(\result_i[7] [4]), .C(y_1_delay[0]), 
         .Z(n33663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15279_3_lut.init = 16'hcaca;
    CCU2C _add_1_998_add_4_14 (.A0(n8581), .B0(n77_adj_7225), .C0(GND_net), 
          .D0(VCC_net), .A1(n8580), .B1(n76_adj_7226), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32288), .COUT(n32289), .S0(op_i_23__N_1310[18]), 
          .S1(op_i_23__N_1310[19]));
    defparam _add_1_998_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_14.INJECT1_1 = "NO";
    LUT4 i4449_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[18]), .D(\result_i[15] [10]), 
         .Z(result_i_ns_0__15__N_517[266])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4449_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_998_add_4_12 (.A0(n8583), .B0(n79_adj_7223), .C0(GND_net), 
          .D0(VCC_net), .A1(n8582), .B1(n78_adj_7224), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32287), .COUT(n32288), .S0(op_i_23__N_1310[16]), 
          .S1(op_i_23__N_1310[17]));
    defparam _add_1_998_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_12.INJECT1_1 = "NO";
    CCU2C add_13626_7 (.A0(n7451), .B0(n34799), .C0(n34692), .D0(rom4_state[0]), 
          .A1(n7450), .B1(n34799), .C1(n34693), .D1(rom4_state[0]), 
          .CIN(n32455), .COUT(n32456), .S0(dout_r_23__N_5203[4]), .S1(dout_r_23__N_5203[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_7.INIT0 = 16'ha9aa;
    defparam add_13626_7.INIT1 = 16'ha9aa;
    defparam add_13626_7.INJECT1_0 = "NO";
    defparam add_13626_7.INJECT1_1 = "NO";
    LUT4 i4441_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[19]), .D(\result_i[15] [11]), 
         .Z(result_i_ns_0__15__N_517[267])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4441_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_998_add_4_10 (.A0(n8585), .B0(n81_adj_7221), .C0(GND_net), 
          .D0(VCC_net), .A1(n8584), .B1(n80_adj_7222), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32286), .COUT(n32287), .S0(op_i_23__N_1310[14]), 
          .S1(op_i_23__N_1310[15]));
    defparam _add_1_998_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_10.INJECT1_1 = "NO";
    LUT4 i4433_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[20]), .D(\result_i[15] [12]), 
         .Z(result_i_ns_0__15__N_517[268])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4433_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_998_add_4_8 (.A0(n8587), .B0(n83_adj_7219), .C0(GND_net), 
          .D0(VCC_net), .A1(n8586), .B1(n82_adj_7220), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32285), .COUT(n32286), .S0(op_i_23__N_1310[12]), 
          .S1(op_i_23__N_1310[13]));
    defparam _add_1_998_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_8.INJECT1_1 = "NO";
    CCU2C add_13626_5 (.A0(n7453), .B0(n34799), .C0(n34695), .D0(rom4_state[0]), 
          .A1(n7452), .B1(n34799), .C1(n34696), .D1(rom4_state[0]), 
          .CIN(n32454), .COUT(n32455), .S0(dout_r_23__N_5203[2]), .S1(dout_r_23__N_5203[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_5.INIT0 = 16'ha9aa;
    defparam add_13626_5.INIT1 = 16'ha9aa;
    defparam add_13626_5.INJECT1_0 = "NO";
    defparam add_13626_5.INJECT1_1 = "NO";
    LUT4 i4425_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[21]), .D(\result_i[15] [13]), 
         .Z(result_i_ns_0__15__N_517[269])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4425_3_lut_4_lut.init = 16'hfb40;
    PFUMX i15794 (.BLUT(n34168), .ALUT(n34169), .C0(y_1_delay[1]), .Z(n34178));
    CCU2C _add_1_998_add_4_6 (.A0(n8589), .B0(n85_adj_7217), .C0(GND_net), 
          .D0(VCC_net), .A1(n8588), .B1(n84_adj_7218), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32284), .COUT(n32285), .S0(op_i_23__N_1310[10]), 
          .S1(op_i_23__N_1310[11]));
    defparam _add_1_998_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_998_add_4_4 (.A0(n8591), .B0(n87_adj_7166), .C0(GND_net), 
          .D0(VCC_net), .A1(n8590), .B1(n86_adj_7216), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32283), .COUT(n32284), .S0(op_i_23__N_1310[8]), 
          .S1(op_i_23__N_1310[9]));
    defparam _add_1_998_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_998_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_4.INJECT1_1 = "NO";
    CCU2C add_13626_3 (.A0(n7455), .B0(n34799), .C0(n34699), .D0(rom4_state[0]), 
          .A1(n7454), .B1(n34799), .C1(n34700), .D1(rom4_state[0]), 
          .CIN(n32453), .COUT(n32454), .S0(dout_r_23__N_5203[0]), .S1(dout_r_23__N_5203[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_3.INIT0 = 16'ha9aa;
    defparam add_13626_3.INIT1 = 16'ha9aa;
    defparam add_13626_3.INJECT1_0 = "NO";
    defparam add_13626_3.INJECT1_1 = "NO";
    CCU2C _add_1_998_add_4_2 (.A0(n8593), .B0(n89_adj_7164), .C0(GND_net), 
          .D0(VCC_net), .A1(n8592), .B1(n88_adj_7165), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32283), .S1(op_i_23__N_1310[7]));
    defparam _add_1_998_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_998_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_998_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_998_add_4_2.INJECT1_1 = "NO";
    CCU2C add_13626_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n29826), .B1(n29827), .C1(n29828), .D1(rom4_state[0]), 
          .COUT(n32453));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13626_1.INIT0 = 16'h0000;
    defparam add_13626_1.INIT1 = 16'hd8ff;
    defparam add_13626_1.INJECT1_0 = "NO";
    defparam add_13626_1.INJECT1_1 = "NO";
    LUT4 i4417_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[22]), .D(\result_i[15] [14]), 
         .Z(result_i_ns_0__15__N_517[270])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4417_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_26 (.A0(n8825), .B0(n65_adj_6772), .C0(GND_net), 
          .D0(VCC_net), .A1(n8824), .B1(n65_adj_6772), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32280), .S0(op_i_23__N_1310_adj_7380[30]), 
          .S1(op_i_23__N_1310_adj_7380[31]));
    defparam _add_1_1039_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1039_add_4_24 (.A0(n8827), .B0(n67_adj_7269), .C0(GND_net), 
          .D0(VCC_net), .A1(n8826), .B1(n66_adj_7268), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32279), .COUT(n32280), .S0(op_i_23__N_1310_adj_7380[28]), 
          .S1(op_i_23__N_1310_adj_7380[29]));
    defparam _add_1_1039_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_24.INJECT1_1 = "NO";
    LUT4 i15525_3_lut (.A(\result_r[2] [11]), .B(\result_r[3] [11]), .C(y_1_delay[0]), 
         .Z(n33909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15525_3_lut.init = 16'hcaca;
    CCU2C _add_1_1039_add_4_22 (.A0(n8829), .B0(n69_adj_7271), .C0(GND_net), 
          .D0(VCC_net), .A1(n8828), .B1(n68_adj_7270), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32278), .COUT(n32279), .S0(op_i_23__N_1310_adj_7380[26]), 
          .S1(op_i_23__N_1310_adj_7380[27]));
    defparam _add_1_1039_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1039_add_4_20 (.A0(n8831), .B0(n71_adj_7273), .C0(GND_net), 
          .D0(VCC_net), .A1(n8830), .B1(n70_adj_7272), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32277), .COUT(n32278), .S0(op_i_23__N_1310_adj_7380[24]), 
          .S1(op_i_23__N_1310_adj_7380[25]));
    defparam _add_1_1039_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_20.INJECT1_1 = "NO";
    LUT4 i4409_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_i[23]), .D(\result_i[15] [15]), 
         .Z(result_i_ns_0__15__N_517[271])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4409_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_18 (.A0(n8833), .B0(n73_adj_7275), .C0(GND_net), 
          .D0(VCC_net), .A1(n8832), .B1(n72_adj_7274), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32276), .COUT(n32277), .S0(op_i_23__N_1310_adj_7380[22]), 
          .S1(op_i_23__N_1310_adj_7380[23]));
    defparam _add_1_1039_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_18.INJECT1_1 = "NO";
    LUT4 i8617_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[8]), .D(\result_r[15] [0]), 
         .Z(result_r_ns_0__15__N_3[256])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8617_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8609_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[9]), .D(\result_r[15] [1]), 
         .Z(result_r_ns_0__15__N_3[257])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8609_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_16 (.A0(n8835), .B0(n75_adj_7277), .C0(GND_net), 
          .D0(VCC_net), .A1(n8834), .B1(n74_adj_7276), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32275), .COUT(n32276), .S0(op_i_23__N_1310_adj_7380[20]), 
          .S1(op_i_23__N_1310_adj_7380[21]));
    defparam _add_1_1039_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_16.INJECT1_1 = "NO";
    CCU2C add_13627_25 (.A0(n7592), .B0(n34799), .C0(n34590), .D0(rom4_state[0]), 
          .A1(n7591), .B1(n34799), .C1(n34589), .D1(rom4_state[0]), 
          .CIN(n32448), .S0(dout_i_23__N_5395[22]), .S1(dout_i_23__N_5395[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_25.INIT0 = 16'ha9aa;
    defparam add_13627_25.INIT1 = 16'ha9aa;
    defparam add_13627_25.INJECT1_0 = "NO";
    defparam add_13627_25.INJECT1_1 = "NO";
    LUT4 i8601_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[10]), .D(\result_r[15] [2]), 
         .Z(result_r_ns_0__15__N_3[258])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8601_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8593_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[11]), .D(\result_r[15] [3]), 
         .Z(result_r_ns_0__15__N_3[259])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8593_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_14 (.A0(n8837), .B0(n77_adj_7279), .C0(GND_net), 
          .D0(VCC_net), .A1(n8836), .B1(n76_adj_7278), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32274), .COUT(n32275), .S0(op_i_23__N_1310_adj_7380[18]), 
          .S1(op_i_23__N_1310_adj_7380[19]));
    defparam _add_1_1039_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_14.INJECT1_1 = "NO";
    LUT4 i8585_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[12]), .D(\result_r[15] [4]), 
         .Z(result_r_ns_0__15__N_3[260])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8585_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8577_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[13]), .D(\result_r[15] [5]), 
         .Z(result_r_ns_0__15__N_3[261])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8577_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_12 (.A0(n8839), .B0(n79_adj_7281), .C0(GND_net), 
          .D0(VCC_net), .A1(n8838), .B1(n78_adj_7280), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32273), .COUT(n32274), .S0(op_i_23__N_1310_adj_7380[16]), 
          .S1(op_i_23__N_1310_adj_7380[17]));
    defparam _add_1_1039_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_12.INJECT1_1 = "NO";
    CCU2C add_13627_23 (.A0(n7594), .B0(n34799), .C0(n34598), .D0(rom4_state[0]), 
          .A1(n7593), .B1(n34799), .C1(n34597), .D1(rom4_state[0]), 
          .CIN(n32447), .COUT(n32448), .S0(dout_i_23__N_5395[20]), .S1(dout_i_23__N_5395[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_23.INIT0 = 16'ha9aa;
    defparam add_13627_23.INIT1 = 16'ha9aa;
    defparam add_13627_23.INJECT1_0 = "NO";
    defparam add_13627_23.INJECT1_1 = "NO";
    PFUMX i15795 (.BLUT(n34170), .ALUT(n34171), .C0(y_1_delay[1]), .Z(n34179));
    LUT4 i15524_3_lut (.A(\result_r[0] [11]), .B(\result_r[1] [11]), .C(y_1_delay[0]), 
         .Z(n33908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15524_3_lut.init = 16'hcaca;
    CCU2C _add_1_1039_add_4_10 (.A0(n8841), .B0(n81_adj_7283), .C0(GND_net), 
          .D0(VCC_net), .A1(n8840), .B1(n80_adj_7282), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32272), .COUT(n32273), .S0(op_i_23__N_1310_adj_7380[14]), 
          .S1(op_i_23__N_1310_adj_7380[15]));
    defparam _add_1_1039_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_10.INJECT1_1 = "NO";
    PFUMX i15670 (.BLUT(n34044), .ALUT(n34045), .C0(y_1_delay[1]), .Z(n34054));
    CCU2C _add_1_1039_add_4_8 (.A0(n8843), .B0(n83_adj_7285), .C0(GND_net), 
          .D0(VCC_net), .A1(n8842), .B1(n82_adj_7284), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32271), .COUT(n32272), .S0(op_i_23__N_1310_adj_7380[12]), 
          .S1(op_i_23__N_1310_adj_7380[13]));
    defparam _add_1_1039_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_8.INJECT1_1 = "NO";
    CCU2C add_13627_21 (.A0(n7596), .B0(n34799), .C0(n34605), .D0(rom4_state[0]), 
          .A1(n7595), .B1(n34799), .C1(n34606), .D1(rom4_state[0]), 
          .CIN(n32446), .COUT(n32447), .S0(dout_i_23__N_5395[18]), .S1(dout_i_23__N_5395[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_21.INIT0 = 16'ha9aa;
    defparam add_13627_21.INIT1 = 16'ha9aa;
    defparam add_13627_21.INJECT1_0 = "NO";
    defparam add_13627_21.INJECT1_1 = "NO";
    CCU2C _add_1_1039_add_4_6 (.A0(n8845), .B0(n85_adj_7287), .C0(GND_net), 
          .D0(VCC_net), .A1(n8844), .B1(n84_adj_7286), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32270), .COUT(n32271), .S0(op_i_23__N_1310_adj_7380[10]), 
          .S1(op_i_23__N_1310_adj_7380[11]));
    defparam _add_1_1039_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_6.INJECT1_1 = "NO";
    LUT4 i8569_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[14]), .D(\result_r[15] [6]), 
         .Z(result_r_ns_0__15__N_3[262])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8569_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_4 (.A0(n8847), .B0(n87_adj_7289), .C0(GND_net), 
          .D0(VCC_net), .A1(n8846), .B1(n86_adj_7288), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32269), .COUT(n32270), .S0(op_i_23__N_1310_adj_7380[8]), 
          .S1(op_i_23__N_1310_adj_7380[9]));
    defparam _add_1_1039_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1039_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_4.INJECT1_1 = "NO";
    CCU2C add_13627_19 (.A0(n7598), .B0(n34799), .C0(n34613), .D0(rom4_state[0]), 
          .A1(n7597), .B1(n34799), .C1(n34614), .D1(rom4_state[0]), 
          .CIN(n32445), .COUT(n32446), .S0(dout_i_23__N_5395[16]), .S1(dout_i_23__N_5395[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_19.INIT0 = 16'ha9aa;
    defparam add_13627_19.INIT1 = 16'ha9aa;
    defparam add_13627_19.INJECT1_0 = "NO";
    defparam add_13627_19.INJECT1_1 = "NO";
    LUT4 i8561_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[15]), .D(\result_r[15] [7]), 
         .Z(result_r_ns_0__15__N_3[263])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8561_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8553_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[16]), .D(\result_r[15] [8]), 
         .Z(result_r_ns_0__15__N_3[264])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8553_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1039_add_4_2 (.A0(n8849), .B0(n89_adj_7291), .C0(GND_net), 
          .D0(VCC_net), .A1(n8848), .B1(n88_adj_7290), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32269), .S1(op_i_23__N_1310_adj_7380[7]));
    defparam _add_1_1039_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1039_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1039_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1039_add_4_2.INJECT1_1 = "NO";
    LUT4 i8545_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[17]), .D(\result_r[15] [9]), 
         .Z(result_r_ns_0__15__N_3[265])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8545_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8537_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[18]), .D(\result_r[15] [10]), 
         .Z(result_r_ns_0__15__N_3[266])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8537_3_lut_4_lut.init = 16'hfb40;
    CCU2C add_13627_17 (.A0(n7600), .B0(n34799), .C0(n34625), .D0(rom4_state[0]), 
          .A1(n7599), .B1(n34799), .C1(n34626), .D1(rom4_state[0]), 
          .CIN(n32444), .COUT(n32445), .S0(dout_i_23__N_5395[14]), .S1(dout_i_23__N_5395[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_17.INIT0 = 16'ha9aa;
    defparam add_13627_17.INIT1 = 16'ha9aa;
    defparam add_13627_17.INJECT1_0 = "NO";
    defparam add_13627_17.INJECT1_1 = "NO";
    LUT4 i15278_3_lut (.A(\result_i[4] [4]), .B(\result_i[5] [4]), .C(y_1_delay[0]), 
         .Z(n33662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15278_3_lut.init = 16'hcaca;
    LUT4 i8529_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[19]), .D(\result_r[15] [11]), 
         .Z(result_r_ns_0__15__N_3[267])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8529_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_32 (.A0(op_r_23__N_1268_adj_7486[30]), .B0(op_r_23__N_1226_adj_7488[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[31]), 
          .B1(op_r_23__N_1226_adj_7488[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32266), .S0(op_r_23__N_1082_adj_7489[30]), .S1(op_r_23__N_1082_adj_7489[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_32.INJECT1_1 = "NO";
    LUT4 i8521_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[20]), .D(\result_r[15] [12]), 
         .Z(result_r_ns_0__15__N_3[268])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8521_3_lut_4_lut.init = 16'hfb40;
    PFUMX i15541 (.BLUT(n33910), .ALUT(n33911), .C0(y_1_delay[1]), .Z(n33925));
    CCU2C _add_1_1089_add_4_30 (.A0(op_r_23__N_1268_adj_7486[28]), .B0(op_r_23__N_1226_adj_7488[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[29]), 
          .B1(op_r_23__N_1226_adj_7488[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32265), .COUT(n32266), .S0(op_r_23__N_1082_adj_7489[28]), 
          .S1(op_r_23__N_1082_adj_7489[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_30.INJECT1_1 = "NO";
    CCU2C add_13627_15 (.A0(n7602), .B0(n34799), .C0(n34637), .D0(rom4_state[0]), 
          .A1(n7601), .B1(n34799), .C1(n34638), .D1(rom4_state[0]), 
          .CIN(n32443), .COUT(n32444), .S0(dout_i_23__N_5395[12]), .S1(dout_i_23__N_5395[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_15.INIT0 = 16'ha9aa;
    defparam add_13627_15.INIT1 = 16'ha9aa;
    defparam add_13627_15.INJECT1_0 = "NO";
    defparam add_13627_15.INJECT1_1 = "NO";
    LUT4 i8513_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[21]), .D(\result_r[15] [13]), 
         .Z(result_r_ns_0__15__N_3[269])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8513_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_28 (.A0(op_r_23__N_1268_adj_7486[26]), .B0(op_r_23__N_1226_adj_7488[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[27]), 
          .B1(op_r_23__N_1226_adj_7488[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32264), .COUT(n32265), .S0(op_r_23__N_1082_adj_7489[26]), 
          .S1(op_r_23__N_1082_adj_7489[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1089_add_4_26 (.A0(op_r_23__N_1268_adj_7486[24]), .B0(op_r_23__N_1226_adj_7488[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[25]), 
          .B1(op_r_23__N_1226_adj_7488[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32263), .COUT(n32264), .S0(op_r_23__N_1082_adj_7489[24]), 
          .S1(op_r_23__N_1082_adj_7489[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_26.INJECT1_1 = "NO";
    CCU2C add_13627_13 (.A0(n7604), .B0(n34799), .C0(n34647), .D0(rom4_state[0]), 
          .A1(n7603), .B1(n34799), .C1(n34648), .D1(rom4_state[0]), 
          .CIN(n32442), .COUT(n32443), .S0(dout_i_23__N_5395[10]), .S1(dout_i_23__N_5395[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_13.INIT0 = 16'ha9aa;
    defparam add_13627_13.INIT1 = 16'ha9aa;
    defparam add_13627_13.INJECT1_0 = "NO";
    defparam add_13627_13.INJECT1_1 = "NO";
    LUT4 i8505_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[22]), .D(\result_r[15] [14]), 
         .Z(result_r_ns_0__15__N_3[270])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8505_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_24 (.A0(op_r_23__N_1268_adj_7486[22]), .B0(op_r_23__N_1226_adj_7488[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[23]), 
          .B1(op_r_23__N_1226_adj_7488[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32262), .COUT(n32263), .S0(op_r_23__N_1082_adj_7489[22]), 
          .S1(op_r_23__N_1082_adj_7489[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_24.INJECT1_1 = "NO";
    LUT4 i8497_3_lut_4_lut (.A(n34720), .B(n34708), .C(out_r[23]), .D(\result_r[15] [15]), 
         .Z(result_r_ns_0__15__N_3[271])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8497_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_22 (.A0(op_r_23__N_1268_adj_7486[20]), .B0(op_r_23__N_1226_adj_7488[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[21]), 
          .B1(op_r_23__N_1226_adj_7488[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32261), .COUT(n32262), .S0(op_r_23__N_1082_adj_7489[20]), 
          .S1(op_r_23__N_1082_adj_7489[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_22.INJECT1_1 = "NO";
    CCU2C add_13627_11 (.A0(n7606), .B0(n34799), .C0(n34657), .D0(rom4_state[0]), 
          .A1(n7605), .B1(n34799), .C1(n34658), .D1(rom4_state[0]), 
          .CIN(n32441), .COUT(n32442), .S0(dout_i_23__N_5395[8]), .S1(dout_i_23__N_5395[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_11.INIT0 = 16'ha9aa;
    defparam add_13627_11.INIT1 = 16'ha9aa;
    defparam add_13627_11.INJECT1_0 = "NO";
    defparam add_13627_11.INJECT1_1 = "NO";
    LUT4 i15783_3_lut (.A(\result_r[22] [3]), .B(\result_r[23] [3]), .C(y_1_delay[0]), 
         .Z(n34167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15783_3_lut.init = 16'hcaca;
    PFUMX i15542 (.BLUT(n33912), .ALUT(n33913), .C0(y_1_delay[1]), .Z(n33926));
    LUT4 i4657_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[8]), .D(\result_i[16] [0]), 
         .Z(result_i_ns_0__15__N_517[240])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4657_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_20 (.A0(op_r_23__N_1268_adj_7486[18]), .B0(op_r_23__N_1226_adj_7488[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[19]), 
          .B1(op_r_23__N_1226_adj_7488[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32260), .COUT(n32261), .S0(op_r_23__N_1082_adj_7489[18]), 
          .S1(op_r_23__N_1082_adj_7489[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_20.INJECT1_1 = "NO";
    LUT4 i4649_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[9]), .D(\result_i[16] [1]), 
         .Z(result_i_ns_0__15__N_517[241])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4649_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4641_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[10]), .D(\result_i[16] [2]), 
         .Z(result_i_ns_0__15__N_517[242])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4641_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_18 (.A0(op_r_23__N_1268_adj_7486[16]), .B0(op_r_23__N_1226_adj_7488[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[17]), 
          .B1(op_r_23__N_1226_adj_7488[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32259), .COUT(n32260), .S0(op_r_23__N_1082_adj_7489[16]), 
          .S1(op_r_23__N_1082_adj_7489[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_18.INJECT1_1 = "NO";
    CCU2C add_13627_9 (.A0(n7608), .B0(n34799), .C0(n34681), .D0(rom4_state[0]), 
          .A1(n7607), .B1(n34799), .C1(n34682), .D1(rom4_state[0]), 
          .CIN(n32440), .COUT(n32441), .S0(dout_i_23__N_5395[6]), .S1(dout_i_23__N_5395[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_9.INIT0 = 16'ha9aa;
    defparam add_13627_9.INIT1 = 16'ha9aa;
    defparam add_13627_9.INJECT1_0 = "NO";
    defparam add_13627_9.INJECT1_1 = "NO";
    LUT4 i4633_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[11]), .D(\result_i[16] [3]), 
         .Z(result_i_ns_0__15__N_517[243])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4633_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4625_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[12]), .D(\result_i[16] [4]), 
         .Z(result_i_ns_0__15__N_517[244])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4625_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_16 (.A0(op_r_23__N_1268_adj_7486[14]), .B0(op_r_23__N_1226_adj_7488[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[15]), 
          .B1(op_r_23__N_1226_adj_7488[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32258), .COUT(n32259));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1089_add_4_14 (.A0(op_r_23__N_1268_adj_7486[12]), .B0(op_r_23__N_1226_adj_7488[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[13]), 
          .B1(op_r_23__N_1226_adj_7488[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32257), .COUT(n32258));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_14.INJECT1_1 = "NO";
    CCU2C add_13627_7 (.A0(n7610), .B0(n34799), .C0(n34694), .D0(rom4_state[0]), 
          .A1(n7609), .B1(n34799), .C1(n34691), .D1(rom4_state[0]), 
          .CIN(n32439), .COUT(n32440), .S0(dout_i_23__N_5395[4]), .S1(dout_i_23__N_5395[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_7.INIT0 = 16'ha9aa;
    defparam add_13627_7.INIT1 = 16'ha9aa;
    defparam add_13627_7.INJECT1_0 = "NO";
    defparam add_13627_7.INJECT1_1 = "NO";
    LUT4 i4617_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[13]), .D(\result_i[16] [5]), 
         .Z(result_i_ns_0__15__N_517[245])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4617_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_12 (.A0(op_r_23__N_1268_adj_7486[10]), .B0(op_r_23__N_1226_adj_7488[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[11]), 
          .B1(op_r_23__N_1226_adj_7488[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32256), .COUT(n32257));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1089_add_4_10 (.A0(op_r_23__N_1268_adj_7486[8]), .B0(op_r_23__N_1226_adj_7488[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[9]), 
          .B1(op_r_23__N_1226_adj_7488[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32255), .COUT(n32256));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_10.INJECT1_1 = "NO";
    CCU2C add_13627_5 (.A0(n7612), .B0(n34799), .C0(n34697), .D0(rom4_state[0]), 
          .A1(n7611), .B1(n34799), .C1(n34698), .D1(rom4_state[0]), 
          .CIN(n32438), .COUT(n32439), .S0(dout_i_23__N_5395[2]), .S1(dout_i_23__N_5395[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_5.INIT0 = 16'ha9aa;
    defparam add_13627_5.INIT1 = 16'ha9aa;
    defparam add_13627_5.INJECT1_0 = "NO";
    defparam add_13627_5.INJECT1_1 = "NO";
    LUT4 i4609_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[14]), .D(\result_i[16] [6]), 
         .Z(result_i_ns_0__15__N_517[246])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4609_3_lut_4_lut.init = 16'hfb40;
    PFUMX i15819 (.BLUT(n34187), .ALUT(n34188), .C0(y_1_delay[1]), .Z(n34203));
    CCU2C _add_1_1089_add_4_8 (.A0(op_r_23__N_1268_adj_7486[6]), .B0(op_r_23__N_1226_adj_7488[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[7]), 
          .B1(op_r_23__N_1226_adj_7488[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32254), .COUT(n32255));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_8.INJECT1_1 = "NO";
    LUT4 i4601_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[15]), .D(\result_i[16] [7]), 
         .Z(result_i_ns_0__15__N_517[247])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4601_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15782_3_lut (.A(\result_r[20] [3]), .B(\result_r[21] [3]), .C(y_1_delay[0]), 
         .Z(n34166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15782_3_lut.init = 16'hcaca;
    CCU2C _add_1_1089_add_4_6 (.A0(op_r_23__N_1268_adj_7486[4]), .B0(op_r_23__N_1226_adj_7488[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[5]), 
          .B1(op_r_23__N_1226_adj_7488[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32253), .COUT(n32254));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_6.INJECT1_1 = "NO";
    CCU2C add_13627_3 (.A0(n7614), .B0(n34799), .C0(n34701), .D0(rom4_state[0]), 
          .A1(n7613), .B1(n34799), .C1(n34702), .D1(rom4_state[0]), 
          .CIN(n32437), .COUT(n32438), .S0(dout_i_23__N_5395[0]), .S1(dout_i_23__N_5395[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_3.INIT0 = 16'ha9aa;
    defparam add_13627_3.INIT1 = 16'ha9aa;
    defparam add_13627_3.INJECT1_0 = "NO";
    defparam add_13627_3.INJECT1_1 = "NO";
    LUT4 i4593_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[16]), .D(\result_i[16] [8]), 
         .Z(result_i_ns_0__15__N_517[248])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4593_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1089_add_4_4 (.A0(op_r_23__N_1268_adj_7486[2]), .B0(op_r_23__N_1226_adj_7488[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[3]), 
          .B1(op_r_23__N_1226_adj_7488[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32252), .COUT(n32253));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1089_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_4.INJECT1_1 = "NO";
    LUT4 i4585_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[17]), .D(\result_i[16] [9]), 
         .Z(result_i_ns_0__15__N_517[249])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4585_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15781_3_lut (.A(\result_r[18] [3]), .B(\result_r[19] [3]), .C(y_1_delay[0]), 
         .Z(n34165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15781_3_lut.init = 16'hcaca;
    CCU2C _add_1_1089_add_4_2 (.A0(op_r_23__N_1268_adj_7486[0]), .B0(op_r_23__N_1226_adj_7488[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7486[1]), 
          .B1(op_r_23__N_1226_adj_7488[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32252));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1089_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1089_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1089_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1089_add_4_2.INJECT1_1 = "NO";
    CCU2C add_13627_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n29826), .B1(n29827), .C1(n29828), .D1(rom4_state[0]), 
          .COUT(n32437));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13627_1.INIT0 = 16'h0000;
    defparam add_13627_1.INIT1 = 16'hd8ff;
    defparam add_13627_1.INJECT1_0 = "NO";
    defparam add_13627_1.INJECT1_1 = "NO";
    LUT4 i15780_3_lut (.A(\result_r[16] [3]), .B(\result_r[17] [3]), .C(y_1_delay[0]), 
         .Z(n34164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15780_3_lut.init = 16'hcaca;
    CCU2C _add_1_1101_add_4_26 (.A0(shift_1_dout_i[23]), .B0(shift_1_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[23]), .B1(shift_1_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32250), .S0(n12088), .S1(n12089));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1101_add_4_24 (.A0(shift_1_dout_i[21]), .B0(shift_1_dout_r[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[22]), .B1(shift_1_dout_r[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32249), .COUT(n32250), .S0(n12086), 
          .S1(n12087));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_24.INJECT1_1 = "NO";
    PFUMX i15820 (.BLUT(n34189), .ALUT(n34190), .C0(y_1_delay[1]), .Z(n34204));
    PFUMX i15671 (.BLUT(n34046), .ALUT(n34047), .C0(y_1_delay[1]), .Z(n34055));
    CCU2C _add_1_1101_add_4_22 (.A0(shift_1_dout_i[19]), .B0(shift_1_dout_r[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[20]), .B1(shift_1_dout_r[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32248), .COUT(n32249), .S0(n12084), 
          .S1(n12085));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1101_add_4_20 (.A0(shift_1_dout_i[17]), .B0(shift_1_dout_r[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[18]), .B1(shift_1_dout_r[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32247), .COUT(n32248), .S0(n12082), 
          .S1(n12083));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_20.INJECT1_1 = "NO";
    LUT4 i4577_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[18]), .D(\result_i[16] [10]), 
         .Z(result_i_ns_0__15__N_517[250])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4577_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_18 (.A0(shift_1_dout_i[15]), .B0(shift_1_dout_r[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[16]), .B1(shift_1_dout_r[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32246), .COUT(n32247), .S0(n12080), 
          .S1(n12081));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_18.INJECT1_1 = "NO";
    LUT4 i4569_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[19]), .D(\result_i[16] [11]), 
         .Z(result_i_ns_0__15__N_517[251])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4569_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_16 (.A0(shift_1_dout_i[13]), .B0(shift_1_dout_r[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[14]), .B1(shift_1_dout_r[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32245), .COUT(n32246), .S0(n12078), 
          .S1(n12079));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_16.INJECT1_1 = "NO";
    CCU2C add_13625_25 (.A0(n7486), .B0(n34794), .C0(n34617), .D0(rom8_state[0]), 
          .A1(n7485), .B1(n34794), .C1(n34618), .D1(rom8_state[0]), 
          .CIN(n32432), .S0(dout_i_23__N_4670[22]), .S1(dout_i_23__N_4670[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_25.INIT0 = 16'ha9aa;
    defparam add_13625_25.INIT1 = 16'ha9aa;
    defparam add_13625_25.INJECT1_0 = "NO";
    defparam add_13625_25.INJECT1_1 = "NO";
    LUT4 i4561_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[20]), .D(\result_i[16] [12]), 
         .Z(result_i_ns_0__15__N_517[252])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4561_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4553_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[21]), .D(\result_i[16] [13]), 
         .Z(result_i_ns_0__15__N_517[253])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4553_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_14 (.A0(shift_1_dout_i[11]), .B0(shift_1_dout_r[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[12]), .B1(shift_1_dout_r[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32244), .COUT(n32245), .S0(n12076), 
          .S1(n12077));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1101_add_4_12 (.A0(shift_1_dout_i[9]), .B0(shift_1_dout_r[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[10]), .B1(shift_1_dout_r[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32243), .COUT(n32244), .S0(n12074), 
          .S1(n12075));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_12.INJECT1_1 = "NO";
    CCU2C add_13625_23 (.A0(n7488), .B0(n34794), .C0(n34629), .D0(rom8_state[0]), 
          .A1(n7487), .B1(n34794), .C1(n34630), .D1(rom8_state[0]), 
          .CIN(n32431), .COUT(n32432), .S0(dout_i_23__N_4670[20]), .S1(dout_i_23__N_4670[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_23.INIT0 = 16'ha9aa;
    defparam add_13625_23.INIT1 = 16'ha9aa;
    defparam add_13625_23.INJECT1_0 = "NO";
    defparam add_13625_23.INJECT1_1 = "NO";
    LUT4 i4545_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[22]), .D(\result_i[16] [14]), 
         .Z(result_i_ns_0__15__N_517[254])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4545_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_10 (.A0(shift_1_dout_i[7]), .B0(shift_1_dout_r[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[8]), .B1(shift_1_dout_r[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32242), .COUT(n32243), .S0(n12072), 
          .S1(n12073));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_10.INJECT1_1 = "NO";
    LUT4 i4537_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_i[23]), .D(\result_i[16] [15]), 
         .Z(result_i_ns_0__15__N_517[255])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4537_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_8 (.A0(shift_1_dout_i[5]), .B0(shift_1_dout_r[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[6]), .B1(shift_1_dout_r[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32241), .COUT(n32242), .S0(n12070), 
          .S1(n12071));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_8.INJECT1_1 = "NO";
    CCU2C add_13625_21 (.A0(n7490), .B0(n34794), .C0(n34641), .D0(rom8_state[0]), 
          .A1(n7489), .B1(n34794), .C1(n34642), .D1(rom8_state[0]), 
          .CIN(n32430), .COUT(n32431), .S0(dout_i_23__N_4670[18]), .S1(dout_i_23__N_4670[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_21.INIT0 = 16'ha9aa;
    defparam add_13625_21.INIT1 = 16'ha9aa;
    defparam add_13625_21.INJECT1_0 = "NO";
    defparam add_13625_21.INJECT1_1 = "NO";
    LUT4 i8745_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[8]), .D(\result_r[16] [0]), 
         .Z(result_r_ns_0__15__N_3[240])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8745_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_6 (.A0(shift_1_dout_i[3]), .B0(shift_1_dout_r[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[4]), .B1(shift_1_dout_r[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32240), .COUT(n32241), .S0(n12068), 
          .S1(n12069));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_6.INJECT1_1 = "NO";
    LUT4 i8737_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[9]), .D(\result_r[16] [1]), 
         .Z(result_r_ns_0__15__N_3[241])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8737_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_4 (.A0(shift_1_dout_i[1]), .B0(shift_1_dout_r[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[2]), .B1(shift_1_dout_r[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32239), .COUT(n32240), .S0(n12066), 
          .S1(n12067));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1101_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_4.INJECT1_1 = "NO";
    CCU2C add_13625_19 (.A0(n7492), .B0(n34794), .C0(n34651), .D0(rom8_state[0]), 
          .A1(n7491), .B1(n34794), .C1(n34652), .D1(rom8_state[0]), 
          .CIN(n32429), .COUT(n32430), .S0(dout_i_23__N_4670[16]), .S1(dout_i_23__N_4670[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_19.INIT0 = 16'ha9aa;
    defparam add_13625_19.INIT1 = 16'ha9aa;
    defparam add_13625_19.INJECT1_0 = "NO";
    defparam add_13625_19.INJECT1_1 = "NO";
    LUT4 i8729_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[10]), .D(\result_r[16] [2]), 
         .Z(result_r_ns_0__15__N_3[242])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8729_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1101_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(shift_1_dout_i[0]), .B1(shift_1_dout_r[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32239), .S1(n12065));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1101_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1101_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1101_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1101_add_4_2.INJECT1_1 = "NO";
    LUT4 i8721_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[11]), .D(\result_r[16] [3]), 
         .Z(result_r_ns_0__15__N_3[243])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8721_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1137_add_4_18 (.A0(din_r_reg[23]), .B0(shift_16_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n32238), .S0(delay_r_23__N_1178[23]));
    defparam _add_1_1137_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_18.INIT1 = 16'h0000;
    defparam _add_1_1137_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_18.INJECT1_1 = "NO";
    CCU2C add_13625_17 (.A0(n7494), .B0(n34794), .C0(n34661), .D0(rom8_state[0]), 
          .A1(n7493), .B1(n34794), .C1(n34662), .D1(rom8_state[0]), 
          .CIN(n32428), .COUT(n32429), .S0(dout_i_23__N_4670[14]), .S1(dout_i_23__N_4670[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_17.INIT0 = 16'ha9aa;
    defparam add_13625_17.INIT1 = 16'ha9aa;
    defparam add_13625_17.INJECT1_0 = "NO";
    defparam add_13625_17.INJECT1_1 = "NO";
    LUT4 i15779_3_lut (.A(\result_r[14] [3]), .B(\result_r[15] [3]), .C(y_1_delay[0]), 
         .Z(n34163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15779_3_lut.init = 16'hcaca;
    LUT4 i8713_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[12]), .D(\result_r[16] [4]), 
         .Z(result_r_ns_0__15__N_3[244])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8713_3_lut_4_lut.init = 16'hfb40;
    PFUMX i15821 (.BLUT(n34191), .ALUT(n34192), .C0(y_1_delay[1]), .Z(n34205));
    CCU2C _add_1_1137_add_4_16 (.A0(din_r_reg[23]), .B0(shift_16_dout_r[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[23]), .B1(shift_16_dout_r[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32237), .COUT(n32238), .S0(delay_r_23__N_1178[21]), 
          .S1(delay_r_23__N_1178[22]));
    defparam _add_1_1137_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1137_add_4_14 (.A0(din_r_reg[23]), .B0(shift_16_dout_r[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[23]), .B1(shift_16_dout_r[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32236), .COUT(n32237), .S0(delay_r_23__N_1178[19]), 
          .S1(delay_r_23__N_1178[20]));
    defparam _add_1_1137_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_14.INJECT1_1 = "NO";
    CCU2C add_13625_15 (.A0(n7496), .B0(n34794), .C0(n34671), .D0(rom8_state[0]), 
          .A1(n7495), .B1(n34794), .C1(n34672), .D1(rom8_state[0]), 
          .CIN(n32427), .COUT(n32428), .S0(dout_i_23__N_4670[12]), .S1(dout_i_23__N_4670[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_15.INIT0 = 16'ha9aa;
    defparam add_13625_15.INIT1 = 16'ha9aa;
    defparam add_13625_15.INJECT1_0 = "NO";
    defparam add_13625_15.INJECT1_1 = "NO";
    CCU2C _add_1_1137_add_4_12 (.A0(din_r_reg[17]), .B0(shift_16_dout_r[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[18]), .B1(shift_16_dout_r[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32235), .COUT(n32236), .S0(delay_r_23__N_1178[17]), 
          .S1(delay_r_23__N_1178[18]));
    defparam _add_1_1137_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1137_add_4_10 (.A0(din_r_reg[15]), .B0(shift_16_dout_r[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[16]), .B1(shift_16_dout_r[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32234), .COUT(n32235), .S0(delay_r_23__N_1178[15]), 
          .S1(delay_r_23__N_1178[16]));
    defparam _add_1_1137_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_10.INJECT1_1 = "NO";
    CCU2C add_13625_13 (.A0(n7498), .B0(n34794), .C0(n34677), .D0(rom8_state[0]), 
          .A1(n7497), .B1(n34794), .C1(n34678), .D1(rom8_state[0]), 
          .CIN(n32426), .COUT(n32427), .S0(dout_i_23__N_4670[10]), .S1(dout_i_23__N_4670[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_13.INIT0 = 16'ha9aa;
    defparam add_13625_13.INIT1 = 16'ha9aa;
    defparam add_13625_13.INJECT1_0 = "NO";
    defparam add_13625_13.INJECT1_1 = "NO";
    CCU2C _add_1_1137_add_4_8 (.A0(din_r_reg[13]), .B0(shift_16_dout_r[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[14]), .B1(shift_16_dout_r[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32233), .COUT(n32234), .S0(delay_r_23__N_1178[13]), 
          .S1(delay_r_23__N_1178[14]));
    defparam _add_1_1137_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1137_add_4_6 (.A0(din_r_reg[11]), .B0(shift_16_dout_r[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[12]), .B1(shift_16_dout_r[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32232), .COUT(n32233), .S0(delay_r_23__N_1178[11]), 
          .S1(delay_r_23__N_1178[12]));
    defparam _add_1_1137_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_6.INJECT1_1 = "NO";
    CCU2C add_13625_11 (.A0(n7500), .B0(n34794), .C0(n34685), .D0(rom8_state[0]), 
          .A1(n7499), .B1(n34794), .C1(n34686), .D1(rom8_state[0]), 
          .CIN(n32425), .COUT(n32426), .S0(dout_i_23__N_4670[8]), .S1(dout_i_23__N_4670[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_11.INIT0 = 16'ha9aa;
    defparam add_13625_11.INIT1 = 16'ha9aa;
    defparam add_13625_11.INJECT1_0 = "NO";
    defparam add_13625_11.INJECT1_1 = "NO";
    LUT4 i8705_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[13]), .D(\result_r[16] [5]), 
         .Z(result_r_ns_0__15__N_3[245])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8705_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1137_add_4_4 (.A0(din_r_reg[9]), .B0(shift_16_dout_r[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(din_r_reg[10]), .B1(shift_16_dout_r[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32231), .COUT(n32232), .S0(delay_r_23__N_1178[9]), 
          .S1(delay_r_23__N_1178[10]));
    defparam _add_1_1137_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1137_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_4.INJECT1_1 = "NO";
    PFUMX i15822 (.BLUT(n34193), .ALUT(n34194), .C0(y_1_delay[1]), .Z(n34206));
    CCU2C _add_1_1137_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(din_r_reg[8]), .B1(shift_16_dout_r[8]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32231), .S1(delay_r_23__N_1178[8]));
    defparam _add_1_1137_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1137_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1137_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1137_add_4_2.INJECT1_1 = "NO";
    CCU2C add_13625_9 (.A0(n7502), .B0(n34794), .C0(radix_no1_op_i[6]), 
          .D0(rom8_state[0]), .A1(n7501), .B1(n34794), .C1(radix_no1_op_i[7]), 
          .D1(rom8_state[0]), .CIN(n32424), .COUT(n32425), .S0(dout_i_23__N_4670[6]), 
          .S1(dout_i_23__N_4670[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_9.INIT0 = 16'ha9aa;
    defparam add_13625_9.INIT1 = 16'ha9aa;
    defparam add_13625_9.INJECT1_0 = "NO";
    defparam add_13625_9.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_32 (.A0(op_r_23__N_1268_adj_7430[30]), .B0(op_i_23__N_1310_adj_7435[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[31]), 
          .B1(op_i_23__N_1310_adj_7435[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32229), .S0(op_i_23__N_1130_adj_7436[30]), .S1(op_i_23__N_1130_adj_7436[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_30 (.A0(op_r_23__N_1268_adj_7430[28]), .B0(op_i_23__N_1310_adj_7435[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[29]), 
          .B1(op_i_23__N_1310_adj_7435[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32228), .COUT(n32229), .S0(op_i_23__N_1130_adj_7436[28]), 
          .S1(op_i_23__N_1130_adj_7436[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_30.INJECT1_1 = "NO";
    CCU2C add_13625_7 (.A0(n7504), .B0(n34794), .C0(radix_no1_op_i[4]), 
          .D0(rom8_state[0]), .A1(n7503), .B1(n34794), .C1(radix_no1_op_i[5]), 
          .D1(rom8_state[0]), .CIN(n32423), .COUT(n32424), .S0(dout_i_23__N_4670[4]), 
          .S1(dout_i_23__N_4670[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_7.INIT0 = 16'ha9aa;
    defparam add_13625_7.INIT1 = 16'ha9aa;
    defparam add_13625_7.INJECT1_0 = "NO";
    defparam add_13625_7.INJECT1_1 = "NO";
    LUT4 i15778_3_lut (.A(\result_r[12] [3]), .B(\result_r[13] [3]), .C(y_1_delay[0]), 
         .Z(n34162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15778_3_lut.init = 16'hcaca;
    CCU2C _add_1_1059_add_4_28 (.A0(op_r_23__N_1268_adj_7430[26]), .B0(op_i_23__N_1310_adj_7435[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[27]), 
          .B1(op_i_23__N_1310_adj_7435[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32227), .COUT(n32228), .S0(op_i_23__N_1130_adj_7436[26]), 
          .S1(op_i_23__N_1130_adj_7436[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_26 (.A0(op_r_23__N_1268_adj_7430[24]), .B0(op_i_23__N_1310_adj_7435[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[25]), 
          .B1(op_i_23__N_1310_adj_7435[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32226), .COUT(n32227), .S0(op_i_23__N_1130_adj_7436[24]), 
          .S1(op_i_23__N_1130_adj_7436[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_26.INJECT1_1 = "NO";
    CCU2C add_13625_5 (.A0(n7506), .B0(n34794), .C0(radix_no1_op_i[2]), 
          .D0(rom8_state[0]), .A1(n7505), .B1(n34794), .C1(radix_no1_op_i[3]), 
          .D1(rom8_state[0]), .CIN(n32422), .COUT(n32423), .S0(dout_i_23__N_4670[2]), 
          .S1(dout_i_23__N_4670[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_5.INIT0 = 16'ha9aa;
    defparam add_13625_5.INIT1 = 16'ha9aa;
    defparam add_13625_5.INJECT1_0 = "NO";
    defparam add_13625_5.INJECT1_1 = "NO";
    LUT4 i15777_3_lut (.A(\result_r[10] [3]), .B(\result_r[11] [3]), .C(y_1_delay[0]), 
         .Z(n34161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15777_3_lut.init = 16'hcaca;
    CCU2C _add_1_1059_add_4_24 (.A0(op_r_23__N_1268_adj_7430[22]), .B0(op_i_23__N_1310_adj_7435[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[23]), 
          .B1(op_i_23__N_1310_adj_7435[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32225), .COUT(n32226), .S0(op_i_23__N_1130_adj_7436[22]), 
          .S1(op_i_23__N_1130_adj_7436[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_24.INJECT1_1 = "NO";
    LUT4 i15776_3_lut (.A(\result_r[8] [3]), .B(\result_r[9] [3]), .C(y_1_delay[0]), 
         .Z(n34160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15776_3_lut.init = 16'hcaca;
    LUT4 i8697_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[14]), .D(\result_r[16] [6]), 
         .Z(result_r_ns_0__15__N_3[246])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8697_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1059_add_4_22 (.A0(op_r_23__N_1268_adj_7430[20]), .B0(op_i_23__N_1310_adj_7435[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[21]), 
          .B1(op_i_23__N_1310_adj_7435[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32224), .COUT(n32225), .S0(op_i_23__N_1130_adj_7436[20]), 
          .S1(op_i_23__N_1130_adj_7436[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_22.INJECT1_1 = "NO";
    CCU2C add_13625_3 (.A0(n7508), .B0(n34794), .C0(radix_no1_op_i[0]), 
          .D0(rom8_state[0]), .A1(n7507), .B1(n34794), .C1(radix_no1_op_i[1]), 
          .D1(rom8_state[0]), .CIN(n32421), .COUT(n32422), .S0(dout_i_23__N_4670[0]), 
          .S1(dout_i_23__N_4670[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_3.INIT0 = 16'ha9aa;
    defparam add_13625_3.INIT1 = 16'ha9aa;
    defparam add_13625_3.INJECT1_0 = "NO";
    defparam add_13625_3.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_20 (.A0(op_r_23__N_1268_adj_7430[18]), .B0(op_i_23__N_1310_adj_7435[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[19]), 
          .B1(op_i_23__N_1310_adj_7435[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32223), .COUT(n32224), .S0(op_i_23__N_1130_adj_7436[18]), 
          .S1(op_i_23__N_1130_adj_7436[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_18 (.A0(op_r_23__N_1268_adj_7430[16]), .B0(op_i_23__N_1310_adj_7435[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[17]), 
          .B1(op_i_23__N_1310_adj_7435[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32222), .COUT(n32223), .S0(op_i_23__N_1130_adj_7436[16]), 
          .S1(op_i_23__N_1130_adj_7436[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_18.INJECT1_1 = "NO";
    CCU2C add_13625_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n29822), .B1(n29823), .C1(n29824), .D1(rom8_state[0]), 
          .COUT(n32421));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13625_1.INIT0 = 16'h0000;
    defparam add_13625_1.INIT1 = 16'hd8ff;
    defparam add_13625_1.INJECT1_0 = "NO";
    defparam add_13625_1.INJECT1_1 = "NO";
    LUT4 i8689_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[15]), .D(\result_r[16] [7]), 
         .Z(result_r_ns_0__15__N_3[247])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8689_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1059_add_4_16 (.A0(op_r_23__N_1268_adj_7430[14]), .B0(op_i_23__N_1310_adj_7435[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[15]), 
          .B1(op_i_23__N_1310_adj_7435[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32221), .COUT(n32222), .S0(op_i_23__N_1130_adj_7436[14]), 
          .S1(op_i_23__N_1130_adj_7436[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_14 (.A0(op_r_23__N_1268_adj_7430[12]), .B0(op_i_23__N_1310_adj_7435[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[13]), 
          .B1(op_i_23__N_1310_adj_7435[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32220), .COUT(n32221), .S0(op_i_23__N_1130_adj_7436[12]), 
          .S1(op_i_23__N_1130_adj_7436[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_14.INJECT1_1 = "NO";
    PFUMX i15823 (.BLUT(n34195), .ALUT(n34196), .C0(y_1_delay[1]), .Z(n34207));
    LUT4 i8681_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[16]), .D(\result_r[16] [8]), 
         .Z(result_r_ns_0__15__N_3[248])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8681_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1059_add_4_12 (.A0(op_r_23__N_1268_adj_7430[10]), .B0(op_i_23__N_1310_adj_7435[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[11]), 
          .B1(op_i_23__N_1310_adj_7435[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32219), .COUT(n32220), .S0(op_i_23__N_1130_adj_7436[10]), 
          .S1(op_i_23__N_1130_adj_7436[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_12.INJECT1_1 = "NO";
    LUT4 i8673_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[17]), .D(\result_r[16] [9]), 
         .Z(result_r_ns_0__15__N_3[249])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8673_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8665_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[18]), .D(\result_r[16] [10]), 
         .Z(result_r_ns_0__15__N_3[250])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8665_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1059_add_4_10 (.A0(op_r_23__N_1268_adj_7430[8]), .B0(op_i_23__N_1310_adj_7435[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[9]), 
          .B1(op_i_23__N_1310_adj_7435[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32218), .COUT(n32219), .S0(op_i_23__N_1130_adj_7436[8]), 
          .S1(op_i_23__N_1130_adj_7436[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_10.INJECT1_1 = "NO";
    LUT4 i8657_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[19]), .D(\result_r[16] [11]), 
         .Z(result_r_ns_0__15__N_3[251])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8657_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8649_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[20]), .D(\result_r[16] [12]), 
         .Z(result_r_ns_0__15__N_3[252])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8649_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1059_add_4_8 (.A0(op_r_23__N_1268_adj_7430[6]), .B0(op_i_23__N_1310_adj_7435[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[7]), 
          .B1(op_i_23__N_1310_adj_7435[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32217), .COUT(n32218));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_8.INJECT1_1 = "NO";
    LUT4 i8641_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[21]), .D(\result_r[16] [13]), 
         .Z(result_r_ns_0__15__N_3[253])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8641_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1059_add_4_6 (.A0(op_r_23__N_1268_adj_7430[4]), .B0(op_i_23__N_1310_adj_7435[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[5]), 
          .B1(op_i_23__N_1310_adj_7435[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32216), .COUT(n32217));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_6.INJECT1_1 = "NO";
    CCU2C add_13628_25 (.A0(n7539), .B0(n34794), .C0(n34615), .D0(rom8_state[0]), 
          .A1(n7538), .B1(n34794), .C1(n34616), .D1(rom8_state[0]), 
          .CIN(n32416), .S0(dout_r_23__N_4286[22]), .S1(dout_r_23__N_4286[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_25.INIT0 = 16'ha9aa;
    defparam add_13628_25.INIT1 = 16'ha9aa;
    defparam add_13628_25.INJECT1_0 = "NO";
    defparam add_13628_25.INJECT1_1 = "NO";
    CCU2C _add_1_1059_add_4_4 (.A0(op_r_23__N_1268_adj_7430[2]), .B0(op_i_23__N_1310_adj_7435[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[3]), 
          .B1(op_i_23__N_1310_adj_7435[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32215), .COUT(n32216));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1059_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_4.INJECT1_1 = "NO";
    PFUMX i15294 (.BLUT(n33664), .ALUT(n33665), .C0(y_1_delay[1]), .Z(n33678));
    CCU2C _add_1_1059_add_4_2 (.A0(op_r_23__N_1268_adj_7430[0]), .B0(op_i_23__N_1310_adj_7435[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7430[1]), 
          .B1(op_i_23__N_1310_adj_7435[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32215));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[14:35])
    defparam _add_1_1059_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1059_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1059_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1059_add_4_2.INJECT1_1 = "NO";
    CCU2C add_13628_23 (.A0(n7541), .B0(n34794), .C0(n34627), .D0(rom8_state[0]), 
          .A1(n7540), .B1(n34794), .C1(n34628), .D1(rom8_state[0]), 
          .CIN(n32415), .COUT(n32416), .S0(dout_r_23__N_4286[20]), .S1(dout_r_23__N_4286[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_23.INIT0 = 16'ha9aa;
    defparam add_13628_23.INIT1 = 16'ha9aa;
    defparam add_13628_23.INJECT1_0 = "NO";
    defparam add_13628_23.INJECT1_1 = "NO";
    LUT4 i8633_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[22]), .D(\result_r[16] [14]), 
         .Z(result_r_ns_0__15__N_3[254])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8633_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8625_3_lut_4_lut (.A(n34720), .B(n34709), .C(out_r[23]), .D(\result_r[16] [15]), 
         .Z(result_r_ns_0__15__N_3[255])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8625_3_lut_4_lut.init = 16'hfb40;
    PFUMX i15824 (.BLUT(n34197), .ALUT(n34198), .C0(y_1_delay[1]), .Z(n34208));
    CCU2C _add_1_1092_add_4_17 (.A0(n31705), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[22]), .A1(n31703), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[23]), .CIN(n32213), .S0(op_r_23__N_1106[22]), 
          .S1(op_r_23__N_1106[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_17.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_17.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_17.INJECT1_1 = "NO";
    CCU2C add_13628_21 (.A0(n7543), .B0(n34794), .C0(n34639), .D0(rom8_state[0]), 
          .A1(n7542), .B1(n34794), .C1(n34640), .D1(rom8_state[0]), 
          .CIN(n32414), .COUT(n32415), .S0(dout_r_23__N_4286[18]), .S1(dout_r_23__N_4286[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_21.INIT0 = 16'ha9aa;
    defparam add_13628_21.INIT1 = 16'ha9aa;
    defparam add_13628_21.INJECT1_0 = "NO";
    defparam add_13628_21.INJECT1_1 = "NO";
    LUT4 i4785_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[8]), .D(\result_i[17] [0]), 
         .Z(result_i_ns_0__15__N_517[224])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4785_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1092_add_4_15 (.A0(n31709), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[20]), .A1(n31707), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[21]), .CIN(n32212), .COUT(n32213), .S0(op_r_23__N_1106[20]), 
          .S1(op_r_23__N_1106[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_15.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_15.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_15.INJECT1_1 = "NO";
    LUT4 i4777_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[9]), .D(\result_i[17] [1]), 
         .Z(result_i_ns_0__15__N_517[225])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4777_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15775_3_lut (.A(\result_r[6] [3]), .B(\result_r[7] [3]), .C(y_1_delay[0]), 
         .Z(n34159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15775_3_lut.init = 16'hcaca;
    CCU2C _add_1_1092_add_4_13 (.A0(n31713), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[18]), .A1(n31711), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[19]), .CIN(n32211), .COUT(n32212), .S0(op_r_23__N_1106[18]), 
          .S1(op_r_23__N_1106[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_13.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_13.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_13.INJECT1_1 = "NO";
    CCU2C add_13628_19 (.A0(n7545), .B0(n34794), .C0(n34649), .D0(rom8_state[0]), 
          .A1(n7544), .B1(n34794), .C1(n34650), .D1(rom8_state[0]), 
          .CIN(n32413), .COUT(n32414), .S0(dout_r_23__N_4286[16]), .S1(dout_r_23__N_4286[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_19.INIT0 = 16'ha9aa;
    defparam add_13628_19.INIT1 = 16'ha9aa;
    defparam add_13628_19.INJECT1_0 = "NO";
    defparam add_13628_19.INJECT1_1 = "NO";
    LUT4 i4769_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[10]), .D(\result_i[17] [2]), 
         .Z(result_i_ns_0__15__N_517[226])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4769_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4761_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[11]), .D(\result_i[17] [3]), 
         .Z(result_i_ns_0__15__N_517[227])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4761_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4753_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[12]), .D(\result_i[17] [4]), 
         .Z(result_i_ns_0__15__N_517[228])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4753_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1092_add_4_11 (.A0(n31717), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[16]), .A1(n31715), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[17]), .CIN(n32210), .COUT(n32211), .S0(op_r_23__N_1106[16]), 
          .S1(op_r_23__N_1106[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_11.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_11.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1092_add_4_9 (.A0(n31721), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[14]), .A1(n31719), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[15]), .CIN(n32209), .COUT(n32210), .S0(op_r_23__N_1106[14]), 
          .S1(op_r_23__N_1106[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_9.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_9.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_9.INJECT1_1 = "NO";
    CCU2C add_13628_17 (.A0(n7547), .B0(n34794), .C0(n34659), .D0(rom8_state[0]), 
          .A1(n7546), .B1(n34794), .C1(n34660), .D1(rom8_state[0]), 
          .CIN(n32412), .COUT(n32413), .S0(dout_r_23__N_4286[14]), .S1(dout_r_23__N_4286[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_17.INIT0 = 16'ha9aa;
    defparam add_13628_17.INIT1 = 16'ha9aa;
    defparam add_13628_17.INJECT1_0 = "NO";
    defparam add_13628_17.INJECT1_1 = "NO";
    CCU2C _add_1_1092_add_4_7 (.A0(n31725), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[12]), .A1(n31723), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[13]), .CIN(n32208), .COUT(n32209), .S0(op_r_23__N_1106[12]), 
          .S1(op_r_23__N_1106[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_7.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_7.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_7.INJECT1_1 = "NO";
    PFUMX i15825 (.BLUT(n34199), .ALUT(n34200), .C0(y_1_delay[1]), .Z(n34209));
    CCU2C _add_1_1092_add_4_5 (.A0(n31729), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[10]), .A1(n31727), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[11]), .CIN(n32207), .COUT(n32208), .S0(op_r_23__N_1106[10]), 
          .S1(op_r_23__N_1106[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_5.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_5.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_5.INJECT1_1 = "NO";
    CCU2C add_13628_15 (.A0(n7549), .B0(n34794), .C0(n34669), .D0(rom8_state[0]), 
          .A1(n7548), .B1(n34794), .C1(n34670), .D1(rom8_state[0]), 
          .CIN(n32411), .COUT(n32412), .S0(dout_r_23__N_4286[12]), .S1(dout_r_23__N_4286[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_15.INIT0 = 16'ha9aa;
    defparam add_13628_15.INIT1 = 16'ha9aa;
    defparam add_13628_15.INJECT1_0 = "NO";
    defparam add_13628_15.INJECT1_1 = "NO";
    CCU2C _add_1_1092_add_4_3 (.A0(n31733), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_r[8]), .A1(n31731), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_r[9]), .CIN(n32206), .COUT(n32207), .S0(op_r_23__N_1106[8]), 
          .S1(op_r_23__N_1106[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_3.INIT0 = 16'h65aa;
    defparam _add_1_1092_add_4_3.INIT1 = 16'h65aa;
    defparam _add_1_1092_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1092_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[5]), .B1(count[4]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32206));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1092_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1092_add_4_1.INIT1 = 16'hfff0;
    defparam _add_1_1092_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1092_add_4_1.INJECT1_1 = "NO";
    CCU2C add_13628_13 (.A0(n7551), .B0(n34794), .C0(n34675), .D0(rom8_state[0]), 
          .A1(n7550), .B1(n34794), .C1(n34676), .D1(rom8_state[0]), 
          .CIN(n32410), .COUT(n32411), .S0(dout_r_23__N_4286[10]), .S1(dout_r_23__N_4286[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_13.INIT0 = 16'ha9aa;
    defparam add_13628_13.INIT1 = 16'ha9aa;
    defparam add_13628_13.INJECT1_0 = "NO";
    defparam add_13628_13.INJECT1_1 = "NO";
    LUT4 i4745_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[13]), .D(\result_i[17] [5]), 
         .Z(result_i_ns_0__15__N_517[229])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4745_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15774_3_lut (.A(\result_r[4] [3]), .B(\result_r[5] [3]), .C(y_1_delay[0]), 
         .Z(n34158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15774_3_lut.init = 16'hcaca;
    LUT4 i4737_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[14]), .D(\result_i[17] [6]), 
         .Z(result_i_ns_0__15__N_517[230])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4737_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_26 (.A0(op_i_23__N_1154_adj_7426[23]), .B0(n34843), 
          .C0(shift_1_dout_i[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n32202), .S0(delay_i_23__N_1202_adj_7484[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_26.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1104_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_26.INJECT1_1 = "NO";
    CCU2C add_13628_11 (.A0(n7553), .B0(n34794), .C0(n34683), .D0(rom8_state[0]), 
          .A1(n7552), .B1(n34794), .C1(n34684), .D1(rom8_state[0]), 
          .CIN(n32409), .COUT(n32410), .S0(dout_r_23__N_4286[8]), .S1(dout_r_23__N_4286[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_11.INIT0 = 16'ha9aa;
    defparam add_13628_11.INIT1 = 16'ha9aa;
    defparam add_13628_11.INJECT1_0 = "NO";
    defparam add_13628_11.INJECT1_1 = "NO";
    LUT4 i4729_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[15]), .D(\result_i[17] [7]), 
         .Z(result_i_ns_0__15__N_517[231])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4729_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4721_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[16]), .D(\result_i[17] [8]), 
         .Z(result_i_ns_0__15__N_517[232])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4721_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_24 (.A0(op_i_23__N_1154_adj_7426[21]), .B0(n34843), 
          .C0(shift_1_dout_i[21]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[22]), 
          .B1(n34843), .C1(shift_1_dout_i[22]), .D1(VCC_net), .CIN(n32201), 
          .COUT(n32202), .S0(delay_i_23__N_1202_adj_7484[21]), .S1(delay_i_23__N_1202_adj_7484[22]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_24.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_24.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_24.INJECT1_1 = "NO";
    LUT4 i15773_3_lut (.A(\result_r[2] [3]), .B(\result_r[3] [3]), .C(y_1_delay[0]), 
         .Z(n34157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15773_3_lut.init = 16'hcaca;
    CCU2C _add_1_1104_add_4_22 (.A0(op_i_23__N_1154_adj_7426[19]), .B0(n34843), 
          .C0(shift_1_dout_i[19]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[20]), 
          .B1(n34843), .C1(shift_1_dout_i[20]), .D1(VCC_net), .CIN(n32200), 
          .COUT(n32201), .S0(delay_i_23__N_1202_adj_7484[19]), .S1(delay_i_23__N_1202_adj_7484[20]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_22.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_22.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_22.INJECT1_1 = "NO";
    CCU2C add_13628_9 (.A0(n7555), .B0(n34794), .C0(radix_no1_op_r[6]), 
          .D0(rom8_state[0]), .A1(n7554), .B1(n34794), .C1(radix_no1_op_r[7]), 
          .D1(rom8_state[0]), .CIN(n32408), .COUT(n32409), .S0(dout_r_23__N_4286[6]), 
          .S1(dout_r_23__N_4286[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_9.INIT0 = 16'ha9aa;
    defparam add_13628_9.INIT1 = 16'ha9aa;
    defparam add_13628_9.INJECT1_0 = "NO";
    defparam add_13628_9.INJECT1_1 = "NO";
    LUT4 i15277_3_lut (.A(\result_i[2] [4]), .B(\result_i[3] [4]), .C(y_1_delay[0]), 
         .Z(n33661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15277_3_lut.init = 16'hcaca;
    CCU2C _add_1_1104_add_4_20 (.A0(op_i_23__N_1154_adj_7426[17]), .B0(n34843), 
          .C0(shift_1_dout_i[17]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[18]), 
          .B1(n34843), .C1(shift_1_dout_i[18]), .D1(VCC_net), .CIN(n32199), 
          .COUT(n32200), .S0(delay_i_23__N_1202_adj_7484[17]), .S1(delay_i_23__N_1202_adj_7484[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_20.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_20.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_20.INJECT1_1 = "NO";
    PFUMX i15826 (.BLUT(n34201), .ALUT(n34202), .C0(y_1_delay[1]), .Z(n34210));
    LUT4 i4713_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[17]), .D(\result_i[17] [9]), 
         .Z(result_i_ns_0__15__N_517[233])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4713_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_18 (.A0(op_i_23__N_1154_adj_7426[15]), .B0(n34843), 
          .C0(shift_1_dout_i[15]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[16]), 
          .B1(n34843), .C1(shift_1_dout_i[16]), .D1(VCC_net), .CIN(n32198), 
          .COUT(n32199), .S0(delay_i_23__N_1202_adj_7484[15]), .S1(delay_i_23__N_1202_adj_7484[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_18.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_18.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_18.INJECT1_1 = "NO";
    CCU2C add_13628_7 (.A0(n7557), .B0(n34794), .C0(radix_no1_op_r[4]), 
          .D0(rom8_state[0]), .A1(n7556), .B1(n34794), .C1(radix_no1_op_r[5]), 
          .D1(rom8_state[0]), .CIN(n32407), .COUT(n32408), .S0(dout_r_23__N_4286[4]), 
          .S1(dout_r_23__N_4286[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_7.INIT0 = 16'ha9aa;
    defparam add_13628_7.INIT1 = 16'ha9aa;
    defparam add_13628_7.INJECT1_0 = "NO";
    defparam add_13628_7.INJECT1_1 = "NO";
    LUT4 i4705_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[18]), .D(\result_i[17] [10]), 
         .Z(result_i_ns_0__15__N_517[234])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4705_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_16 (.A0(op_i_23__N_1154_adj_7426[13]), .B0(n34843), 
          .C0(shift_1_dout_i[13]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[14]), 
          .B1(n34843), .C1(shift_1_dout_i[14]), .D1(VCC_net), .CIN(n32197), 
          .COUT(n32198), .S0(delay_i_23__N_1202_adj_7484[13]), .S1(delay_i_23__N_1202_adj_7484[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_16.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_16.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1104_add_4_14 (.A0(op_i_23__N_1154_adj_7426[11]), .B0(n34843), 
          .C0(shift_1_dout_i[11]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[12]), 
          .B1(n34843), .C1(shift_1_dout_i[12]), .D1(VCC_net), .CIN(n32196), 
          .COUT(n32197), .S0(delay_i_23__N_1202_adj_7484[11]), .S1(delay_i_23__N_1202_adj_7484[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_14.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_14.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_14.INJECT1_1 = "NO";
    CCU2C add_13628_5 (.A0(n7559), .B0(n34794), .C0(radix_no1_op_r[2]), 
          .D0(rom8_state[0]), .A1(n7558), .B1(n34794), .C1(radix_no1_op_r[3]), 
          .D1(rom8_state[0]), .CIN(n32406), .COUT(n32407), .S0(dout_r_23__N_4286[2]), 
          .S1(dout_r_23__N_4286[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_5.INIT0 = 16'ha9aa;
    defparam add_13628_5.INIT1 = 16'ha9aa;
    defparam add_13628_5.INJECT1_0 = "NO";
    defparam add_13628_5.INJECT1_1 = "NO";
    CCU2C _add_1_1104_add_4_12 (.A0(op_i_23__N_1154_adj_7426[9]), .B0(n34843), 
          .C0(shift_1_dout_i[9]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[10]), 
          .B1(n34843), .C1(shift_1_dout_i[10]), .D1(VCC_net), .CIN(n32195), 
          .COUT(n32196), .S0(delay_i_23__N_1202_adj_7484[9]), .S1(delay_i_23__N_1202_adj_7484[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_12.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_12.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_12.INJECT1_1 = "NO";
    LUT4 i4697_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[19]), .D(\result_i[17] [11]), 
         .Z(result_i_ns_0__15__N_517[235])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4697_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_10 (.A0(op_i_23__N_1154_adj_7426[7]), .B0(n34843), 
          .C0(shift_1_dout_i[7]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[8]), 
          .B1(n34843), .C1(shift_1_dout_i[8]), .D1(VCC_net), .CIN(n32194), 
          .COUT(n32195), .S0(delay_i_23__N_1202_adj_7484[7]), .S1(delay_i_23__N_1202_adj_7484[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_10.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_10.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_10.INJECT1_1 = "NO";
    CCU2C add_13628_3 (.A0(n7561), .B0(n34794), .C0(radix_no1_op_r[0]), 
          .D0(rom8_state[0]), .A1(n7560), .B1(n34794), .C1(radix_no1_op_r[1]), 
          .D1(rom8_state[0]), .CIN(n32405), .COUT(n32406), .S0(dout_r_23__N_4286[0]), 
          .S1(dout_r_23__N_4286[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_3.INIT0 = 16'ha9aa;
    defparam add_13628_3.INIT1 = 16'ha9aa;
    defparam add_13628_3.INJECT1_0 = "NO";
    defparam add_13628_3.INJECT1_1 = "NO";
    LUT4 i15772_3_lut (.A(\result_r[0] [3]), .B(\result_r[1] [3]), .C(y_1_delay[0]), 
         .Z(n34156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15772_3_lut.init = 16'hcaca;
    LUT4 i4689_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[20]), .D(\result_i[17] [12]), 
         .Z(result_i_ns_0__15__N_517[236])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4689_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_8 (.A0(op_i_23__N_1154_adj_7426[5]), .B0(n34843), 
          .C0(shift_1_dout_i[5]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[6]), 
          .B1(n34843), .C1(shift_1_dout_i[6]), .D1(VCC_net), .CIN(n32193), 
          .COUT(n32194), .S0(delay_i_23__N_1202_adj_7484[5]), .S1(delay_i_23__N_1202_adj_7484[6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_8.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_8.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1104_add_4_6 (.A0(op_i_23__N_1154_adj_7426[3]), .B0(n34843), 
          .C0(shift_1_dout_i[3]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[4]), 
          .B1(n34843), .C1(shift_1_dout_i[4]), .D1(VCC_net), .CIN(n32192), 
          .COUT(n32193), .S0(delay_i_23__N_1202_adj_7484[3]), .S1(delay_i_23__N_1202_adj_7484[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_6.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_6.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_6.INJECT1_1 = "NO";
    CCU2C add_13628_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n29822), .B1(n29823), .C1(n29824), .D1(rom8_state[0]), 
          .COUT(n32405));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam add_13628_1.INIT0 = 16'h0000;
    defparam add_13628_1.INIT1 = 16'hd8ff;
    defparam add_13628_1.INJECT1_0 = "NO";
    defparam add_13628_1.INJECT1_1 = "NO";
    LUT4 i4681_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[21]), .D(\result_i[17] [13]), 
         .Z(result_i_ns_0__15__N_517[237])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4681_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_4 (.A0(op_i_23__N_1154_adj_7426[1]), .B0(n34843), 
          .C0(shift_1_dout_i[1]), .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[2]), 
          .B1(n34843), .C1(shift_1_dout_i[2]), .D1(VCC_net), .CIN(n32191), 
          .COUT(n32192), .S0(delay_i_23__N_1202_adj_7484[1]), .S1(delay_i_23__N_1202_adj_7484[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_4.INIT0 = 16'h8787;
    defparam _add_1_1104_add_4_4.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_4.INJECT1_1 = "NO";
    LUT4 i4673_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[22]), .D(\result_i[17] [14]), 
         .Z(result_i_ns_0__15__N_517[238])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4673_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1104_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(op_i_23__N_1154_adj_7426[0]), .B1(n34843), 
          .C1(shift_1_dout_i[0]), .D1(VCC_net), .COUT(n32191), .S1(delay_i_23__N_1202_adj_7484[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(37[9:28])
    defparam _add_1_1104_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1104_add_4_2.INIT1 = 16'h8787;
    defparam _add_1_1104_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1104_add_4_2.INJECT1_1 = "NO";
    PFUMX i15543 (.BLUT(n33914), .ALUT(n33915), .C0(y_1_delay[1]), .Z(n33927));
    CCU2C _add_1_985_add_4_17 (.A0(n31672), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[22]), .A1(n31670), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[23]), .CIN(n32189), .S0(op_i_23__N_1154[22]), 
          .S1(op_i_23__N_1154[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_17.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_17.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_985_add_4_15 (.A0(n31676), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[20]), .A1(n31674), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[21]), .CIN(n32188), .COUT(n32189), .S0(op_i_23__N_1154[20]), 
          .S1(op_i_23__N_1154[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_15.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_15.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_15.INJECT1_1 = "NO";
    PFUMX i15295 (.BLUT(n33666), .ALUT(n33667), .C0(y_1_delay[1]), .Z(n33679));
    CCU2C _add_1_985_add_4_13 (.A0(n31680), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[18]), .A1(n31678), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[19]), .CIN(n32187), .COUT(n32188), .S0(op_i_23__N_1154[18]), 
          .S1(op_i_23__N_1154[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_13.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_13.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_13.INJECT1_1 = "NO";
    LUT4 i4665_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_i[23]), .D(\result_i[17] [15]), 
         .Z(result_i_ns_0__15__N_517[239])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4665_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8873_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[8]), .D(\result_r[17] [0]), 
         .Z(result_r_ns_0__15__N_3[224])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8873_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_985_add_4_11 (.A0(n31684), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[16]), .A1(n31682), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[17]), .CIN(n32186), .COUT(n32187), .S0(op_i_23__N_1154[16]), 
          .S1(op_i_23__N_1154[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_11.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_11.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_11.INJECT1_1 = "NO";
    PFUMX i15199 (.BLUT(n33567), .ALUT(n33568), .C0(y_1_delay[1]), .Z(n33583));
    CCU2C _add_1_985_add_4_9 (.A0(n31688), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[14]), .A1(n31686), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[15]), .CIN(n32185), .COUT(n32186), .S0(op_i_23__N_1154[14]), 
          .S1(op_i_23__N_1154[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_9.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_9.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_9.INJECT1_1 = "NO";
    LUT4 i8865_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[9]), .D(\result_r[17] [1]), 
         .Z(result_r_ns_0__15__N_3[225])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8865_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_985_add_4_7 (.A0(n31692), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[12]), .A1(n31690), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[13]), .CIN(n32184), .COUT(n32185), .S0(op_i_23__N_1154[12]), 
          .S1(op_i_23__N_1154[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_7.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_7.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_985_add_4_5 (.A0(n31696), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[10]), .A1(n31694), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[11]), .CIN(n32183), .COUT(n32184), .S0(op_i_23__N_1154[10]), 
          .S1(op_i_23__N_1154[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_5.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_5.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_5.INJECT1_1 = "NO";
    LUT4 i8857_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[10]), .D(\result_r[17] [2]), 
         .Z(result_r_ns_0__15__N_3[226])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8857_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_985_add_4_3 (.A0(n31700), .B0(count[4]), .C0(count[5]), 
          .D0(shift_16_dout_i[8]), .A1(n31698), .B1(count[4]), .C1(count[5]), 
          .D1(shift_16_dout_i[9]), .CIN(n32182), .COUT(n32183), .S0(op_i_23__N_1154[8]), 
          .S1(op_i_23__N_1154[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_3.INIT0 = 16'h65aa;
    defparam _add_1_985_add_4_3.INIT1 = 16'h65aa;
    defparam _add_1_985_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_3.INJECT1_1 = "NO";
    LUT4 i8849_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[11]), .D(\result_r[17] [3]), 
         .Z(result_r_ns_0__15__N_3[227])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8849_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_985_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[5]), .B1(count[4]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32182));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(34[9:26])
    defparam _add_1_985_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_985_add_4_1.INIT1 = 16'hfff0;
    defparam _add_1_985_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_985_add_4_1.INJECT1_1 = "NO";
    LUT4 i8841_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[12]), .D(\result_r[17] [4]), 
         .Z(result_r_ns_0__15__N_3[228])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8841_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15508_3_lut (.A(\result_r[30] [12]), .B(\result_r[31] [12]), .C(y_1_delay[0]), 
         .Z(n33892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15508_3_lut.init = 16'hcaca;
    CCU2C _add_1_1107_add_4_26 (.A0(op_r_23__N_1106_adj_7425[23]), .B0(n34843), 
          .C0(shift_1_dout_r[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n32178), .S0(delay_r_23__N_1178_adj_7483[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_26.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1107_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_26.INJECT1_1 = "NO";
    LUT4 i8833_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[13]), .D(\result_r[17] [5]), 
         .Z(result_r_ns_0__15__N_3[229])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8833_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8825_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[14]), .D(\result_r[17] [6]), 
         .Z(result_r_ns_0__15__N_3[230])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8825_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1107_add_4_24 (.A0(op_r_23__N_1106_adj_7425[21]), .B0(n34843), 
          .C0(shift_1_dout_r[21]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[22]), 
          .B1(n34843), .C1(shift_1_dout_r[22]), .D1(VCC_net), .CIN(n32177), 
          .COUT(n32178), .S0(delay_r_23__N_1178_adj_7483[21]), .S1(delay_r_23__N_1178_adj_7483[22]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_24.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_24.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_24.INJECT1_1 = "NO";
    LUT4 i15507_3_lut (.A(\result_r[28] [12]), .B(\result_r[29] [12]), .C(y_1_delay[0]), 
         .Z(n33891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15507_3_lut.init = 16'hcaca;
    CCU2C _add_1_1107_add_4_22 (.A0(op_r_23__N_1106_adj_7425[19]), .B0(n34843), 
          .C0(shift_1_dout_r[19]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[20]), 
          .B1(n34843), .C1(shift_1_dout_r[20]), .D1(VCC_net), .CIN(n32176), 
          .COUT(n32177), .S0(delay_r_23__N_1178_adj_7483[19]), .S1(delay_r_23__N_1178_adj_7483[20]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_22.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_22.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_22.INJECT1_1 = "NO";
    LUT4 i8817_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[15]), .D(\result_r[17] [7]), 
         .Z(result_r_ns_0__15__N_3[231])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8817_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1107_add_4_20 (.A0(op_r_23__N_1106_adj_7425[17]), .B0(n34843), 
          .C0(shift_1_dout_r[17]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[18]), 
          .B1(n34843), .C1(shift_1_dout_r[18]), .D1(VCC_net), .CIN(n32175), 
          .COUT(n32176), .S0(delay_r_23__N_1178_adj_7483[17]), .S1(delay_r_23__N_1178_adj_7483[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_20.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_20.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_20.INJECT1_1 = "NO";
    PFUMX i15200 (.BLUT(n33569), .ALUT(n33570), .C0(y_1_delay[1]), .Z(n33584));
    CCU2C _add_1_1107_add_4_18 (.A0(op_r_23__N_1106_adj_7425[15]), .B0(n34843), 
          .C0(shift_1_dout_r[15]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[16]), 
          .B1(n34843), .C1(shift_1_dout_r[16]), .D1(VCC_net), .CIN(n32174), 
          .COUT(n32175), .S0(delay_r_23__N_1178_adj_7483[15]), .S1(delay_r_23__N_1178_adj_7483[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_18.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_18.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_18.INJECT1_1 = "NO";
    LUT4 i8809_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[16]), .D(\result_r[17] [8]), 
         .Z(result_r_ns_0__15__N_3[232])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8809_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1107_add_4_16 (.A0(op_r_23__N_1106_adj_7425[13]), .B0(n34843), 
          .C0(shift_1_dout_r[13]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[14]), 
          .B1(n34843), .C1(shift_1_dout_r[14]), .D1(VCC_net), .CIN(n32173), 
          .COUT(n32174), .S0(delay_r_23__N_1178_adj_7483[13]), .S1(delay_r_23__N_1178_adj_7483[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_16.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_16.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1107_add_4_14 (.A0(op_r_23__N_1106_adj_7425[11]), .B0(n34843), 
          .C0(shift_1_dout_r[11]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[12]), 
          .B1(n34843), .C1(shift_1_dout_r[12]), .D1(VCC_net), .CIN(n32172), 
          .COUT(n32173), .S0(delay_r_23__N_1178_adj_7483[11]), .S1(delay_r_23__N_1178_adj_7483[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_14.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_14.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1107_add_4_12 (.A0(op_r_23__N_1106_adj_7425[9]), .B0(n34843), 
          .C0(shift_1_dout_r[9]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[10]), 
          .B1(n34843), .C1(shift_1_dout_r[10]), .D1(VCC_net), .CIN(n32171), 
          .COUT(n32172), .S0(delay_r_23__N_1178_adj_7483[9]), .S1(delay_r_23__N_1178_adj_7483[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_12.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_12.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1107_add_4_10 (.A0(op_r_23__N_1106_adj_7425[7]), .B0(n34843), 
          .C0(shift_1_dout_r[7]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[8]), 
          .B1(n34843), .C1(shift_1_dout_r[8]), .D1(VCC_net), .CIN(n32170), 
          .COUT(n32171), .S0(delay_r_23__N_1178_adj_7483[7]), .S1(delay_r_23__N_1178_adj_7483[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_10.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_10.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_10.INJECT1_1 = "NO";
    LUT4 i8801_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[17]), .D(\result_r[17] [9]), 
         .Z(result_r_ns_0__15__N_3[233])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8801_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1107_add_4_8 (.A0(op_r_23__N_1106_adj_7425[5]), .B0(n34843), 
          .C0(shift_1_dout_r[5]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[6]), 
          .B1(n34843), .C1(shift_1_dout_r[6]), .D1(VCC_net), .CIN(n32169), 
          .COUT(n32170), .S0(delay_r_23__N_1178_adj_7483[5]), .S1(delay_r_23__N_1178_adj_7483[6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_8.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_8.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_8.INJECT1_1 = "NO";
    LUT4 i8793_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[18]), .D(\result_r[17] [10]), 
         .Z(result_r_ns_0__15__N_3[234])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8793_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1107_add_4_6 (.A0(op_r_23__N_1106_adj_7425[3]), .B0(n34843), 
          .C0(shift_1_dout_r[3]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[4]), 
          .B1(n34843), .C1(shift_1_dout_r[4]), .D1(VCC_net), .CIN(n32168), 
          .COUT(n32169), .S0(delay_r_23__N_1178_adj_7483[3]), .S1(delay_r_23__N_1178_adj_7483[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_6.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_6.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1107_add_4_4 (.A0(op_r_23__N_1106_adj_7425[1]), .B0(n34843), 
          .C0(shift_1_dout_r[1]), .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[2]), 
          .B1(n34843), .C1(shift_1_dout_r[2]), .D1(VCC_net), .CIN(n32167), 
          .COUT(n32168), .S0(delay_r_23__N_1178_adj_7483[1]), .S1(delay_r_23__N_1178_adj_7483[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_4.INIT0 = 16'h8787;
    defparam _add_1_1107_add_4_4.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_4.INJECT1_1 = "NO";
    LUT4 i8785_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[19]), .D(\result_r[17] [11]), 
         .Z(result_r_ns_0__15__N_3[235])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8785_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1107_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(op_r_23__N_1106_adj_7425[0]), .B1(n34843), 
          .C1(shift_1_dout_r[0]), .D1(VCC_net), .COUT(n32167), .S1(delay_r_23__N_1178_adj_7483[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(36[9:28])
    defparam _add_1_1107_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1107_add_4_2.INIT1 = 16'h8787;
    defparam _add_1_1107_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1107_add_4_2.INJECT1_1 = "NO";
    LUT4 i15276_3_lut (.A(\result_i[0] [4]), .B(\result_i[1] [4]), .C(y_1_delay[0]), 
         .Z(n33660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15276_3_lut.init = 16'hcaca;
    PFUMX i15544 (.BLUT(n33916), .ALUT(n33917), .C0(y_1_delay[1]), .Z(n33928));
    CCU2C _add_1_1020_add_4_32 (.A0(op_r_23__N_1268_adj_7324[30]), .B0(op_r_23__N_1226_adj_7326[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[31]), 
          .B1(op_r_23__N_1226_adj_7326[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32165), .S0(op_r_23__N_1082_adj_7327[30]), .S1(op_r_23__N_1082_adj_7327[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_32.INJECT1_1 = "NO";
    LUT4 i8777_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[20]), .D(\result_r[17] [12]), 
         .Z(result_r_ns_0__15__N_3[236])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8777_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_30 (.A0(op_r_23__N_1268_adj_7324[28]), .B0(op_r_23__N_1226_adj_7326[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[29]), 
          .B1(op_r_23__N_1226_adj_7326[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32164), .COUT(n32165), .S0(op_r_23__N_1082_adj_7327[28]), 
          .S1(op_r_23__N_1082_adj_7327[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_30.INJECT1_1 = "NO";
    CCU2C count_y_689_add_4_7 (.A0(count_y[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32392), .S0(n30));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689_add_4_7.INIT0 = 16'haaa0;
    defparam count_y_689_add_4_7.INIT1 = 16'h0000;
    defparam count_y_689_add_4_7.INJECT1_0 = "NO";
    defparam count_y_689_add_4_7.INJECT1_1 = "NO";
    LUT4 i8769_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[21]), .D(\result_r[17] [13]), 
         .Z(result_r_ns_0__15__N_3[237])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8769_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_28 (.A0(op_r_23__N_1268_adj_7324[26]), .B0(op_r_23__N_1226_adj_7326[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[27]), 
          .B1(op_r_23__N_1226_adj_7326[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32163), .COUT(n32164), .S0(op_r_23__N_1082_adj_7327[26]), 
          .S1(op_r_23__N_1082_adj_7327[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_28.INJECT1_1 = "NO";
    LUT4 i8761_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[22]), .D(\result_r[17] [14]), 
         .Z(result_r_ns_0__15__N_3[238])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8761_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_26 (.A0(op_r_23__N_1268_adj_7324[24]), .B0(op_r_23__N_1226_adj_7326[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[25]), 
          .B1(op_r_23__N_1226_adj_7326[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32162), .COUT(n32163), .S0(op_r_23__N_1082_adj_7327[24]), 
          .S1(op_r_23__N_1082_adj_7327[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_26.INJECT1_1 = "NO";
    CCU2C count_y_689_add_4_5 (.A0(count_y[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_y[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32391), .COUT(n32392), .S0(n32), .S1(n31));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689_add_4_5.INIT0 = 16'haaa0;
    defparam count_y_689_add_4_5.INIT1 = 16'haaa0;
    defparam count_y_689_add_4_5.INJECT1_0 = "NO";
    defparam count_y_689_add_4_5.INJECT1_1 = "NO";
    LUT4 i8753_3_lut_4_lut (.A(n34720), .B(n34710), .C(out_r[23]), .D(\result_r[17] [15]), 
         .Z(result_r_ns_0__15__N_3[239])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8753_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4913_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[8]), .D(\result_i[18] [0]), 
         .Z(result_i_ns_0__15__N_517[208])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4913_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_24 (.A0(op_r_23__N_1268_adj_7324[22]), .B0(op_r_23__N_1226_adj_7326[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[23]), 
          .B1(op_r_23__N_1226_adj_7326[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32161), .COUT(n32162), .S0(op_r_23__N_1082_adj_7327[22]), 
          .S1(op_r_23__N_1082_adj_7327[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_22 (.A0(op_r_23__N_1268_adj_7324[20]), .B0(op_r_23__N_1226_adj_7326[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[21]), 
          .B1(op_r_23__N_1226_adj_7326[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32160), .COUT(n32161), .S0(op_r_23__N_1082_adj_7327[20]), 
          .S1(op_r_23__N_1082_adj_7327[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_22.INJECT1_1 = "NO";
    CCU2C count_y_689_add_4_3 (.A0(count_y[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_y[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32390), .COUT(n32391), .S0(n34), .S1(n33));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689_add_4_3.INIT0 = 16'haaa0;
    defparam count_y_689_add_4_3.INIT1 = 16'haaa0;
    defparam count_y_689_add_4_3.INJECT1_0 = "NO";
    defparam count_y_689_add_4_3.INJECT1_1 = "NO";
    LUT4 i4905_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[9]), .D(\result_i[18] [1]), 
         .Z(result_i_ns_0__15__N_517[209])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4905_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_20 (.A0(op_r_23__N_1268_adj_7324[18]), .B0(op_r_23__N_1226_adj_7326[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[19]), 
          .B1(op_r_23__N_1226_adj_7326[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32159), .COUT(n32160), .S0(op_r_23__N_1082_adj_7327[18]), 
          .S1(op_r_23__N_1082_adj_7327[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_18 (.A0(op_r_23__N_1268_adj_7324[16]), .B0(op_r_23__N_1226_adj_7326[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[17]), 
          .B1(op_r_23__N_1226_adj_7326[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32158), .COUT(n32159), .S0(op_r_23__N_1082_adj_7327[16]), 
          .S1(op_r_23__N_1082_adj_7327[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_18.INJECT1_1 = "NO";
    CCU2C count_y_689_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_y[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n32390), .S1(n35));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689_add_4_1.INIT0 = 16'h0000;
    defparam count_y_689_add_4_1.INIT1 = 16'h555f;
    defparam count_y_689_add_4_1.INJECT1_0 = "NO";
    defparam count_y_689_add_4_1.INJECT1_1 = "NO";
    PFUMX i15201 (.BLUT(n33571), .ALUT(n33572), .C0(y_1_delay[1]), .Z(n33585));
    CCU2C _add_1_1020_add_4_16 (.A0(op_r_23__N_1268_adj_7324[14]), .B0(op_r_23__N_1226_adj_7326[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[15]), 
          .B1(op_r_23__N_1226_adj_7326[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32157), .COUT(n32158), .S0(op_r_23__N_1082_adj_7327[14]), 
          .S1(op_r_23__N_1082_adj_7327[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_14 (.A0(op_r_23__N_1268_adj_7324[12]), .B0(op_r_23__N_1226_adj_7326[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[13]), 
          .B1(op_r_23__N_1226_adj_7326[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32156), .COUT(n32157), .S0(op_r_23__N_1082_adj_7327[12]), 
          .S1(op_r_23__N_1082_adj_7327[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_12 (.A0(op_r_23__N_1268_adj_7324[10]), .B0(op_r_23__N_1226_adj_7326[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[11]), 
          .B1(op_r_23__N_1226_adj_7326[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32155), .COUT(n32156), .S0(op_r_23__N_1082_adj_7327[10]), 
          .S1(op_r_23__N_1082_adj_7327[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_10 (.A0(op_r_23__N_1268_adj_7324[8]), .B0(op_r_23__N_1226_adj_7326[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[9]), 
          .B1(op_r_23__N_1226_adj_7326[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32154), .COUT(n32155), .S0(op_r_23__N_1082_adj_7327[8]), 
          .S1(op_r_23__N_1082_adj_7327[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_10.INJECT1_1 = "NO";
    LUT4 i4897_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[10]), .D(\result_i[18] [2]), 
         .Z(result_i_ns_0__15__N_517[210])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4897_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_8 (.A0(op_r_23__N_1268_adj_7324[6]), .B0(op_r_23__N_1226_adj_7326[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[7]), 
          .B1(op_r_23__N_1226_adj_7326[7]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32153), .COUT(n32154));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_6 (.A0(op_r_23__N_1268_adj_7324[4]), .B0(op_r_23__N_1226_adj_7326[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[5]), 
          .B1(op_r_23__N_1226_adj_7326[5]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32152), .COUT(n32153));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_6.INJECT1_1 = "NO";
    LUT4 i4889_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[11]), .D(\result_i[18] [3]), 
         .Z(result_i_ns_0__15__N_517[211])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4889_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1020_add_4_4 (.A0(op_r_23__N_1268_adj_7324[2]), .B0(op_r_23__N_1226_adj_7326[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[3]), 
          .B1(op_r_23__N_1226_adj_7326[3]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32151), .COUT(n32152));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_2 (.A0(op_r_23__N_1268_adj_7324[0]), .B0(op_r_23__N_1226_adj_7326[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_r_23__N_1268_adj_7324[1]), 
          .B1(op_r_23__N_1226_adj_7326[1]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32151));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:35])
    defparam _add_1_1020_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1020_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1020_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_2.INJECT1_1 = "NO";
    LUT4 i4881_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[12]), .D(\result_i[18] [4]), 
         .Z(result_i_ns_0__15__N_517[212])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4881_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4873_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[13]), .D(\result_i[18] [5]), 
         .Z(result_i_ns_0__15__N_517[213])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4873_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4865_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[14]), .D(\result_i[18] [6]), 
         .Z(result_i_ns_0__15__N_517[214])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4865_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1051_add_4_25 (.A0(shift_2_dout_r[22]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[30]), .D0(n34578), .A1(shift_2_dout_r[23]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[31]), .D1(n34577), 
          .CIN(n32149), .S0(op_r_23__N_1106_adj_7425[22]), .S1(op_r_23__N_1106_adj_7425[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_25 (.A0(shift_1_dout_r[23]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[23]), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n32386), .S0(op_r_23__N_1106_adj_7481[23]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_25.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_25.INIT1 = 16'h0000;
    defparam _add_1_1073_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_25.INJECT1_1 = "NO";
    LUT4 i4857_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[15]), .D(\result_i[18] [7]), 
         .Z(result_i_ns_0__15__N_517[215])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4857_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1051_add_4_23 (.A0(shift_2_dout_r[20]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[28]), .D0(n34582), .A1(shift_2_dout_r[21]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[29]), .D1(n34581), 
          .CIN(n32148), .COUT(n32149), .S0(op_r_23__N_1106_adj_7425[20]), 
          .S1(op_r_23__N_1106_adj_7425[21]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_23.INJECT1_1 = "NO";
    LUT4 i4849_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[16]), .D(\result_i[18] [8]), 
         .Z(result_i_ns_0__15__N_517[216])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4849_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1051_add_4_21 (.A0(shift_2_dout_r[18]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[26]), .D0(n34586), .A1(shift_2_dout_r[19]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[27]), .D1(n34585), 
          .CIN(n32147), .COUT(n32148), .S0(op_r_23__N_1106_adj_7425[18]), 
          .S1(op_r_23__N_1106_adj_7425[19]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_23 (.A0(shift_1_dout_r[21]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[21]), .A1(shift_1_dout_r[22]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[22]), .CIN(n32385), 
          .COUT(n32386), .S0(op_r_23__N_1106_adj_7481[21]), .S1(op_r_23__N_1106_adj_7481[22]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_23.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_23.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_23.INJECT1_1 = "NO";
    LUT4 i4841_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[17]), .D(\result_i[18] [9]), 
         .Z(result_i_ns_0__15__N_517[217])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4841_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4833_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[18]), .D(\result_i[18] [10]), 
         .Z(result_i_ns_0__15__N_517[218])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4833_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1051_add_4_19 (.A0(shift_2_dout_r[16]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[24]), .D0(n34594), .A1(shift_2_dout_r[17]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[25]), .D1(n34593), 
          .CIN(n32146), .COUT(n32147), .S0(op_r_23__N_1106_adj_7425[16]), 
          .S1(op_r_23__N_1106_adj_7425[17]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_19.INJECT1_1 = "NO";
    LUT4 i4825_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[19]), .D(\result_i[18] [11]), 
         .Z(result_i_ns_0__15__N_517[219])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4825_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1051_add_4_17 (.A0(shift_2_dout_r[14]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[22]), .D0(n34602), .A1(shift_2_dout_r[15]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[23]), .D1(n34601), 
          .CIN(n32145), .COUT(n32146), .S0(op_r_23__N_1106_adj_7425[14]), 
          .S1(op_r_23__N_1106_adj_7425[15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_21 (.A0(shift_1_dout_r[19]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[19]), .A1(shift_1_dout_r[20]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[20]), .CIN(n32384), 
          .COUT(n32385), .S0(op_r_23__N_1106_adj_7481[19]), .S1(op_r_23__N_1106_adj_7481[20]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_21.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_21.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_21.INJECT1_1 = "NO";
    PFUMX i15202 (.BLUT(n33573), .ALUT(n33574), .C0(y_1_delay[1]), .Z(n33586));
    CCU2C _add_1_1051_add_4_15 (.A0(shift_2_dout_r[12]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[20]), .D0(n34610), .A1(shift_2_dout_r[13]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[21]), .D1(n34609), 
          .CIN(n32144), .COUT(n32145), .S0(op_r_23__N_1106_adj_7425[12]), 
          .S1(op_r_23__N_1106_adj_7425[13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1051_add_4_13 (.A0(shift_2_dout_r[10]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[18]), .D0(n34622), .A1(shift_2_dout_r[11]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[19]), .D1(n34621), 
          .CIN(n32143), .COUT(n32144), .S0(op_r_23__N_1106_adj_7425[10]), 
          .S1(op_r_23__N_1106_adj_7425[11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_19 (.A0(shift_1_dout_r[17]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[17]), .A1(shift_1_dout_r[18]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[18]), .CIN(n32383), 
          .COUT(n32384), .S0(op_r_23__N_1106_adj_7481[17]), .S1(op_r_23__N_1106_adj_7481[18]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_19.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_19.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1051_add_4_11 (.A0(shift_2_dout_r[8]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[16]), .D0(n34634), .A1(shift_2_dout_r[9]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[17]), .D1(n34633), 
          .CIN(n32142), .COUT(n32143), .S0(op_r_23__N_1106_adj_7425[8]), 
          .S1(op_r_23__N_1106_adj_7425[9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1051_add_4_9 (.A0(shift_2_dout_r[6]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[14]), .D0(n34666), .A1(shift_2_dout_r[7]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[15]), .D1(n34665), 
          .CIN(n32141), .COUT(n32142), .S0(op_r_23__N_1106_adj_7425[6]), 
          .S1(op_r_23__N_1106_adj_7425[7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_17 (.A0(shift_1_dout_r[15]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[15]), .A1(shift_1_dout_r[16]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[16]), .CIN(n32382), 
          .COUT(n32383), .S0(op_r_23__N_1106_adj_7481[15]), .S1(op_r_23__N_1106_adj_7481[16]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_17.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_17.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_17.INJECT1_1 = "NO";
    PFUMX i15296 (.BLUT(n33668), .ALUT(n33669), .C0(y_1_delay[1]), .Z(n33680));
    CCU2C _add_1_1051_add_4_7 (.A0(shift_2_dout_r[4]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[12]), .D0(n34674), .A1(shift_2_dout_r[5]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[13]), .D1(n34673), 
          .CIN(n32140), .COUT(n32141), .S0(op_r_23__N_1106_adj_7425[4]), 
          .S1(op_r_23__N_1106_adj_7425[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1051_add_4_5 (.A0(shift_2_dout_r[2]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[10]), .D0(n34680), .A1(shift_2_dout_r[3]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[11]), .D1(n34679), 
          .CIN(n32139), .COUT(n32140), .S0(op_r_23__N_1106_adj_7425[2]), 
          .S1(op_r_23__N_1106_adj_7425[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_15 (.A0(shift_1_dout_r[13]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[13]), .A1(shift_1_dout_r[14]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[14]), .CIN(n32381), 
          .COUT(n32382), .S0(op_r_23__N_1106_adj_7481[13]), .S1(op_r_23__N_1106_adj_7481[14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_15.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_15.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_15.INJECT1_1 = "NO";
    LUT4 i4817_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[20]), .D(\result_i[18] [12]), 
         .Z(result_i_ns_0__15__N_517[220])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4817_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4809_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[21]), .D(\result_i[18] [13]), 
         .Z(result_i_ns_0__15__N_517[221])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4809_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1051_add_4_3 (.A0(shift_2_dout_r[0]), .B0(state_1__N_5843[1]), 
          .C0(op_r_23__N_1082_adj_7433[8]), .D0(n34690), .A1(shift_2_dout_r[1]), 
          .B1(state_1__N_5843[1]), .C1(op_r_23__N_1082_adj_7433[9]), .D1(n34689), 
          .CIN(n32138), .COUT(n32139), .S0(op_r_23__N_1106_adj_7425[0]), 
          .S1(op_r_23__N_1106_adj_7425[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1051_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1051_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_3.INJECT1_1 = "NO";
    PFUMX i15545 (.BLUT(n33918), .ALUT(n33919), .C0(y_1_delay[1]), .Z(n33929));
    CCU2C _add_1_1051_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n34800), .B1(n34801), .C1(count_adj_7456[1]), 
          .D1(s_count_adj_7458[1]), .COUT(n32138));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1051_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1051_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1051_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1051_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_13 (.A0(shift_1_dout_r[11]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[11]), .A1(shift_1_dout_r[12]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[12]), .CIN(n32380), 
          .COUT(n32381), .S0(op_r_23__N_1106_adj_7481[11]), .S1(op_r_23__N_1106_adj_7481[12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_13.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_13.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_13.INJECT1_1 = "NO";
    LUT4 i4801_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[22]), .D(\result_i[18] [14]), 
         .Z(result_i_ns_0__15__N_517[222])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4801_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4793_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_i[23]), .D(\result_i[18] [15]), 
         .Z(result_i_ns_0__15__N_517[223])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4793_3_lut_4_lut.init = 16'hfb40;
    LUT4 i9001_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[8]), .D(\result_r[18] [0]), 
         .Z(result_r_ns_0__15__N_3[208])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9001_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_26 (.A0(shift_16_dout_i[23]), .B0(shift_16_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[23]), .B1(shift_16_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32133), .S0(n12337), .S1(n12338));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_11 (.A0(shift_1_dout_r[9]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[9]), .A1(shift_1_dout_r[10]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[10]), .CIN(n32379), 
          .COUT(n32380), .S0(op_r_23__N_1106_adj_7481[9]), .S1(op_r_23__N_1106_adj_7481[10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_11.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_11.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_11.INJECT1_1 = "NO";
    LUT4 i15506_3_lut (.A(\result_r[26] [12]), .B(\result_r[27] [12]), .C(y_1_delay[0]), 
         .Z(n33890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15506_3_lut.init = 16'hcaca;
    LUT4 i8993_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[9]), .D(\result_r[18] [1]), 
         .Z(result_r_ns_0__15__N_3[209])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8993_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_24 (.A0(shift_16_dout_i[21]), .B0(shift_16_dout_r[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[22]), .B1(shift_16_dout_r[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32132), .COUT(n32133), .S0(n12335), 
          .S1(n12336));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_24.INJECT1_1 = "NO";
    LUT4 i8985_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[10]), .D(\result_r[18] [2]), 
         .Z(result_r_ns_0__15__N_3[210])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8985_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15505_3_lut (.A(\result_r[24] [12]), .B(\result_r[25] [12]), .C(y_1_delay[0]), 
         .Z(n33889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15505_3_lut.init = 16'hcaca;
    CCU2C _add_1_1128_add_4_22 (.A0(shift_16_dout_i[19]), .B0(shift_16_dout_r[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[20]), .B1(shift_16_dout_r[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32131), .COUT(n32132), .S0(n12333), 
          .S1(n12334));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_9 (.A0(shift_1_dout_r[7]), .B0(n34769), .C0(n34839), 
          .D0(op_r_23__N_1106_adj_7425[7]), .A1(shift_1_dout_r[8]), .B1(n34769), 
          .C1(n34839), .D1(op_r_23__N_1106_adj_7425[8]), .CIN(n32378), 
          .COUT(n32379), .S1(op_r_23__N_1106_adj_7481[8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_9.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_9.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_9.INJECT1_1 = "NO";
    LUT4 i8977_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[11]), .D(\result_r[18] [3]), 
         .Z(result_r_ns_0__15__N_3[211])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8977_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8969_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[12]), .D(\result_r[18] [4]), 
         .Z(result_r_ns_0__15__N_3[212])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8969_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_20 (.A0(shift_16_dout_i[17]), .B0(shift_16_dout_r[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[18]), .B1(shift_16_dout_r[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32130), .COUT(n32131), .S0(n12331), 
          .S1(n12332));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_20.INJECT1_1 = "NO";
    LUT4 i8961_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[13]), .D(\result_r[18] [5]), 
         .Z(result_r_ns_0__15__N_3[213])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8961_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_18 (.A0(shift_16_dout_i[15]), .B0(shift_16_dout_r[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[16]), .B1(shift_16_dout_r[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32129), .COUT(n32130), .S0(n12329), 
          .S1(n12330));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_7 (.A0(shift_1_dout_r[5]), .B0(n34769), .C0(count_adj_7456[1]), 
          .D0(op_r_23__N_1106_adj_7425[5]), .A1(shift_1_dout_r[6]), .B1(n34769), 
          .C1(count_adj_7456[1]), .D1(op_r_23__N_1106_adj_7425[6]), .CIN(n32377), 
          .COUT(n32378));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_7.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_7.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_7.INJECT1_1 = "NO";
    LUT4 i8953_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[14]), .D(\result_r[18] [6]), 
         .Z(result_r_ns_0__15__N_3[214])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8953_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8945_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[15]), .D(\result_r[18] [7]), 
         .Z(result_r_ns_0__15__N_3[215])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8945_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8937_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[16]), .D(\result_r[18] [8]), 
         .Z(result_r_ns_0__15__N_3[216])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8937_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_16 (.A0(shift_16_dout_i[13]), .B0(shift_16_dout_r[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[14]), .B1(shift_16_dout_r[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32128), .COUT(n32129), .S0(n12327), 
          .S1(n12328));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_16.INJECT1_1 = "NO";
    LUT4 i8929_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[17]), .D(\result_r[18] [9]), 
         .Z(result_r_ns_0__15__N_3[217])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8929_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8921_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[18]), .D(\result_r[18] [10]), 
         .Z(result_r_ns_0__15__N_3[218])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8921_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_14 (.A0(shift_16_dout_i[11]), .B0(shift_16_dout_r[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[12]), .B1(shift_16_dout_r[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32127), .COUT(n32128), .S0(n12325), 
          .S1(n12326));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_5 (.A0(shift_1_dout_r[3]), .B0(n34769), .C0(count_adj_7456[1]), 
          .D0(op_r_23__N_1106_adj_7425[3]), .A1(shift_1_dout_r[4]), .B1(n34769), 
          .C1(count_adj_7456[1]), .D1(op_r_23__N_1106_adj_7425[4]), .CIN(n32376), 
          .COUT(n32377));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_5.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_5.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_5.INJECT1_1 = "NO";
    LUT4 i8913_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[19]), .D(\result_r[18] [11]), 
         .Z(result_r_ns_0__15__N_3[219])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8913_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8905_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[20]), .D(\result_r[18] [12]), 
         .Z(result_r_ns_0__15__N_3[220])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8905_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_12 (.A0(shift_16_dout_i[9]), .B0(shift_16_dout_r[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[10]), .B1(shift_16_dout_r[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32126), .COUT(n32127), .S0(n12323), 
          .S1(n12324));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_12.INJECT1_1 = "NO";
    LUT4 i8897_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[21]), .D(\result_r[18] [13]), 
         .Z(result_r_ns_0__15__N_3[221])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8897_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_10 (.A0(op_i_23__N_1154[7]), .B0(op_r_23__N_1106[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_16_dout_i[8]), .B1(shift_16_dout_r[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32125), .COUT(n32126), .S0(n12321), 
          .S1(n12322));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_3 (.A0(shift_1_dout_r[1]), .B0(n34769), .C0(count_adj_7456[1]), 
          .D0(op_r_23__N_1106_adj_7425[1]), .A1(shift_1_dout_r[2]), .B1(n34769), 
          .C1(count_adj_7456[1]), .D1(op_r_23__N_1106_adj_7425[2]), .CIN(n32375), 
          .COUT(n32376));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_3.INIT0 = 16'h56aa;
    defparam _add_1_1073_add_4_3.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_3.INJECT1_1 = "NO";
    LUT4 i8889_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[22]), .D(\result_r[18] [14]), 
         .Z(result_r_ns_0__15__N_3[222])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8889_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8881_3_lut_4_lut (.A(n34720), .B(n34711), .C(out_r[23]), .D(\result_r[18] [15]), 
         .Z(result_r_ns_0__15__N_3[223])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i8881_3_lut_4_lut.init = 16'hfb40;
    CCU2C _add_1_1128_add_4_8 (.A0(op_i_23__N_1154[5]), .B0(op_r_23__N_1106[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[6]), .B1(op_r_23__N_1106[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32124), .COUT(n32125), .S0(n12319), 
          .S1(n12320));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_8.INJECT1_1 = "NO";
    LUT4 i5041_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[8]), .D(\result_i[19] [0]), 
         .Z(result_i_ns_0__15__N_517[192])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5041_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_1128_add_4_6 (.A0(op_i_23__N_1154[3]), .B0(op_r_23__N_1106[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[4]), .B1(op_r_23__N_1106[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32123), .COUT(n32124), .S0(n12317), 
          .S1(n12318));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(shift_1_dout_r[0]), .B1(n34769), .C1(count_adj_7456[1]), 
          .D1(op_r_23__N_1106_adj_7425[0]), .COUT(n32375));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(33[9:26])
    defparam _add_1_1073_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1073_add_4_1.INIT1 = 16'h56aa;
    defparam _add_1_1073_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_1.INJECT1_1 = "NO";
    LUT4 i5033_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[9]), .D(\result_i[19] [1]), 
         .Z(result_i_ns_0__15__N_517[193])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5033_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_1128_add_4_4 (.A0(op_i_23__N_1154[1]), .B0(op_r_23__N_1106[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(op_i_23__N_1154[2]), .B1(op_r_23__N_1106[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32122), .COUT(n32123), .S0(n12315), 
          .S1(n12316));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1128_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_4.INJECT1_1 = "NO";
    LUT4 i5025_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[10]), .D(\result_i[19] [2]), 
         .Z(result_i_ns_0__15__N_517[194])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5025_3_lut_4_lut.init = 16'hf780;
    LUT4 i5017_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[11]), .D(\result_i[19] [3]), 
         .Z(result_i_ns_0__15__N_517[195])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5017_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_1128_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(op_i_23__N_1154[0]), .B1(op_r_23__N_1106[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n32122), .S1(n12314));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1128_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1128_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1128_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1128_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_26 (.A0(shift_1_dout_i[23]), .B0(shift_1_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n32374), .S0(n319_adj_7163));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_26.INIT1 = 16'h0000;
    defparam _add_1_1070_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_26.INJECT1_1 = "NO";
    LUT4 i5009_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[12]), .D(\result_i[19] [4]), 
         .Z(result_i_ns_0__15__N_517[196])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5009_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_1110_add_4_26 (.A0(shift_2_dout_i[23]), .B0(shift_2_dout_r[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[23]), .B1(shift_2_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32120), .S0(n12175), .S1(n12176));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1110_add_4_24 (.A0(shift_2_dout_i[21]), .B0(shift_2_dout_r[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[22]), .B1(shift_2_dout_r[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32119), .COUT(n32120), .S0(n12173), 
          .S1(n12174));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_24 (.A0(shift_1_dout_i[22]), .B0(shift_1_dout_r[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[23]), .B1(shift_1_dout_r[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32373), .COUT(n32374), .S0(n11578), 
          .S1(n11579));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_24.INJECT1_1 = "NO";
    LUT4 i5001_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[13]), .D(\result_i[19] [5]), 
         .Z(result_i_ns_0__15__N_517[197])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5001_3_lut_4_lut.init = 16'hf780;
    LUT4 i4993_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[14]), .D(\result_i[19] [6]), 
         .Z(result_i_ns_0__15__N_517[198])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4993_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_1110_add_4_22 (.A0(shift_2_dout_i[19]), .B0(shift_2_dout_r[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[20]), .B1(shift_2_dout_r[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32118), .COUT(n32119), .S0(n12171), 
          .S1(n12172));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_22.INJECT1_1 = "NO";
    PFUMX i15664 (.BLUT(n34032), .ALUT(n34033), .C0(y_1_delay[1]), .Z(n34048));
    CCU2C _add_1_1110_add_4_20 (.A0(shift_2_dout_i[17]), .B0(shift_2_dout_r[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_2_dout_i[18]), .B1(shift_2_dout_r[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32117), .COUT(n32118), .S0(n12169), 
          .S1(n12170));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[20:27])
    defparam _add_1_1110_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1110_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1110_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1110_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_22 (.A0(shift_1_dout_i[20]), .B0(shift_1_dout_r[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(shift_1_dout_i[21]), .B1(shift_1_dout_r[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n32372), .COUT(n32373), .S0(n11576), 
          .S1(n11577));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(54[20:27])
    defparam _add_1_1070_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1070_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1070_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_22.INJECT1_1 = "NO";
    LUT4 i4985_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[15]), .D(\result_i[19] [7]), 
         .Z(result_i_ns_0__15__N_517[199])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4985_3_lut_4_lut.init = 16'hf780;
    LUT4 i4977_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[16]), .D(\result_i[19] [8]), 
         .Z(result_i_ns_0__15__N_517[200])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4977_3_lut_4_lut.init = 16'hf780;
    LUT4 i4969_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[17]), .D(\result_i[19] [9]), 
         .Z(result_i_ns_0__15__N_517[201])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4969_3_lut_4_lut.init = 16'hf780;
    LUT4 i4961_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[18]), .D(\result_i[19] [10]), 
         .Z(result_i_ns_0__15__N_517[202])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4961_3_lut_4_lut.init = 16'hf780;
    LUT4 i4953_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[19]), .D(\result_i[19] [11]), 
         .Z(result_i_ns_0__15__N_517[203])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4953_3_lut_4_lut.init = 16'hf780;
    LUT4 i4945_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[20]), .D(\result_i[19] [12]), 
         .Z(result_i_ns_0__15__N_517[204])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4945_3_lut_4_lut.init = 16'hf780;
    LUT4 i4937_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[21]), .D(\result_i[19] [13]), 
         .Z(result_i_ns_0__15__N_517[205])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4937_3_lut_4_lut.init = 16'hf780;
    LUT4 i4929_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[22]), .D(\result_i[19] [14]), 
         .Z(result_i_ns_0__15__N_517[206])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4929_3_lut_4_lut.init = 16'hf780;
    LUT4 i4921_3_lut_4_lut (.A(n6), .B(n34708), .C(out_i[23]), .D(\result_i[19] [15]), 
         .Z(result_i_ns_0__15__N_517[207])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i4921_3_lut_4_lut.init = 16'hf780;
    LUT4 i9129_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[8]), .D(\result_r[19] [0]), 
         .Z(result_r_ns_0__15__N_3[192])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9129_3_lut_4_lut.init = 16'hf780;
    LUT4 i9121_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[9]), .D(\result_r[19] [1]), 
         .Z(result_r_ns_0__15__N_3[193])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9121_3_lut_4_lut.init = 16'hf780;
    LUT4 i9113_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[10]), .D(\result_r[19] [2]), 
         .Z(result_r_ns_0__15__N_3[194])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9113_3_lut_4_lut.init = 16'hf780;
    LUT4 i9105_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[11]), .D(\result_r[19] [3]), 
         .Z(result_r_ns_0__15__N_3[195])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9105_3_lut_4_lut.init = 16'hf780;
    LUT4 i9097_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[12]), .D(\result_r[19] [4]), 
         .Z(result_r_ns_0__15__N_3[196])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9097_3_lut_4_lut.init = 16'hf780;
    LUT4 i9089_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[13]), .D(\result_r[19] [5]), 
         .Z(result_r_ns_0__15__N_3[197])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9089_3_lut_4_lut.init = 16'hf780;
    LUT4 i9081_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[14]), .D(\result_r[19] [6]), 
         .Z(result_r_ns_0__15__N_3[198])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9081_3_lut_4_lut.init = 16'hf780;
    LUT4 i9073_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[15]), .D(\result_r[19] [7]), 
         .Z(result_r_ns_0__15__N_3[199])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9073_3_lut_4_lut.init = 16'hf780;
    LUT4 i9065_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[16]), .D(\result_r[19] [8]), 
         .Z(result_r_ns_0__15__N_3[200])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9065_3_lut_4_lut.init = 16'hf780;
    LUT4 i9057_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[17]), .D(\result_r[19] [9]), 
         .Z(result_r_ns_0__15__N_3[201])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9057_3_lut_4_lut.init = 16'hf780;
    LUT4 i9049_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[18]), .D(\result_r[19] [10]), 
         .Z(result_r_ns_0__15__N_3[202])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9049_3_lut_4_lut.init = 16'hf780;
    LUT4 i9041_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[19]), .D(\result_r[19] [11]), 
         .Z(result_r_ns_0__15__N_3[203])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9041_3_lut_4_lut.init = 16'hf780;
    LUT4 i9033_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[20]), .D(\result_r[19] [12]), 
         .Z(result_r_ns_0__15__N_3[204])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9033_3_lut_4_lut.init = 16'hf780;
    LUT4 i9025_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[21]), .D(\result_r[19] [13]), 
         .Z(result_r_ns_0__15__N_3[205])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9025_3_lut_4_lut.init = 16'hf780;
    LUT4 i15504_3_lut (.A(\result_r[22] [12]), .B(\result_r[23] [12]), .C(y_1_delay[0]), 
         .Z(n33888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15504_3_lut.init = 16'hcaca;
    LUT4 i9017_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[22]), .D(\result_r[19] [14]), 
         .Z(result_r_ns_0__15__N_3[206])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9017_3_lut_4_lut.init = 16'hf780;
    LUT4 i9009_3_lut_4_lut (.A(n6), .B(n34708), .C(out_r[23]), .D(\result_r[19] [15]), 
         .Z(result_r_ns_0__15__N_3[207])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9009_3_lut_4_lut.init = 16'hf780;
    LUT4 i5169_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[8]), .D(\result_i[20] [0]), 
         .Z(result_i_ns_0__15__N_517[176])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5169_3_lut_4_lut.init = 16'hf780;
    LUT4 i5161_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[9]), .D(\result_i[20] [1]), 
         .Z(result_i_ns_0__15__N_517[177])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5161_3_lut_4_lut.init = 16'hf780;
    LUT4 i15503_3_lut (.A(\result_r[20] [12]), .B(\result_r[21] [12]), .C(y_1_delay[0]), 
         .Z(n33887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15503_3_lut.init = 16'hcaca;
    LUT4 i5153_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[10]), .D(\result_i[20] [2]), 
         .Z(result_i_ns_0__15__N_517[178])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5153_3_lut_4_lut.init = 16'hf780;
    LUT4 i5145_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[11]), .D(\result_i[20] [3]), 
         .Z(result_i_ns_0__15__N_517[179])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5145_3_lut_4_lut.init = 16'hf780;
    LUT4 i5137_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[12]), .D(\result_i[20] [4]), 
         .Z(result_i_ns_0__15__N_517[180])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5137_3_lut_4_lut.init = 16'hf780;
    LUT4 i5129_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[13]), .D(\result_i[20] [5]), 
         .Z(result_i_ns_0__15__N_517[181])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5129_3_lut_4_lut.init = 16'hf780;
    LUT4 i5121_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[14]), .D(\result_i[20] [6]), 
         .Z(result_i_ns_0__15__N_517[182])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5121_3_lut_4_lut.init = 16'hf780;
    LUT4 i15659_3_lut (.A(\result_r[22] [7]), .B(\result_r[23] [7]), .C(y_1_delay[0]), 
         .Z(n34043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15659_3_lut.init = 16'hcaca;
    LUT4 i5113_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[15]), .D(\result_i[20] [7]), 
         .Z(result_i_ns_0__15__N_517[183])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5113_3_lut_4_lut.init = 16'hf780;
    LUT4 i5105_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[16]), .D(\result_i[20] [8]), 
         .Z(result_i_ns_0__15__N_517[184])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5105_3_lut_4_lut.init = 16'hf780;
    LUT4 i5097_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[17]), .D(\result_i[20] [9]), 
         .Z(result_i_ns_0__15__N_517[185])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5097_3_lut_4_lut.init = 16'hf780;
    LUT4 i5089_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[18]), .D(\result_i[20] [10]), 
         .Z(result_i_ns_0__15__N_517[186])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5089_3_lut_4_lut.init = 16'hf780;
    LUT4 i5081_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[19]), .D(\result_i[20] [11]), 
         .Z(result_i_ns_0__15__N_517[187])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5081_3_lut_4_lut.init = 16'hf780;
    LUT4 i5073_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[20]), .D(\result_i[20] [12]), 
         .Z(result_i_ns_0__15__N_517[188])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5073_3_lut_4_lut.init = 16'hf780;
    LUT4 i5065_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[21]), .D(\result_i[20] [13]), 
         .Z(result_i_ns_0__15__N_517[189])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5065_3_lut_4_lut.init = 16'hf780;
    LUT4 i5057_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[22]), .D(\result_i[20] [14]), 
         .Z(result_i_ns_0__15__N_517[190])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5057_3_lut_4_lut.init = 16'hf780;
    LUT4 i5049_3_lut_4_lut (.A(n6), .B(n34709), .C(out_i[23]), .D(\result_i[20] [15]), 
         .Z(result_i_ns_0__15__N_517[191])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5049_3_lut_4_lut.init = 16'hf780;
    LUT4 i9257_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[8]), .D(\result_r[20] [0]), 
         .Z(result_r_ns_0__15__N_3[176])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9257_3_lut_4_lut.init = 16'hf780;
    LUT4 i9249_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[9]), .D(\result_r[20] [1]), 
         .Z(result_r_ns_0__15__N_3[177])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9249_3_lut_4_lut.init = 16'hf780;
    LUT4 i9241_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[10]), .D(\result_r[20] [2]), 
         .Z(result_r_ns_0__15__N_3[178])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9241_3_lut_4_lut.init = 16'hf780;
    LUT4 i9233_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[11]), .D(\result_r[20] [3]), 
         .Z(result_r_ns_0__15__N_3[179])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9233_3_lut_4_lut.init = 16'hf780;
    LUT4 i9225_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[12]), .D(\result_r[20] [4]), 
         .Z(result_r_ns_0__15__N_3[180])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9225_3_lut_4_lut.init = 16'hf780;
    LUT4 i9217_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[13]), .D(\result_r[20] [5]), 
         .Z(result_r_ns_0__15__N_3[181])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9217_3_lut_4_lut.init = 16'hf780;
    LUT4 i9209_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[14]), .D(\result_r[20] [6]), 
         .Z(result_r_ns_0__15__N_3[182])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9209_3_lut_4_lut.init = 16'hf780;
    LUT4 i15502_3_lut (.A(\result_r[18] [12]), .B(\result_r[19] [12]), .C(y_1_delay[0]), 
         .Z(n33886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15502_3_lut.init = 16'hcaca;
    LUT4 i9201_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[15]), .D(\result_r[20] [7]), 
         .Z(result_r_ns_0__15__N_3[183])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9201_3_lut_4_lut.init = 16'hf780;
    LUT4 i9193_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[16]), .D(\result_r[20] [8]), 
         .Z(result_r_ns_0__15__N_3[184])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9193_3_lut_4_lut.init = 16'hf780;
    LUT4 i9185_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[17]), .D(\result_r[20] [9]), 
         .Z(result_r_ns_0__15__N_3[185])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9185_3_lut_4_lut.init = 16'hf780;
    LUT4 i9177_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[18]), .D(\result_r[20] [10]), 
         .Z(result_r_ns_0__15__N_3[186])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9177_3_lut_4_lut.init = 16'hf780;
    LUT4 i9169_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[19]), .D(\result_r[20] [11]), 
         .Z(result_r_ns_0__15__N_3[187])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9169_3_lut_4_lut.init = 16'hf780;
    LUT4 i9161_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[20]), .D(\result_r[20] [12]), 
         .Z(result_r_ns_0__15__N_3[188])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9161_3_lut_4_lut.init = 16'hf780;
    LUT4 i9153_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[21]), .D(\result_r[20] [13]), 
         .Z(result_r_ns_0__15__N_3[189])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9153_3_lut_4_lut.init = 16'hf780;
    LUT4 i9145_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[22]), .D(\result_r[20] [14]), 
         .Z(result_r_ns_0__15__N_3[190])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9145_3_lut_4_lut.init = 16'hf780;
    LUT4 i9137_3_lut_4_lut (.A(n6), .B(n34709), .C(out_r[23]), .D(\result_r[20] [15]), 
         .Z(result_r_ns_0__15__N_3[191])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9137_3_lut_4_lut.init = 16'hf780;
    LUT4 i5297_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[8]), .D(\result_i[21] [0]), 
         .Z(result_i_ns_0__15__N_517[160])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5297_3_lut_4_lut.init = 16'hf780;
    LUT4 i5289_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[9]), .D(\result_i[21] [1]), 
         .Z(result_i_ns_0__15__N_517[161])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5289_3_lut_4_lut.init = 16'hf780;
    LUT4 i5281_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[10]), .D(\result_i[21] [2]), 
         .Z(result_i_ns_0__15__N_517[162])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5281_3_lut_4_lut.init = 16'hf780;
    LUT4 i5273_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[11]), .D(\result_i[21] [3]), 
         .Z(result_i_ns_0__15__N_517[163])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5273_3_lut_4_lut.init = 16'hf780;
    LUT4 i5265_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[12]), .D(\result_i[21] [4]), 
         .Z(result_i_ns_0__15__N_517[164])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5265_3_lut_4_lut.init = 16'hf780;
    LUT4 i5257_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[13]), .D(\result_i[21] [5]), 
         .Z(result_i_ns_0__15__N_517[165])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5257_3_lut_4_lut.init = 16'hf780;
    LUT4 i5249_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[14]), .D(\result_i[21] [6]), 
         .Z(result_i_ns_0__15__N_517[166])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5249_3_lut_4_lut.init = 16'hf780;
    LUT4 i5241_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[15]), .D(\result_i[21] [7]), 
         .Z(result_i_ns_0__15__N_517[167])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5241_3_lut_4_lut.init = 16'hf780;
    LUT4 i5233_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[16]), .D(\result_i[21] [8]), 
         .Z(result_i_ns_0__15__N_517[168])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5233_3_lut_4_lut.init = 16'hf780;
    LUT4 i5225_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[17]), .D(\result_i[21] [9]), 
         .Z(result_i_ns_0__15__N_517[169])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5225_3_lut_4_lut.init = 16'hf780;
    LUT4 i5217_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[18]), .D(\result_i[21] [10]), 
         .Z(result_i_ns_0__15__N_517[170])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5217_3_lut_4_lut.init = 16'hf780;
    LUT4 i15501_3_lut (.A(\result_r[16] [12]), .B(\result_r[17] [12]), .C(y_1_delay[0]), 
         .Z(n33885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15501_3_lut.init = 16'hcaca;
    LUT4 i5209_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[19]), .D(\result_i[21] [11]), 
         .Z(result_i_ns_0__15__N_517[171])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5209_3_lut_4_lut.init = 16'hf780;
    LUT4 i5201_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[20]), .D(\result_i[21] [12]), 
         .Z(result_i_ns_0__15__N_517[172])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5201_3_lut_4_lut.init = 16'hf780;
    LUT4 i5193_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[21]), .D(\result_i[21] [13]), 
         .Z(result_i_ns_0__15__N_517[173])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5193_3_lut_4_lut.init = 16'hf780;
    LUT4 i5185_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[22]), .D(\result_i[21] [14]), 
         .Z(result_i_ns_0__15__N_517[174])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5185_3_lut_4_lut.init = 16'hf780;
    LUT4 i5177_3_lut_4_lut (.A(n6), .B(n34710), .C(out_i[23]), .D(\result_i[21] [15]), 
         .Z(result_i_ns_0__15__N_517[175])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5177_3_lut_4_lut.init = 16'hf780;
    LUT4 i9385_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[8]), .D(\result_r[21] [0]), 
         .Z(result_r_ns_0__15__N_3[160])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9385_3_lut_4_lut.init = 16'hf780;
    LUT4 i9377_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[9]), .D(\result_r[21] [1]), 
         .Z(result_r_ns_0__15__N_3[161])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9377_3_lut_4_lut.init = 16'hf780;
    LUT4 i9369_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[10]), .D(\result_r[21] [2]), 
         .Z(result_r_ns_0__15__N_3[162])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9369_3_lut_4_lut.init = 16'hf780;
    LUT4 i9361_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[11]), .D(\result_r[21] [3]), 
         .Z(result_r_ns_0__15__N_3[163])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9361_3_lut_4_lut.init = 16'hf780;
    LUT4 i9353_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[12]), .D(\result_r[21] [4]), 
         .Z(result_r_ns_0__15__N_3[164])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9353_3_lut_4_lut.init = 16'hf780;
    LUT4 i9345_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[13]), .D(\result_r[21] [5]), 
         .Z(result_r_ns_0__15__N_3[165])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9345_3_lut_4_lut.init = 16'hf780;
    LUT4 i9337_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[14]), .D(\result_r[21] [6]), 
         .Z(result_r_ns_0__15__N_3[166])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9337_3_lut_4_lut.init = 16'hf780;
    LUT4 i9329_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[15]), .D(\result_r[21] [7]), 
         .Z(result_r_ns_0__15__N_3[167])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9329_3_lut_4_lut.init = 16'hf780;
    LUT4 i15500_3_lut (.A(\result_r[14] [12]), .B(\result_r[15] [12]), .C(y_1_delay[0]), 
         .Z(n33884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15500_3_lut.init = 16'hcaca;
    LUT4 i9321_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[16]), .D(\result_r[21] [8]), 
         .Z(result_r_ns_0__15__N_3[168])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9321_3_lut_4_lut.init = 16'hf780;
    LUT4 i9313_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[17]), .D(\result_r[21] [9]), 
         .Z(result_r_ns_0__15__N_3[169])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9313_3_lut_4_lut.init = 16'hf780;
    LUT4 i9305_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[18]), .D(\result_r[21] [10]), 
         .Z(result_r_ns_0__15__N_3[170])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9305_3_lut_4_lut.init = 16'hf780;
    LUT4 i9297_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[19]), .D(\result_r[21] [11]), 
         .Z(result_r_ns_0__15__N_3[171])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9297_3_lut_4_lut.init = 16'hf780;
    LUT4 i9289_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[20]), .D(\result_r[21] [12]), 
         .Z(result_r_ns_0__15__N_3[172])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9289_3_lut_4_lut.init = 16'hf780;
    LUT4 i9281_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[21]), .D(\result_r[21] [13]), 
         .Z(result_r_ns_0__15__N_3[173])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9281_3_lut_4_lut.init = 16'hf780;
    LUT4 i9273_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[22]), .D(\result_r[21] [14]), 
         .Z(result_r_ns_0__15__N_3[174])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9273_3_lut_4_lut.init = 16'hf780;
    LUT4 i9265_3_lut_4_lut (.A(n6), .B(n34710), .C(out_r[23]), .D(\result_r[21] [15]), 
         .Z(result_r_ns_0__15__N_3[175])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9265_3_lut_4_lut.init = 16'hf780;
    LUT4 i5425_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[8]), .D(\result_i[22] [0]), 
         .Z(result_i_ns_0__15__N_517[144])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5425_3_lut_4_lut.init = 16'hf780;
    LUT4 i5417_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[9]), .D(\result_i[22] [1]), 
         .Z(result_i_ns_0__15__N_517[145])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5417_3_lut_4_lut.init = 16'hf780;
    LUT4 i5409_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[10]), .D(\result_i[22] [2]), 
         .Z(result_i_ns_0__15__N_517[146])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5409_3_lut_4_lut.init = 16'hf780;
    LUT4 i5401_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[11]), .D(\result_i[22] [3]), 
         .Z(result_i_ns_0__15__N_517[147])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5401_3_lut_4_lut.init = 16'hf780;
    LUT4 i5393_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[12]), .D(\result_i[22] [4]), 
         .Z(result_i_ns_0__15__N_517[148])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5393_3_lut_4_lut.init = 16'hf780;
    LUT4 i5385_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[13]), .D(\result_i[22] [5]), 
         .Z(result_i_ns_0__15__N_517[149])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5385_3_lut_4_lut.init = 16'hf780;
    LUT4 i5377_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[14]), .D(\result_i[22] [6]), 
         .Z(result_i_ns_0__15__N_517[150])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5377_3_lut_4_lut.init = 16'hf780;
    LUT4 i5369_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[15]), .D(\result_i[22] [7]), 
         .Z(result_i_ns_0__15__N_517[151])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5369_3_lut_4_lut.init = 16'hf780;
    LUT4 i5361_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[16]), .D(\result_i[22] [8]), 
         .Z(result_i_ns_0__15__N_517[152])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5361_3_lut_4_lut.init = 16'hf780;
    LUT4 i5353_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[17]), .D(\result_i[22] [9]), 
         .Z(result_i_ns_0__15__N_517[153])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5353_3_lut_4_lut.init = 16'hf780;
    LUT4 i5345_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[18]), .D(\result_i[22] [10]), 
         .Z(result_i_ns_0__15__N_517[154])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5345_3_lut_4_lut.init = 16'hf780;
    LUT4 i5337_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[19]), .D(\result_i[22] [11]), 
         .Z(result_i_ns_0__15__N_517[155])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5337_3_lut_4_lut.init = 16'hf780;
    LUT4 i5329_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[20]), .D(\result_i[22] [12]), 
         .Z(result_i_ns_0__15__N_517[156])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5329_3_lut_4_lut.init = 16'hf780;
    LUT4 i5321_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[21]), .D(\result_i[22] [13]), 
         .Z(result_i_ns_0__15__N_517[157])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5321_3_lut_4_lut.init = 16'hf780;
    LUT4 i5313_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[22]), .D(\result_i[22] [14]), 
         .Z(result_i_ns_0__15__N_517[158])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5313_3_lut_4_lut.init = 16'hf780;
    LUT4 i5305_3_lut_4_lut (.A(n6), .B(n34711), .C(out_i[23]), .D(\result_i[22] [15]), 
         .Z(result_i_ns_0__15__N_517[159])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5305_3_lut_4_lut.init = 16'hf780;
    LUT4 i9513_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[8]), .D(\result_r[22] [0]), 
         .Z(result_r_ns_0__15__N_3[144])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9513_3_lut_4_lut.init = 16'hf780;
    LUT4 i9505_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[9]), .D(\result_r[22] [1]), 
         .Z(result_r_ns_0__15__N_3[145])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9505_3_lut_4_lut.init = 16'hf780;
    LUT4 i9497_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[10]), .D(\result_r[22] [2]), 
         .Z(result_r_ns_0__15__N_3[146])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9497_3_lut_4_lut.init = 16'hf780;
    LUT4 i9489_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[11]), .D(\result_r[22] [3]), 
         .Z(result_r_ns_0__15__N_3[147])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9489_3_lut_4_lut.init = 16'hf780;
    LUT4 i15499_3_lut (.A(\result_r[12] [12]), .B(\result_r[13] [12]), .C(y_1_delay[0]), 
         .Z(n33883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15499_3_lut.init = 16'hcaca;
    LUT4 i9481_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[12]), .D(\result_r[22] [4]), 
         .Z(result_r_ns_0__15__N_3[148])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9481_3_lut_4_lut.init = 16'hf780;
    LUT4 i9473_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[13]), .D(\result_r[22] [5]), 
         .Z(result_r_ns_0__15__N_3[149])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9473_3_lut_4_lut.init = 16'hf780;
    LUT4 i9465_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[14]), .D(\result_r[22] [6]), 
         .Z(result_r_ns_0__15__N_3[150])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9465_3_lut_4_lut.init = 16'hf780;
    LUT4 i9457_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[15]), .D(\result_r[22] [7]), 
         .Z(result_r_ns_0__15__N_3[151])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9457_3_lut_4_lut.init = 16'hf780;
    LUT4 i9449_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[16]), .D(\result_r[22] [8]), 
         .Z(result_r_ns_0__15__N_3[152])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9449_3_lut_4_lut.init = 16'hf780;
    LUT4 i9441_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[17]), .D(\result_r[22] [9]), 
         .Z(result_r_ns_0__15__N_3[153])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9441_3_lut_4_lut.init = 16'hf780;
    LUT4 i9433_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[18]), .D(\result_r[22] [10]), 
         .Z(result_r_ns_0__15__N_3[154])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9433_3_lut_4_lut.init = 16'hf780;
    LUT4 i9425_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[19]), .D(\result_r[22] [11]), 
         .Z(result_r_ns_0__15__N_3[155])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9425_3_lut_4_lut.init = 16'hf780;
    LUT4 i9417_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[20]), .D(\result_r[22] [12]), 
         .Z(result_r_ns_0__15__N_3[156])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9417_3_lut_4_lut.init = 16'hf780;
    LUT4 i9409_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[21]), .D(\result_r[22] [13]), 
         .Z(result_r_ns_0__15__N_3[157])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9409_3_lut_4_lut.init = 16'hf780;
    LUT4 i9401_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[22]), .D(\result_r[22] [14]), 
         .Z(result_r_ns_0__15__N_3[158])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9401_3_lut_4_lut.init = 16'hf780;
    LUT4 i9393_3_lut_4_lut (.A(n6), .B(n34711), .C(out_r[23]), .D(\result_r[22] [15]), 
         .Z(result_r_ns_0__15__N_3[159])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9393_3_lut_4_lut.init = 16'hf780;
    LUT4 i5553_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[8]), .D(\result_i[23] [0]), 
         .Z(result_i_ns_0__15__N_517[128])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5553_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5545_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[9]), .D(\result_i[23] [1]), 
         .Z(result_i_ns_0__15__N_517[129])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5545_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5537_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[10]), .D(\result_i[23] [2]), 
         .Z(result_i_ns_0__15__N_517[130])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5537_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5529_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[11]), .D(\result_i[23] [3]), 
         .Z(result_i_ns_0__15__N_517[131])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5529_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5521_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[12]), .D(\result_i[23] [4]), 
         .Z(result_i_ns_0__15__N_517[132])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5521_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5513_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[13]), .D(\result_i[23] [5]), 
         .Z(result_i_ns_0__15__N_517[133])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5513_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5505_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[14]), .D(\result_i[23] [6]), 
         .Z(result_i_ns_0__15__N_517[134])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5505_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5497_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[15]), .D(\result_i[23] [7]), 
         .Z(result_i_ns_0__15__N_517[135])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5497_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5489_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[16]), .D(\result_i[23] [8]), 
         .Z(result_i_ns_0__15__N_517[136])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5489_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5481_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[17]), .D(\result_i[23] [9]), 
         .Z(result_i_ns_0__15__N_517[137])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5481_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5473_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[18]), .D(\result_i[23] [10]), 
         .Z(result_i_ns_0__15__N_517[138])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5473_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5465_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[19]), .D(\result_i[23] [11]), 
         .Z(result_i_ns_0__15__N_517[139])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5465_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5457_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[20]), .D(\result_i[23] [12]), 
         .Z(result_i_ns_0__15__N_517[140])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5457_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5449_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[21]), .D(\result_i[23] [13]), 
         .Z(result_i_ns_0__15__N_517[141])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5449_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5441_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[22]), .D(\result_i[23] [14]), 
         .Z(result_i_ns_0__15__N_517[142])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5441_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5433_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_i[23]), .D(\result_i[23] [15]), 
         .Z(result_i_ns_0__15__N_517[143])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5433_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9641_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[8]), .D(\result_r[23] [0]), 
         .Z(result_r_ns_0__15__N_3[128])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9641_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9633_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[9]), .D(\result_r[23] [1]), 
         .Z(result_r_ns_0__15__N_3[129])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9633_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9625_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[10]), .D(\result_r[23] [2]), 
         .Z(result_r_ns_0__15__N_3[130])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9625_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9617_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[11]), .D(\result_r[23] [3]), 
         .Z(result_r_ns_0__15__N_3[131])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9617_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9609_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[12]), .D(\result_r[23] [4]), 
         .Z(result_r_ns_0__15__N_3[132])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9609_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9601_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[13]), .D(\result_r[23] [5]), 
         .Z(result_r_ns_0__15__N_3[133])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9601_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9593_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[14]), .D(\result_r[23] [6]), 
         .Z(result_r_ns_0__15__N_3[134])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9593_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9585_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[15]), .D(\result_r[23] [7]), 
         .Z(result_r_ns_0__15__N_3[135])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9585_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9577_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[16]), .D(\result_r[23] [8]), 
         .Z(result_r_ns_0__15__N_3[136])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9577_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9569_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[17]), .D(\result_r[23] [9]), 
         .Z(result_r_ns_0__15__N_3[137])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9569_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9561_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[18]), .D(\result_r[23] [10]), 
         .Z(result_r_ns_0__15__N_3[138])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9561_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9553_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[19]), .D(\result_r[23] [11]), 
         .Z(result_r_ns_0__15__N_3[139])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9553_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9545_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[20]), .D(\result_r[23] [12]), 
         .Z(result_r_ns_0__15__N_3[140])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9545_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9537_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[21]), .D(\result_r[23] [13]), 
         .Z(result_r_ns_0__15__N_3[141])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9537_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9529_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[22]), .D(\result_r[23] [14]), 
         .Z(result_r_ns_0__15__N_3[142])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9529_3_lut_4_lut.init = 16'hfd20;
    LUT4 i9521_3_lut_4_lut (.A(n34714), .B(n34725), .C(out_r[23]), .D(\result_r[23] [15]), 
         .Z(result_r_ns_0__15__N_3[143])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9521_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5681_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[8]), .D(\result_i[24] [0]), 
         .Z(result_i_ns_0__15__N_517[112])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5681_3_lut_4_lut.init = 16'hf780;
    LUT4 i5673_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[9]), .D(\result_i[24] [1]), 
         .Z(result_i_ns_0__15__N_517[113])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5673_3_lut_4_lut.init = 16'hf780;
    LUT4 i5665_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[10]), .D(\result_i[24] [2]), 
         .Z(result_i_ns_0__15__N_517[114])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5665_3_lut_4_lut.init = 16'hf780;
    LUT4 i5657_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[11]), .D(\result_i[24] [3]), 
         .Z(result_i_ns_0__15__N_517[115])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5657_3_lut_4_lut.init = 16'hf780;
    LUT4 i5649_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[12]), .D(\result_i[24] [4]), 
         .Z(result_i_ns_0__15__N_517[116])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5649_3_lut_4_lut.init = 16'hf780;
    LUT4 i5641_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[13]), .D(\result_i[24] [5]), 
         .Z(result_i_ns_0__15__N_517[117])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5641_3_lut_4_lut.init = 16'hf780;
    LUT4 i5633_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[14]), .D(\result_i[24] [6]), 
         .Z(result_i_ns_0__15__N_517[118])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5633_3_lut_4_lut.init = 16'hf780;
    LUT4 i5625_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[15]), .D(\result_i[24] [7]), 
         .Z(result_i_ns_0__15__N_517[119])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5625_3_lut_4_lut.init = 16'hf780;
    LUT4 i5617_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[16]), .D(\result_i[24] [8]), 
         .Z(result_i_ns_0__15__N_517[120])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5617_3_lut_4_lut.init = 16'hf780;
    LUT4 i5609_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[17]), .D(\result_i[24] [9]), 
         .Z(result_i_ns_0__15__N_517[121])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5609_3_lut_4_lut.init = 16'hf780;
    LUT4 i5601_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[18]), .D(\result_i[24] [10]), 
         .Z(result_i_ns_0__15__N_517[122])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5601_3_lut_4_lut.init = 16'hf780;
    LUT4 i5593_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[19]), .D(\result_i[24] [11]), 
         .Z(result_i_ns_0__15__N_517[123])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5593_3_lut_4_lut.init = 16'hf780;
    LUT4 i5585_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[20]), .D(\result_i[24] [12]), 
         .Z(result_i_ns_0__15__N_517[124])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5585_3_lut_4_lut.init = 16'hf780;
    LUT4 i5577_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[21]), .D(\result_i[24] [13]), 
         .Z(result_i_ns_0__15__N_517[125])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5577_3_lut_4_lut.init = 16'hf780;
    LUT4 i5569_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[22]), .D(\result_i[24] [14]), 
         .Z(result_i_ns_0__15__N_517[126])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5569_3_lut_4_lut.init = 16'hf780;
    LUT4 i5561_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_i[23]), .D(\result_i[24] [15]), 
         .Z(result_i_ns_0__15__N_517[127])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5561_3_lut_4_lut.init = 16'hf780;
    LUT4 i9769_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[8]), .D(\result_r[24] [0]), 
         .Z(result_r_ns_0__15__N_3[112])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9769_3_lut_4_lut.init = 16'hf780;
    LUT4 i9761_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[9]), .D(\result_r[24] [1]), 
         .Z(result_r_ns_0__15__N_3[113])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9761_3_lut_4_lut.init = 16'hf780;
    LUT4 i9753_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[10]), .D(\result_r[24] [2]), 
         .Z(result_r_ns_0__15__N_3[114])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9753_3_lut_4_lut.init = 16'hf780;
    LUT4 i9745_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[11]), .D(\result_r[24] [3]), 
         .Z(result_r_ns_0__15__N_3[115])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9745_3_lut_4_lut.init = 16'hf780;
    LUT4 i9737_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[12]), .D(\result_r[24] [4]), 
         .Z(result_r_ns_0__15__N_3[116])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9737_3_lut_4_lut.init = 16'hf780;
    LUT4 i9729_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[13]), .D(\result_r[24] [5]), 
         .Z(result_r_ns_0__15__N_3[117])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9729_3_lut_4_lut.init = 16'hf780;
    LUT4 i9721_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[14]), .D(\result_r[24] [6]), 
         .Z(result_r_ns_0__15__N_3[118])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9721_3_lut_4_lut.init = 16'hf780;
    LUT4 i9713_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[15]), .D(\result_r[24] [7]), 
         .Z(result_r_ns_0__15__N_3[119])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9713_3_lut_4_lut.init = 16'hf780;
    LUT4 i9705_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[16]), .D(\result_r[24] [8]), 
         .Z(result_r_ns_0__15__N_3[120])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9705_3_lut_4_lut.init = 16'hf780;
    LUT4 i9697_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[17]), .D(\result_r[24] [9]), 
         .Z(result_r_ns_0__15__N_3[121])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9697_3_lut_4_lut.init = 16'hf780;
    LUT4 i9689_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[18]), .D(\result_r[24] [10]), 
         .Z(result_r_ns_0__15__N_3[122])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9689_3_lut_4_lut.init = 16'hf780;
    LUT4 i9681_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[19]), .D(\result_r[24] [11]), 
         .Z(result_r_ns_0__15__N_3[123])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9681_3_lut_4_lut.init = 16'hf780;
    LUT4 i9673_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[20]), .D(\result_r[24] [12]), 
         .Z(result_r_ns_0__15__N_3[124])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9673_3_lut_4_lut.init = 16'hf780;
    LUT4 i9665_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[21]), .D(\result_r[24] [13]), 
         .Z(result_r_ns_0__15__N_3[125])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9665_3_lut_4_lut.init = 16'hf780;
    LUT4 i9657_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[22]), .D(\result_r[24] [14]), 
         .Z(result_r_ns_0__15__N_3[126])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9657_3_lut_4_lut.init = 16'hf780;
    LUT4 i9649_3_lut_4_lut (.A(n34714), .B(n34724), .C(out_r[23]), .D(\result_r[24] [15]), 
         .Z(result_r_ns_0__15__N_3[127])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9649_3_lut_4_lut.init = 16'hf780;
    LUT4 i5809_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[8]), .D(\result_i[25] [0]), 
         .Z(result_i_ns_0__15__N_517[96])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5809_3_lut_4_lut.init = 16'hf780;
    LUT4 i5801_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[9]), .D(\result_i[25] [1]), 
         .Z(result_i_ns_0__15__N_517[97])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5801_3_lut_4_lut.init = 16'hf780;
    LUT4 i5793_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[10]), .D(\result_i[25] [2]), 
         .Z(result_i_ns_0__15__N_517[98])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5793_3_lut_4_lut.init = 16'hf780;
    LUT4 i5785_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[11]), .D(\result_i[25] [3]), 
         .Z(result_i_ns_0__15__N_517[99])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5785_3_lut_4_lut.init = 16'hf780;
    LUT4 i5777_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[12]), .D(\result_i[25] [4]), 
         .Z(result_i_ns_0__15__N_517[100])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5777_3_lut_4_lut.init = 16'hf780;
    LUT4 i5769_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[13]), .D(\result_i[25] [5]), 
         .Z(result_i_ns_0__15__N_517[101])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5769_3_lut_4_lut.init = 16'hf780;
    LUT4 i5761_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[14]), .D(\result_i[25] [6]), 
         .Z(result_i_ns_0__15__N_517[102])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5761_3_lut_4_lut.init = 16'hf780;
    LUT4 i5753_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[15]), .D(\result_i[25] [7]), 
         .Z(result_i_ns_0__15__N_517[103])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5753_3_lut_4_lut.init = 16'hf780;
    LUT4 i5745_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[16]), .D(\result_i[25] [8]), 
         .Z(result_i_ns_0__15__N_517[104])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5745_3_lut_4_lut.init = 16'hf780;
    LUT4 i5737_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[17]), .D(\result_i[25] [9]), 
         .Z(result_i_ns_0__15__N_517[105])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5737_3_lut_4_lut.init = 16'hf780;
    LUT4 i5729_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[18]), .D(\result_i[25] [10]), 
         .Z(result_i_ns_0__15__N_517[106])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5729_3_lut_4_lut.init = 16'hf780;
    LUT4 i5721_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[19]), .D(\result_i[25] [11]), 
         .Z(result_i_ns_0__15__N_517[107])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5721_3_lut_4_lut.init = 16'hf780;
    LUT4 i5713_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[20]), .D(\result_i[25] [12]), 
         .Z(result_i_ns_0__15__N_517[108])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5713_3_lut_4_lut.init = 16'hf780;
    LUT4 i5705_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[21]), .D(\result_i[25] [13]), 
         .Z(result_i_ns_0__15__N_517[109])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5705_3_lut_4_lut.init = 16'hf780;
    LUT4 i5697_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[22]), .D(\result_i[25] [14]), 
         .Z(result_i_ns_0__15__N_517[110])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5697_3_lut_4_lut.init = 16'hf780;
    LUT4 i5689_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_i[23]), .D(\result_i[25] [15]), 
         .Z(result_i_ns_0__15__N_517[111])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5689_3_lut_4_lut.init = 16'hf780;
    LUT4 i9897_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[8]), .D(\result_r[25] [0]), 
         .Z(result_r_ns_0__15__N_3[96])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9897_3_lut_4_lut.init = 16'hf780;
    LUT4 i9889_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[9]), .D(\result_r[25] [1]), 
         .Z(result_r_ns_0__15__N_3[97])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9889_3_lut_4_lut.init = 16'hf780;
    LUT4 i9881_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[10]), .D(\result_r[25] [2]), 
         .Z(result_r_ns_0__15__N_3[98])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9881_3_lut_4_lut.init = 16'hf780;
    LUT4 i9873_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[11]), .D(\result_r[25] [3]), 
         .Z(result_r_ns_0__15__N_3[99])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9873_3_lut_4_lut.init = 16'hf780;
    LUT4 i9865_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[12]), .D(\result_r[25] [4]), 
         .Z(result_r_ns_0__15__N_3[100])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9865_3_lut_4_lut.init = 16'hf780;
    LUT4 i9857_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[13]), .D(\result_r[25] [5]), 
         .Z(result_r_ns_0__15__N_3[101])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9857_3_lut_4_lut.init = 16'hf780;
    LUT4 i9849_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[14]), .D(\result_r[25] [6]), 
         .Z(result_r_ns_0__15__N_3[102])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9849_3_lut_4_lut.init = 16'hf780;
    LUT4 i9841_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[15]), .D(\result_r[25] [7]), 
         .Z(result_r_ns_0__15__N_3[103])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9841_3_lut_4_lut.init = 16'hf780;
    LUT4 i9833_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[16]), .D(\result_r[25] [8]), 
         .Z(result_r_ns_0__15__N_3[104])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9833_3_lut_4_lut.init = 16'hf780;
    LUT4 i9825_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[17]), .D(\result_r[25] [9]), 
         .Z(result_r_ns_0__15__N_3[105])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9825_3_lut_4_lut.init = 16'hf780;
    LUT4 i9817_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[18]), .D(\result_r[25] [10]), 
         .Z(result_r_ns_0__15__N_3[106])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9817_3_lut_4_lut.init = 16'hf780;
    LUT4 i9809_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[19]), .D(\result_r[25] [11]), 
         .Z(result_r_ns_0__15__N_3[107])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9809_3_lut_4_lut.init = 16'hf780;
    LUT4 i9801_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[20]), .D(\result_r[25] [12]), 
         .Z(result_r_ns_0__15__N_3[108])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9801_3_lut_4_lut.init = 16'hf780;
    LUT4 i9793_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[21]), .D(\result_r[25] [13]), 
         .Z(result_r_ns_0__15__N_3[109])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9793_3_lut_4_lut.init = 16'hf780;
    LUT4 i9785_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[22]), .D(\result_r[25] [14]), 
         .Z(result_r_ns_0__15__N_3[110])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9785_3_lut_4_lut.init = 16'hf780;
    LUT4 i9777_3_lut_4_lut (.A(n34714), .B(n34723), .C(out_r[23]), .D(\result_r[25] [15]), 
         .Z(result_r_ns_0__15__N_3[111])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9777_3_lut_4_lut.init = 16'hf780;
    LUT4 i6201_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[23]), .D(\result_i[29] [15]), 
         .Z(result_i_ns_0__15__N_517[47])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6201_3_lut_4_lut.init = 16'hf780;
    LUT4 i6209_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[22]), .D(\result_i[29] [14]), 
         .Z(result_i_ns_0__15__N_517[46])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6209_3_lut_4_lut.init = 16'hf780;
    LUT4 i6217_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[21]), .D(\result_i[29] [13]), 
         .Z(result_i_ns_0__15__N_517[45])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6217_3_lut_4_lut.init = 16'hf780;
    LUT4 i6225_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[20]), .D(\result_i[29] [12]), 
         .Z(result_i_ns_0__15__N_517[44])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6225_3_lut_4_lut.init = 16'hf780;
    LUT4 i6233_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[19]), .D(\result_i[29] [11]), 
         .Z(result_i_ns_0__15__N_517[43])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6233_3_lut_4_lut.init = 16'hf780;
    LUT4 i6241_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[18]), .D(\result_i[29] [10]), 
         .Z(result_i_ns_0__15__N_517[42])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6241_3_lut_4_lut.init = 16'hf780;
    LUT4 i6249_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[17]), .D(\result_i[29] [9]), 
         .Z(result_i_ns_0__15__N_517[41])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6249_3_lut_4_lut.init = 16'hf780;
    LUT4 i6257_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[16]), .D(\result_i[29] [8]), 
         .Z(result_i_ns_0__15__N_517[40])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6257_3_lut_4_lut.init = 16'hf780;
    LUT4 i6265_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[15]), .D(\result_i[29] [7]), 
         .Z(result_i_ns_0__15__N_517[39])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6265_3_lut_4_lut.init = 16'hf780;
    LUT4 i6273_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[14]), .D(\result_i[29] [6]), 
         .Z(result_i_ns_0__15__N_517[38])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6273_3_lut_4_lut.init = 16'hf780;
    LUT4 i6281_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[13]), .D(\result_i[29] [5]), 
         .Z(result_i_ns_0__15__N_517[37])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6281_3_lut_4_lut.init = 16'hf780;
    LUT4 i6289_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[12]), .D(\result_i[29] [4]), 
         .Z(result_i_ns_0__15__N_517[36])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6289_3_lut_4_lut.init = 16'hf780;
    LUT4 i6297_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[11]), .D(\result_i[29] [3]), 
         .Z(result_i_ns_0__15__N_517[35])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6297_3_lut_4_lut.init = 16'hf780;
    LUT4 i6305_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[10]), .D(\result_i[29] [2]), 
         .Z(result_i_ns_0__15__N_517[34])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6305_3_lut_4_lut.init = 16'hf780;
    LUT4 i6313_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[9]), .D(\result_i[29] [1]), 
         .Z(result_i_ns_0__15__N_517[33])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6313_3_lut_4_lut.init = 16'hf780;
    LUT4 i6321_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_i[8]), .D(\result_i[29] [0]), 
         .Z(result_i_ns_0__15__N_517[32])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6321_3_lut_4_lut.init = 16'hf780;
    LUT4 i10409_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[8]), .D(\result_r[29] [0]), 
         .Z(result_r_ns_0__15__N_3[32])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10409_3_lut_4_lut.init = 16'hf780;
    LUT4 i10401_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[9]), .D(\result_r[29] [1]), 
         .Z(result_r_ns_0__15__N_3[33])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10401_3_lut_4_lut.init = 16'hf780;
    LUT4 i10393_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[10]), .D(\result_r[29] [2]), 
         .Z(result_r_ns_0__15__N_3[34])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10393_3_lut_4_lut.init = 16'hf780;
    LUT4 i10385_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[11]), .D(\result_r[29] [3]), 
         .Z(result_r_ns_0__15__N_3[35])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10385_3_lut_4_lut.init = 16'hf780;
    LUT4 i10377_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[12]), .D(\result_r[29] [4]), 
         .Z(result_r_ns_0__15__N_3[36])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10377_3_lut_4_lut.init = 16'hf780;
    LUT4 i10369_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[13]), .D(\result_r[29] [5]), 
         .Z(result_r_ns_0__15__N_3[37])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10369_3_lut_4_lut.init = 16'hf780;
    LUT4 i10361_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[14]), .D(\result_r[29] [6]), 
         .Z(result_r_ns_0__15__N_3[38])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10361_3_lut_4_lut.init = 16'hf780;
    LUT4 i10353_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[15]), .D(\result_r[29] [7]), 
         .Z(result_r_ns_0__15__N_3[39])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10353_3_lut_4_lut.init = 16'hf780;
    LUT4 i10345_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[16]), .D(\result_r[29] [8]), 
         .Z(result_r_ns_0__15__N_3[40])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10345_3_lut_4_lut.init = 16'hf780;
    LUT4 i10337_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[17]), .D(\result_r[29] [9]), 
         .Z(result_r_ns_0__15__N_3[41])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10337_3_lut_4_lut.init = 16'hf780;
    LUT4 i10329_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[18]), .D(\result_r[29] [10]), 
         .Z(result_r_ns_0__15__N_3[42])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10329_3_lut_4_lut.init = 16'hf780;
    LUT4 i10321_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[19]), .D(\result_r[29] [11]), 
         .Z(result_r_ns_0__15__N_3[43])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10321_3_lut_4_lut.init = 16'hf780;
    LUT4 i10313_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[20]), .D(\result_r[29] [12]), 
         .Z(result_r_ns_0__15__N_3[44])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10313_3_lut_4_lut.init = 16'hf780;
    LUT4 i10305_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[21]), .D(\result_r[29] [13]), 
         .Z(result_r_ns_0__15__N_3[45])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10305_3_lut_4_lut.init = 16'hf780;
    LUT4 i10297_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[22]), .D(\result_r[29] [14]), 
         .Z(result_r_ns_0__15__N_3[46])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10297_3_lut_4_lut.init = 16'hf780;
    LUT4 i10289_3_lut_4_lut (.A(n34712), .B(n34723), .C(out_r[23]), .D(\result_r[29] [15]), 
         .Z(result_r_ns_0__15__N_3[47])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10289_3_lut_4_lut.init = 16'hf780;
    LUT4 i6073_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[23]), .D(\result_i[28] [15]), 
         .Z(result_i_ns_0__15__N_517[63])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6073_3_lut_4_lut.init = 16'hf780;
    LUT4 i6081_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[22]), .D(\result_i[28] [14]), 
         .Z(result_i_ns_0__15__N_517[62])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6081_3_lut_4_lut.init = 16'hf780;
    LUT4 i6089_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[21]), .D(\result_i[28] [13]), 
         .Z(result_i_ns_0__15__N_517[61])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6089_3_lut_4_lut.init = 16'hf780;
    LUT4 i6097_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[20]), .D(\result_i[28] [12]), 
         .Z(result_i_ns_0__15__N_517[60])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6097_3_lut_4_lut.init = 16'hf780;
    LUT4 i6105_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[19]), .D(\result_i[28] [11]), 
         .Z(result_i_ns_0__15__N_517[59])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6105_3_lut_4_lut.init = 16'hf780;
    LUT4 i6113_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[18]), .D(\result_i[28] [10]), 
         .Z(result_i_ns_0__15__N_517[58])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6113_3_lut_4_lut.init = 16'hf780;
    LUT4 i6121_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[17]), .D(\result_i[28] [9]), 
         .Z(result_i_ns_0__15__N_517[57])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6121_3_lut_4_lut.init = 16'hf780;
    LUT4 i6129_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[16]), .D(\result_i[28] [8]), 
         .Z(result_i_ns_0__15__N_517[56])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6129_3_lut_4_lut.init = 16'hf780;
    LUT4 i6137_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[15]), .D(\result_i[28] [7]), 
         .Z(result_i_ns_0__15__N_517[55])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6137_3_lut_4_lut.init = 16'hf780;
    LUT4 i6145_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[14]), .D(\result_i[28] [6]), 
         .Z(result_i_ns_0__15__N_517[54])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6145_3_lut_4_lut.init = 16'hf780;
    LUT4 i6153_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[13]), .D(\result_i[28] [5]), 
         .Z(result_i_ns_0__15__N_517[53])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6153_3_lut_4_lut.init = 16'hf780;
    LUT4 i6161_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[12]), .D(\result_i[28] [4]), 
         .Z(result_i_ns_0__15__N_517[52])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6161_3_lut_4_lut.init = 16'hf780;
    LUT4 i6169_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[11]), .D(\result_i[28] [3]), 
         .Z(result_i_ns_0__15__N_517[51])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6169_3_lut_4_lut.init = 16'hf780;
    LUT4 i6177_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[10]), .D(\result_i[28] [2]), 
         .Z(result_i_ns_0__15__N_517[50])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6177_3_lut_4_lut.init = 16'hf780;
    LUT4 i6185_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[9]), .D(\result_i[28] [1]), 
         .Z(result_i_ns_0__15__N_517[49])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6185_3_lut_4_lut.init = 16'hf780;
    LUT4 i6193_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_i[8]), .D(\result_i[28] [0]), 
         .Z(result_i_ns_0__15__N_517[48])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6193_3_lut_4_lut.init = 16'hf780;
    LUT4 i10281_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[8]), .D(\result_r[28] [0]), 
         .Z(result_r_ns_0__15__N_3[48])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10281_3_lut_4_lut.init = 16'hf780;
    LUT4 i10273_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[9]), .D(\result_r[28] [1]), 
         .Z(result_r_ns_0__15__N_3[49])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10273_3_lut_4_lut.init = 16'hf780;
    LUT4 i10265_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[10]), .D(\result_r[28] [2]), 
         .Z(result_r_ns_0__15__N_3[50])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10265_3_lut_4_lut.init = 16'hf780;
    LUT4 i10257_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[11]), .D(\result_r[28] [3]), 
         .Z(result_r_ns_0__15__N_3[51])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10257_3_lut_4_lut.init = 16'hf780;
    LUT4 i10249_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[12]), .D(\result_r[28] [4]), 
         .Z(result_r_ns_0__15__N_3[52])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10249_3_lut_4_lut.init = 16'hf780;
    LUT4 i10241_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[13]), .D(\result_r[28] [5]), 
         .Z(result_r_ns_0__15__N_3[53])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10241_3_lut_4_lut.init = 16'hf780;
    LUT4 i10233_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[14]), .D(\result_r[28] [6]), 
         .Z(result_r_ns_0__15__N_3[54])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10233_3_lut_4_lut.init = 16'hf780;
    LUT4 i10225_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[15]), .D(\result_r[28] [7]), 
         .Z(result_r_ns_0__15__N_3[55])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10225_3_lut_4_lut.init = 16'hf780;
    LUT4 i10217_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[16]), .D(\result_r[28] [8]), 
         .Z(result_r_ns_0__15__N_3[56])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10217_3_lut_4_lut.init = 16'hf780;
    LUT4 i10209_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[17]), .D(\result_r[28] [9]), 
         .Z(result_r_ns_0__15__N_3[57])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10209_3_lut_4_lut.init = 16'hf780;
    LUT4 i10201_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[18]), .D(\result_r[28] [10]), 
         .Z(result_r_ns_0__15__N_3[58])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10201_3_lut_4_lut.init = 16'hf780;
    LUT4 i10193_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[19]), .D(\result_r[28] [11]), 
         .Z(result_r_ns_0__15__N_3[59])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10193_3_lut_4_lut.init = 16'hf780;
    LUT4 i10185_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[20]), .D(\result_r[28] [12]), 
         .Z(result_r_ns_0__15__N_3[60])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10185_3_lut_4_lut.init = 16'hf780;
    LUT4 i10177_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[21]), .D(\result_r[28] [13]), 
         .Z(result_r_ns_0__15__N_3[61])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10177_3_lut_4_lut.init = 16'hf780;
    LUT4 i10169_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[22]), .D(\result_r[28] [14]), 
         .Z(result_r_ns_0__15__N_3[62])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10169_3_lut_4_lut.init = 16'hf780;
    LUT4 i10161_3_lut_4_lut (.A(n34712), .B(n34724), .C(out_r[23]), .D(\result_r[28] [15]), 
         .Z(result_r_ns_0__15__N_3[63])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10161_3_lut_4_lut.init = 16'hf780;
    LUT4 i6329_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[23]), .D(\result_i[30] [15]), 
         .Z(result_i_ns_0__15__N_517[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6329_3_lut_4_lut.init = 16'hf780;
    LUT4 i6337_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[22]), .D(\result_i[30] [14]), 
         .Z(result_i_ns_0__15__N_517[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6337_3_lut_4_lut.init = 16'hf780;
    LUT4 i6345_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[21]), .D(\result_i[30] [13]), 
         .Z(result_i_ns_0__15__N_517[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6345_3_lut_4_lut.init = 16'hf780;
    LUT4 i6353_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[20]), .D(\result_i[30] [12]), 
         .Z(result_i_ns_0__15__N_517[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6353_3_lut_4_lut.init = 16'hf780;
    LUT4 i6361_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[19]), .D(\result_i[30] [11]), 
         .Z(result_i_ns_0__15__N_517[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6361_3_lut_4_lut.init = 16'hf780;
    LUT4 i6369_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[18]), .D(\result_i[30] [10]), 
         .Z(result_i_ns_0__15__N_517[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6369_3_lut_4_lut.init = 16'hf780;
    LUT4 i6377_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[17]), .D(\result_i[30] [9]), 
         .Z(result_i_ns_0__15__N_517[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6377_3_lut_4_lut.init = 16'hf780;
    LUT4 i6385_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[16]), .D(\result_i[30] [8]), 
         .Z(result_i_ns_0__15__N_517[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6385_3_lut_4_lut.init = 16'hf780;
    LUT4 i6393_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[15]), .D(\result_i[30] [7]), 
         .Z(result_i_ns_0__15__N_517[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6393_3_lut_4_lut.init = 16'hf780;
    LUT4 i6401_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[14]), .D(\result_i[30] [6]), 
         .Z(result_i_ns_0__15__N_517[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6401_3_lut_4_lut.init = 16'hf780;
    LUT4 i6409_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[13]), .D(\result_i[30] [5]), 
         .Z(result_i_ns_0__15__N_517[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6409_3_lut_4_lut.init = 16'hf780;
    LUT4 i6417_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[12]), .D(\result_i[30] [4]), 
         .Z(result_i_ns_0__15__N_517[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6417_3_lut_4_lut.init = 16'hf780;
    LUT4 i6425_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[11]), .D(\result_i[30] [3]), 
         .Z(result_i_ns_0__15__N_517[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6425_3_lut_4_lut.init = 16'hf780;
    LUT4 i6433_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[10]), .D(\result_i[30] [2]), 
         .Z(result_i_ns_0__15__N_517[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6433_3_lut_4_lut.init = 16'hf780;
    LUT4 i6441_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[9]), .D(\result_i[30] [1]), 
         .Z(result_i_ns_0__15__N_517[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6441_3_lut_4_lut.init = 16'hf780;
    LUT4 i6449_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_i[8]), .D(\result_i[30] [0]), 
         .Z(result_i_ns_0__15__N_517[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6449_3_lut_4_lut.init = 16'hf780;
    LUT4 i10537_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[8]), .D(\result_r[30] [0]), 
         .Z(result_r_ns_0__15__N_3[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10537_3_lut_4_lut.init = 16'hf780;
    LUT4 i10529_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[9]), .D(\result_r[30] [1]), 
         .Z(result_r_ns_0__15__N_3[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10529_3_lut_4_lut.init = 16'hf780;
    LUT4 i10521_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[10]), .D(\result_r[30] [2]), 
         .Z(result_r_ns_0__15__N_3[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10521_3_lut_4_lut.init = 16'hf780;
    LUT4 i10513_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[11]), .D(\result_r[30] [3]), 
         .Z(result_r_ns_0__15__N_3[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10513_3_lut_4_lut.init = 16'hf780;
    LUT4 i10505_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[12]), .D(\result_r[30] [4]), 
         .Z(result_r_ns_0__15__N_3[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10505_3_lut_4_lut.init = 16'hf780;
    LUT4 i10497_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[13]), .D(\result_r[30] [5]), 
         .Z(result_r_ns_0__15__N_3[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10497_3_lut_4_lut.init = 16'hf780;
    LUT4 i10489_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[14]), .D(\result_r[30] [6]), 
         .Z(result_r_ns_0__15__N_3[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10489_3_lut_4_lut.init = 16'hf780;
    LUT4 i10481_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[15]), .D(\result_r[30] [7]), 
         .Z(result_r_ns_0__15__N_3[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10481_3_lut_4_lut.init = 16'hf780;
    LUT4 i10473_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[16]), .D(\result_r[30] [8]), 
         .Z(result_r_ns_0__15__N_3[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10473_3_lut_4_lut.init = 16'hf780;
    LUT4 i10465_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[17]), .D(\result_r[30] [9]), 
         .Z(result_r_ns_0__15__N_3[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10465_3_lut_4_lut.init = 16'hf780;
    LUT4 i10457_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[18]), .D(\result_r[30] [10]), 
         .Z(result_r_ns_0__15__N_3[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10457_3_lut_4_lut.init = 16'hf780;
    LUT4 i10449_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[19]), .D(\result_r[30] [11]), 
         .Z(result_r_ns_0__15__N_3[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10449_3_lut_4_lut.init = 16'hf780;
    LUT4 i10441_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[20]), .D(\result_r[30] [12]), 
         .Z(result_r_ns_0__15__N_3[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10441_3_lut_4_lut.init = 16'hf780;
    LUT4 i10433_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[21]), .D(\result_r[30] [13]), 
         .Z(result_r_ns_0__15__N_3[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10433_3_lut_4_lut.init = 16'hf780;
    LUT4 i10425_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[22]), .D(\result_r[30] [14]), 
         .Z(result_r_ns_0__15__N_3[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10425_3_lut_4_lut.init = 16'hf780;
    LUT4 i10417_3_lut_4_lut (.A(n34712), .B(n32944), .C(out_r[23]), .D(\result_r[30] [15]), 
         .Z(result_r_ns_0__15__N_3[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10417_3_lut_4_lut.init = 16'hf780;
    LUT4 i5945_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[23]), .D(\result_i[27] [15]), 
         .Z(result_i_ns_0__15__N_517[79])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5945_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5953_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[22]), .D(\result_i[27] [14]), 
         .Z(result_i_ns_0__15__N_517[78])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5953_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5961_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[21]), .D(\result_i[27] [13]), 
         .Z(result_i_ns_0__15__N_517[77])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5961_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5969_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[20]), .D(\result_i[27] [12]), 
         .Z(result_i_ns_0__15__N_517[76])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5969_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5977_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[19]), .D(\result_i[27] [11]), 
         .Z(result_i_ns_0__15__N_517[75])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5977_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5985_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[18]), .D(\result_i[27] [10]), 
         .Z(result_i_ns_0__15__N_517[74])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5985_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5993_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[17]), .D(\result_i[27] [9]), 
         .Z(result_i_ns_0__15__N_517[73])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5993_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6001_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[16]), .D(\result_i[27] [8]), 
         .Z(result_i_ns_0__15__N_517[72])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6001_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6009_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[15]), .D(\result_i[27] [7]), 
         .Z(result_i_ns_0__15__N_517[71])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6009_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6017_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[14]), .D(\result_i[27] [6]), 
         .Z(result_i_ns_0__15__N_517[70])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6017_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6025_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[13]), .D(\result_i[27] [5]), 
         .Z(result_i_ns_0__15__N_517[69])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6025_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6033_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[12]), .D(\result_i[27] [4]), 
         .Z(result_i_ns_0__15__N_517[68])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6033_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6041_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[11]), .D(\result_i[27] [3]), 
         .Z(result_i_ns_0__15__N_517[67])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6041_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6049_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[10]), .D(\result_i[27] [2]), 
         .Z(result_i_ns_0__15__N_517[66])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6049_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6057_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[9]), .D(\result_i[27] [1]), 
         .Z(result_i_ns_0__15__N_517[65])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6057_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6065_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_i[8]), .D(\result_i[27] [0]), 
         .Z(result_i_ns_0__15__N_517[64])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6065_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10153_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[8]), .D(\result_r[27] [0]), 
         .Z(result_r_ns_0__15__N_3[64])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10153_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10145_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[9]), .D(\result_r[27] [1]), 
         .Z(result_r_ns_0__15__N_3[65])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10145_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10137_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[10]), .D(\result_r[27] [2]), 
         .Z(result_r_ns_0__15__N_3[66])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10137_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10129_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[11]), .D(\result_r[27] [3]), 
         .Z(result_r_ns_0__15__N_3[67])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10129_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10121_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[12]), .D(\result_r[27] [4]), 
         .Z(result_r_ns_0__15__N_3[68])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10121_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10113_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[13]), .D(\result_r[27] [5]), 
         .Z(result_r_ns_0__15__N_3[69])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10113_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10105_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[14]), .D(\result_r[27] [6]), 
         .Z(result_r_ns_0__15__N_3[70])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10105_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10097_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[15]), .D(\result_r[27] [7]), 
         .Z(result_r_ns_0__15__N_3[71])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10097_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10089_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[16]), .D(\result_r[27] [8]), 
         .Z(result_r_ns_0__15__N_3[72])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10089_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10081_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[17]), .D(\result_r[27] [9]), 
         .Z(result_r_ns_0__15__N_3[73])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10081_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10073_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[18]), .D(\result_r[27] [10]), 
         .Z(result_r_ns_0__15__N_3[74])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10073_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10065_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[19]), .D(\result_r[27] [11]), 
         .Z(result_r_ns_0__15__N_3[75])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10065_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10057_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[20]), .D(\result_r[27] [12]), 
         .Z(result_r_ns_0__15__N_3[76])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10057_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10049_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[21]), .D(\result_r[27] [13]), 
         .Z(result_r_ns_0__15__N_3[77])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10049_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10041_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[22]), .D(\result_r[27] [14]), 
         .Z(result_r_ns_0__15__N_3[78])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10041_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10033_3_lut_4_lut (.A(n34712), .B(n34725), .C(out_r[23]), .D(\result_r[27] [15]), 
         .Z(result_r_ns_0__15__N_3[79])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10033_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5897_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[13]), .D(\result_i[26] [5]), 
         .Z(result_i_ns_0__15__N_517[85])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5897_3_lut_4_lut.init = 16'hf780;
    LUT4 i5905_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[12]), .D(\result_i[26] [4]), 
         .Z(result_i_ns_0__15__N_517[84])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5905_3_lut_4_lut.init = 16'hf780;
    LUT4 i5913_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[11]), .D(\result_i[26] [3]), 
         .Z(result_i_ns_0__15__N_517[83])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5913_3_lut_4_lut.init = 16'hf780;
    LUT4 i5921_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[10]), .D(\result_i[26] [2]), 
         .Z(result_i_ns_0__15__N_517[82])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5921_3_lut_4_lut.init = 16'hf780;
    LUT4 i5929_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[9]), .D(\result_i[26] [1]), 
         .Z(result_i_ns_0__15__N_517[81])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5929_3_lut_4_lut.init = 16'hf780;
    LUT4 i5937_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[8]), .D(\result_i[26] [0]), 
         .Z(result_i_ns_0__15__N_517[80])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5937_3_lut_4_lut.init = 16'hf780;
    LUT4 i5889_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[14]), .D(\result_i[26] [6]), 
         .Z(result_i_ns_0__15__N_517[86])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5889_3_lut_4_lut.init = 16'hf780;
    LUT4 i5881_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[15]), .D(\result_i[26] [7]), 
         .Z(result_i_ns_0__15__N_517[87])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5881_3_lut_4_lut.init = 16'hf780;
    LUT4 i5873_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[16]), .D(\result_i[26] [8]), 
         .Z(result_i_ns_0__15__N_517[88])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5873_3_lut_4_lut.init = 16'hf780;
    LUT4 i5865_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[17]), .D(\result_i[26] [9]), 
         .Z(result_i_ns_0__15__N_517[89])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5865_3_lut_4_lut.init = 16'hf780;
    LUT4 i5857_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[18]), .D(\result_i[26] [10]), 
         .Z(result_i_ns_0__15__N_517[90])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5857_3_lut_4_lut.init = 16'hf780;
    LUT4 i5849_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[19]), .D(\result_i[26] [11]), 
         .Z(result_i_ns_0__15__N_517[91])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5849_3_lut_4_lut.init = 16'hf780;
    LUT4 i5841_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[20]), .D(\result_i[26] [12]), 
         .Z(result_i_ns_0__15__N_517[92])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5841_3_lut_4_lut.init = 16'hf780;
    LUT4 i5833_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[21]), .D(\result_i[26] [13]), 
         .Z(result_i_ns_0__15__N_517[93])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5833_3_lut_4_lut.init = 16'hf780;
    LUT4 i5825_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[22]), .D(\result_i[26] [14]), 
         .Z(result_i_ns_0__15__N_517[94])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5825_3_lut_4_lut.init = 16'hf780;
    LUT4 i5817_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_i[23]), .D(\result_i[26] [15]), 
         .Z(result_i_ns_0__15__N_517[95])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i5817_3_lut_4_lut.init = 16'hf780;
    LUT4 i10025_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[8]), .D(\result_r[26] [0]), 
         .Z(result_r_ns_0__15__N_3[80])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10025_3_lut_4_lut.init = 16'hf780;
    LUT4 i10017_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[9]), .D(\result_r[26] [1]), 
         .Z(result_r_ns_0__15__N_3[81])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10017_3_lut_4_lut.init = 16'hf780;
    LUT4 i10009_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[10]), .D(\result_r[26] [2]), 
         .Z(result_r_ns_0__15__N_3[82])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10009_3_lut_4_lut.init = 16'hf780;
    LUT4 i10001_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[11]), .D(\result_r[26] [3]), 
         .Z(result_r_ns_0__15__N_3[83])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10001_3_lut_4_lut.init = 16'hf780;
    LUT4 i9993_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[12]), .D(\result_r[26] [4]), 
         .Z(result_r_ns_0__15__N_3[84])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9993_3_lut_4_lut.init = 16'hf780;
    LUT4 i9985_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[13]), .D(\result_r[26] [5]), 
         .Z(result_r_ns_0__15__N_3[85])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9985_3_lut_4_lut.init = 16'hf780;
    LUT4 i9977_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[14]), .D(\result_r[26] [6]), 
         .Z(result_r_ns_0__15__N_3[86])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9977_3_lut_4_lut.init = 16'hf780;
    LUT4 i9969_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[15]), .D(\result_r[26] [7]), 
         .Z(result_r_ns_0__15__N_3[87])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9969_3_lut_4_lut.init = 16'hf780;
    LUT4 i9961_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[16]), .D(\result_r[26] [8]), 
         .Z(result_r_ns_0__15__N_3[88])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9961_3_lut_4_lut.init = 16'hf780;
    LUT4 i9953_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[17]), .D(\result_r[26] [9]), 
         .Z(result_r_ns_0__15__N_3[89])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9953_3_lut_4_lut.init = 16'hf780;
    LUT4 i9945_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[18]), .D(\result_r[26] [10]), 
         .Z(result_r_ns_0__15__N_3[90])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9945_3_lut_4_lut.init = 16'hf780;
    LUT4 i9937_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[19]), .D(\result_r[26] [11]), 
         .Z(result_r_ns_0__15__N_3[91])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9937_3_lut_4_lut.init = 16'hf780;
    LUT4 i9929_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[20]), .D(\result_r[26] [12]), 
         .Z(result_r_ns_0__15__N_3[92])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9929_3_lut_4_lut.init = 16'hf780;
    LUT4 i9921_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[21]), .D(\result_r[26] [13]), 
         .Z(result_r_ns_0__15__N_3[93])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9921_3_lut_4_lut.init = 16'hf780;
    LUT4 i9913_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[22]), .D(\result_r[26] [14]), 
         .Z(result_r_ns_0__15__N_3[94])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9913_3_lut_4_lut.init = 16'hf780;
    LUT4 i9905_3_lut_4_lut (.A(n34714), .B(n32944), .C(out_r[23]), .D(\result_r[26] [15]), 
         .Z(result_r_ns_0__15__N_3[95])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i9905_3_lut_4_lut.init = 16'hf780;
    LUT4 i2459_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2459_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10646_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10646_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6457_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6457_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6465_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6465_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6473_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6473_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6481_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6481_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6489_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6489_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6497_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6497_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6505_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6505_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6513_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6513_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6521_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6521_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6529_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6529_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6537_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6537_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6545_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6545_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6553_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6553_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6561_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6561_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6569_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[31] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6569_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10687_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10687_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10675_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10675_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10651_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10651_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10633_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10633_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10625_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10625_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10617_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10617_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10609_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10609_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10601_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10601_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10593_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10593_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10585_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10585_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10577_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10577_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10569_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10569_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10561_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10561_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10553_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10553_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10545_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[31] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i10545_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12804_2_lut_3_lut_4_lut (.A(n34739), .B(n34731), .C(over), .D(n32944), 
         .Z(next_over_N_1081)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i12804_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_341_4_lut (.A(n34740), .B(n34739), .C(n34812), .D(n34811), 
         .Z(n34703)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i1_2_lut_rep_341_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_353_4_lut (.A(n34740), .B(n34739), .C(n34812), .D(n34811), 
         .Z(n34715)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i1_2_lut_rep_353_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_rep_354_4_lut (.A(count_y[2]), .B(n34751), .C(n34802), 
         .D(n34812), .Z(n34716)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A ((C+(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i2_2_lut_rep_354_4_lut.init = 16'hff59;
    LUT4 i12793_2_lut_4_lut (.A(count_y[2]), .B(n34751), .C(n34802), .D(n34812), 
         .Z(n30503)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A !((C+!(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i12793_2_lut_4_lut.init = 16'ha600;
    LUT4 i12783_2_lut_rep_358_4_lut (.A(count_y[2]), .B(n34751), .C(n34802), 
         .D(n34812), .Z(n34720)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i12783_2_lut_rep_358_4_lut.init = 16'hffa6;
    LUT4 i2_2_lut_rep_355_4_lut (.A(count_y[2]), .B(n34751), .C(n34802), 
         .D(n34812), .Z(n34717)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A !(B (C (D))+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i2_2_lut_rep_355_4_lut.init = 16'ha6ff;
    LUT4 i2_2_lut_4_lut (.A(count_y[2]), .B(n34751), .C(n34802), .D(n34812), 
         .Z(n6)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A ((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i2_2_lut_4_lut.init = 16'h00a6;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34706)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B+(C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'hf6ff;
    LUT4 i1_2_lut_rep_352_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34739), 
         .D(n34812), .Z(n34714)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_352_3_lut_4_lut.init = 16'h0600;
    LUT4 i1_2_lut_rep_350_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34739), 
         .D(n34812), .Z(n34712)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_350_3_lut_4_lut.init = 16'h6000;
    LUT4 i1_2_lut_rep_349_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34711)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_349_3_lut_4_lut.init = 16'h6000;
    LUT4 i1_2_lut_rep_348_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34710)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_348_3_lut_4_lut.init = 16'h0600;
    LUT4 i1_2_lut_rep_347_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34709)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_347_3_lut_4_lut.init = 16'h0060;
    LUT4 i1_2_lut_rep_346_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34708)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_346_3_lut_4_lut.init = 16'h0006;
    LUT4 i1_2_lut_rep_345_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34707)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+!(C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_345_3_lut_4_lut.init = 16'h6fff;
    LUT4 i1_2_lut_rep_343_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34705)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B+((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_343_3_lut_4_lut.init = 16'hff6f;
    LUT4 i1_2_lut_rep_342_3_lut_4_lut (.A(count_y[0]), .B(n34751), .C(n34811), 
         .D(n34741), .Z(n34704)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_342_3_lut_4_lut.init = 16'hfff6;
    LUT4 i856_3_lut_rep_377_4_lut (.A(count_y[3]), .B(n34771), .C(n34802), 
         .D(count_y[2]), .Z(n34739)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i856_3_lut_rep_377_4_lut.init = 16'hf10e;
    LUT4 i15498_3_lut (.A(\result_r[10] [12]), .B(\result_r[11] [12]), .C(y_1_delay[0]), 
         .Z(n33882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15498_3_lut.init = 16'hcaca;
    LUT4 i15658_3_lut (.A(\result_r[20] [7]), .B(\result_r[21] [7]), .C(y_1_delay[0]), 
         .Z(n34042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15658_3_lut.init = 16'hcaca;
    LUT4 i15497_3_lut (.A(\result_r[8] [12]), .B(\result_r[9] [12]), .C(y_1_delay[0]), 
         .Z(n33881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15497_3_lut.init = 16'hcaca;
    LUT4 i15648_3_lut (.A(\result_r[0] [7]), .B(\result_r[1] [7]), .C(y_1_delay[0]), 
         .Z(n34032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15648_3_lut.init = 16'hcaca;
    LUT4 i15496_3_lut (.A(\result_r[6] [12]), .B(\result_r[7] [12]), .C(y_1_delay[0]), 
         .Z(n33880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15496_3_lut.init = 16'hcaca;
    LUT4 i15495_3_lut (.A(\result_r[4] [12]), .B(\result_r[5] [12]), .C(y_1_delay[0]), 
         .Z(n33879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15495_3_lut.init = 16'hcaca;
    LUT4 i15494_3_lut (.A(\result_r[2] [12]), .B(\result_r[3] [12]), .C(y_1_delay[0]), 
         .Z(n33878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15494_3_lut.init = 16'hcaca;
    LUT4 i15493_3_lut (.A(\result_r[0] [12]), .B(\result_r[1] [12]), .C(y_1_delay[0]), 
         .Z(n33877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15493_3_lut.init = 16'hcaca;
    LUT4 i15756_3_lut (.A(\result_r[30] [4]), .B(\result_r[31] [4]), .C(y_1_delay[0]), 
         .Z(n34140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15756_3_lut.init = 16'hcaca;
    LUT4 i15755_3_lut (.A(\result_r[28] [4]), .B(\result_r[29] [4]), .C(y_1_delay[0]), 
         .Z(n34139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15755_3_lut.init = 16'hcaca;
    LUT4 i15754_3_lut (.A(\result_r[26] [4]), .B(\result_r[27] [4]), .C(y_1_delay[0]), 
         .Z(n34138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15754_3_lut.init = 16'hcaca;
    LUT4 i15753_3_lut (.A(\result_r[24] [4]), .B(\result_r[25] [4]), .C(y_1_delay[0]), 
         .Z(n34137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15753_3_lut.init = 16'hcaca;
    radix2_U2 radix_no2 (.op_r_23__N_1106({op_r_23__N_1106_adj_7319}), .n34842(n34842), 
            .n3(n3), .shift_4_dout_r({shift_4_dout_r}), .n7431({n7432, 
            n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, 
            n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, 
            n7449, n7450, n7451, n7452, n7453, n7454, n7455}), 
            .n6514(n6514), .\op_r_23__N_1082[29] (op_r_23__N_1082_adj_7378[29]), 
            .n31429(n31429), .op_i_23__N_1154({op_i_23__N_1154_adj_7320}), 
            .shift_4_dout_i({shift_4_dout_i}), .n7590({n7591, n7592, n7593, 
            n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, 
            n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, 
            n7610, n7611, n7612, n7613, n7614}), .\op_i_23__N_1130[26] (op_i_23__N_1130_adj_7381[26]), 
            .n31484(n31484), .GND_net(GND_net), .\op_i_23__N_1310[0] (op_i_23__N_1310_adj_7329[0]), 
            .\op_i_23__N_1310[1] (op_i_23__N_1310_adj_7329[1]), .\op_i_23__N_1310[2] (op_i_23__N_1310_adj_7329[2]), 
            .\op_i_23__N_1310[3] (op_i_23__N_1310_adj_7329[3]), .\op_i_23__N_1310[4] (op_i_23__N_1310_adj_7329[4]), 
            .\op_i_23__N_1310[5] (op_i_23__N_1310_adj_7329[5]), .n89(n89), 
            .n88(n88), .n87(n87), .n86(n86), .n85(n85), .n84(n84), 
            .n83(n83), .n82(n82), .n81(n81), .n80(n80), .n79(n79), 
            .n78(n78), .n77(n77), .n76(n76), .n75(n75), .n74(n74), 
            .n73(n73), .n72(n72), .n71(n71), .n70(n70), .n69(n69), 
            .n68(n68), .n67(n67), .n66(n66), .n65(n65_adj_6358), .VCC_net(VCC_net), 
            .\rom8_w_i[12] (rom8_w_i[12]), .n11148(n11148), .n11149(n11149), 
            .n11150(n11150), .n11151(n11151), .n11152(n11152), .n11153(n11153), 
            .\op_i_23__N_1130[27] (op_i_23__N_1130_adj_7381[27]), .n31482(n31482), 
            .\rom8_w_i[0] (rom8_w_i[0]), .\rom8_w_i[1] (rom8_w_i[1]), .\rom8_w_i[2] (rom8_w_i[2]), 
            .\rom8_w_i[3] (rom8_w_i[3]), .\rom8_w_i[4] (rom8_w_i[4]), .\rom8_w_i[6] (rom8_w_i[6]), 
            .\op_r_23__N_1082[26] (op_r_23__N_1082_adj_7378[26]), .n31435(n31435), 
            .\op_r_23__N_1082[27] (op_r_23__N_1082_adj_7378[27]), .n31433(n31433), 
            .shift_8_dout_i({shift_8_dout_i}), .n119(n119), .\op_r_23__N_1268[0] (op_r_23__N_1268_adj_7324[0]), 
            .\op_r_23__N_1268[1] (op_r_23__N_1268_adj_7324[1]), .\op_r_23__N_1268[2] (op_r_23__N_1268_adj_7324[2]), 
            .\op_r_23__N_1268[3] (op_r_23__N_1268_adj_7324[3]), .\op_r_23__N_1268[4] (op_r_23__N_1268_adj_7324[4]), 
            .\op_r_23__N_1268[5] (op_r_23__N_1268_adj_7324[5]), .\op_r_23__N_1268[6] (op_r_23__N_1268_adj_7324[6]), 
            .\op_r_23__N_1268[7] (op_r_23__N_1268_adj_7324[7]), .\op_r_23__N_1268[8] (op_r_23__N_1268_adj_7324[8]), 
            .\op_r_23__N_1268[9] (op_r_23__N_1268_adj_7324[9]), .\op_r_23__N_1268[10] (op_r_23__N_1268_adj_7324[10]), 
            .\op_r_23__N_1268[11] (op_r_23__N_1268_adj_7324[11]), .\op_r_23__N_1268[12] (op_r_23__N_1268_adj_7324[12]), 
            .\op_r_23__N_1268[13] (op_r_23__N_1268_adj_7324[13]), .\op_r_23__N_1268[14] (op_r_23__N_1268_adj_7324[14]), 
            .\op_r_23__N_1268[15] (op_r_23__N_1268_adj_7324[15]), .\op_r_23__N_1268[16] (op_r_23__N_1268_adj_7324[16]), 
            .\op_r_23__N_1268[17] (op_r_23__N_1268_adj_7324[17]), .\op_r_23__N_1268[18] (op_r_23__N_1268_adj_7324[18]), 
            .\op_r_23__N_1268[19] (op_r_23__N_1268_adj_7324[19]), .\op_r_23__N_1268[20] (op_r_23__N_1268_adj_7324[20]), 
            .\op_r_23__N_1268[21] (op_r_23__N_1268_adj_7324[21]), .\op_r_23__N_1268[22] (op_r_23__N_1268_adj_7324[22]), 
            .\op_r_23__N_1268[23] (op_r_23__N_1268_adj_7324[23]), .\op_r_23__N_1268[24] (op_r_23__N_1268_adj_7324[24]), 
            .\op_r_23__N_1268[25] (op_r_23__N_1268_adj_7324[25]), .\op_r_23__N_1268[26] (op_r_23__N_1268_adj_7324[26]), 
            .\op_r_23__N_1268[27] (op_r_23__N_1268_adj_7324[27]), .\op_r_23__N_1268[28] (op_r_23__N_1268_adj_7324[28]), 
            .\op_r_23__N_1268[29] (op_r_23__N_1268_adj_7324[29]), .\op_r_23__N_1268[30] (op_r_23__N_1268_adj_7324[30]), 
            .\op_r_23__N_1268[31] (op_r_23__N_1268_adj_7324[31]), .\op_r_23__N_1226[0] (op_r_23__N_1226_adj_7326[0]), 
            .\op_r_23__N_1226[1] (op_r_23__N_1226_adj_7326[1]), .\op_r_23__N_1226[2] (op_r_23__N_1226_adj_7326[2]), 
            .\op_r_23__N_1226[3] (op_r_23__N_1226_adj_7326[3]), .\op_r_23__N_1226[4] (op_r_23__N_1226_adj_7326[4]), 
            .\op_r_23__N_1226[5] (op_r_23__N_1226_adj_7326[5]), .\op_r_23__N_1226[6] (op_r_23__N_1226_adj_7326[6]), 
            .\op_r_23__N_1226[7] (op_r_23__N_1226_adj_7326[7]), .\op_r_23__N_1226[8] (op_r_23__N_1226_adj_7326[8]), 
            .\op_r_23__N_1226[9] (op_r_23__N_1226_adj_7326[9]), .\op_r_23__N_1226[10] (op_r_23__N_1226_adj_7326[10]), 
            .\op_r_23__N_1226[11] (op_r_23__N_1226_adj_7326[11]), .\op_r_23__N_1226[12] (op_r_23__N_1226_adj_7326[12]), 
            .\op_r_23__N_1226[13] (op_r_23__N_1226_adj_7326[13]), .\op_r_23__N_1226[14] (op_r_23__N_1226_adj_7326[14]), 
            .\op_r_23__N_1226[15] (op_r_23__N_1226_adj_7326[15]), .\op_r_23__N_1226[16] (op_r_23__N_1226_adj_7326[16]), 
            .\op_r_23__N_1226[17] (op_r_23__N_1226_adj_7326[17]), .\op_r_23__N_1226[18] (op_r_23__N_1226_adj_7326[18]), 
            .\op_r_23__N_1226[19] (op_r_23__N_1226_adj_7326[19]), .\op_r_23__N_1226[20] (op_r_23__N_1226_adj_7326[20]), 
            .\op_r_23__N_1226[21] (op_r_23__N_1226_adj_7326[21]), .\op_r_23__N_1226[22] (op_r_23__N_1226_adj_7326[22]), 
            .\op_r_23__N_1226[23] (op_r_23__N_1226_adj_7326[23]), .\op_r_23__N_1226[24] (op_r_23__N_1226_adj_7326[24]), 
            .\op_r_23__N_1226[25] (op_r_23__N_1226_adj_7326[25]), .\op_r_23__N_1226[26] (op_r_23__N_1226_adj_7326[26]), 
            .\op_r_23__N_1226[27] (op_r_23__N_1226_adj_7326[27]), .\op_r_23__N_1226[28] (op_r_23__N_1226_adj_7326[28]), 
            .\op_r_23__N_1226[29] (op_r_23__N_1226_adj_7326[29]), .\op_r_23__N_1226[30] (op_r_23__N_1226_adj_7326[30]), 
            .\op_r_23__N_1226[31] (op_r_23__N_1226_adj_7326[31]), .\op_i_23__N_1130[24] (op_i_23__N_1130_adj_7381[24]), 
            .n31488(n31488), .\rom8_w_r[0] (rom8_w_r[0]), .\rom8_w_r[1] (rom8_w_r[1]), 
            .\rom8_w_r[7] (rom8_w_r[7]), .\rom8_w_r[3] (rom8_w_r[3]), .\rom8_w_r[4] (rom8_w_r[4]), 
            .\rom8_w_r[5] (rom8_w_r[5]), .\rom8_w_r[6] (rom8_w_r[6]), .\rom8_w_r[8] (rom8_w_r[8]), 
            .\rom8_w_r[10] (rom8_w_r[10]), .n12270(n12270), .n12271(n12271), 
            .n12272(n12272), .n12273(n12273), .n12274(n12274), .n12275(n12275), 
            .n12276(n12276), .n12277(n12277), .n12278(n12278), .n12279(n12279), 
            .n12280(n12280), .n12281(n12281), .n12282(n12282), .n12283(n12283), 
            .n12284(n12284), .n12285(n12285), .n12286(n12286), .n12287(n12287), 
            .n8721(n8721), .n8720(n8720), .n8719(n8719), .n8718(n8718), 
            .n8717(n8717), .n8716(n8716), .n8715(n8715), .n8714(n8714), 
            .n8713(n8713), .n8712(n8712), .n8711(n8711), .n8710(n8710), 
            .n8709(n8709), .n8708(n8708), .n8707(n8707), .n8706(n8706), 
            .n8705(n8705), .n8704(n8704), .n8703(n8703), .n8702(n8702), 
            .n8701(n8701), .n8700(n8700), .n8699(n8699), .n8698(n8698), 
            .n8697(n8697), .n8696(n8696), .n319(n319_adj_6495), .n11154(n11154), 
            .n11155(n11155), .n11156(n11156), .n11157(n11157), .n11158(n11158), 
            .n11159(n11159), .n11160(n11160), .n11161(n11161), .n11162(n11162), 
            .n11163(n11163), .n11164(n11164), .n11165(n11165), .n11166(n11166), 
            .n11167(n11167), .n11168(n11168), .n11169(n11169), .n11170(n11170), 
            .n11171(n11171), .n12444(n12444), .n12445(n12445), .n12446(n12446), 
            .n12447(n12447), .n12448(n12448), .n12449(n12449), .n12450(n12450), 
            .n12451(n12451), .n12452(n12452), .n12453(n12453), .n12288(n12288), 
            .n12289(n12289), .n12290(n12290), .n12291(n12291), .n12292(n12292), 
            .n12293(n12293), .n12294(n12294), .\op_i_23__N_1130[25] (op_i_23__N_1130_adj_7381[25]), 
            .n31486(n31486), .\op_r_23__N_1082[24] (op_r_23__N_1082_adj_7378[24]), 
            .n31439(n31439), .\op_r_23__N_1082[25] (op_r_23__N_1082_adj_7378[25]), 
            .n31437(n31437), .\op_i_23__N_1130[22] (op_i_23__N_1130_adj_7381[22]), 
            .n31492(n31492), .\op_i_23__N_1130[23] (op_i_23__N_1130_adj_7381[23]), 
            .n31490(n31490), .\op_r_23__N_1082[22] (op_r_23__N_1082_adj_7378[22]), 
            .n31443(n31443), .\op_r_23__N_1082[23] (op_r_23__N_1082_adj_7378[23]), 
            .n31441(n31441), .\op_i_23__N_1130[20] (op_i_23__N_1130_adj_7381[20]), 
            .n31496(n31496), .\op_i_23__N_1130[21] (op_i_23__N_1130_adj_7381[21]), 
            .n31494(n31494), .\op_r_23__N_1082[20] (op_r_23__N_1082_adj_7378[20]), 
            .n31447(n31447), .\op_r_23__N_1082[21] (op_r_23__N_1082_adj_7378[21]), 
            .n31445(n31445), .\op_i_23__N_1130[18] (op_i_23__N_1130_adj_7381[18]), 
            .n31500(n31500), .\op_i_23__N_1130[19] (op_i_23__N_1130_adj_7381[19]), 
            .n31498(n31498), .\op_r_23__N_1082[18] (op_r_23__N_1082_adj_7378[18]), 
            .n31451(n31451), .\op_r_23__N_1082[19] (op_r_23__N_1082_adj_7378[19]), 
            .n31449(n31449), .\op_i_23__N_1130[16] (op_i_23__N_1130_adj_7381[16]), 
            .n31504(n31504), .\op_i_23__N_1130[17] (op_i_23__N_1130_adj_7381[17]), 
            .n31502(n31502), .\op_i_23__N_1130[31] (op_i_23__N_1130_adj_7381[31]), 
            .n31474(n31474), .\op_r_23__N_1082[16] (op_r_23__N_1082_adj_7378[16]), 
            .n31455(n31455), .\op_r_23__N_1082[17] (op_r_23__N_1082_adj_7378[17]), 
            .n31453(n31453), .\op_r_23__N_1082[30] (op_r_23__N_1082_adj_7378[30]), 
            .n31427(n31427), .\op_i_23__N_1130[30] (op_i_23__N_1130_adj_7381[30]), 
            .n31476(n31476), .\op_r_23__N_1082[31] (op_r_23__N_1082_adj_7378[31]), 
            .n31425(n31425), .\rom8_state[0] (rom8_state[0]), .n34794(n34794), 
            .\radix_no1_op_i[1] (radix_no1_op_i[1]), .n7507(n7507), .\radix_no1_op_i[0] (radix_no1_op_i[0]), 
            .n7508(n7508), .\radix_no1_op_i[3] (radix_no1_op_i[3]), .n7505(n7505), 
            .\radix_no1_op_i[2] (radix_no1_op_i[2]), .n7506(n7506), .\radix_no1_op_i[5] (radix_no1_op_i[5]), 
            .n7503(n7503), .\radix_no1_op_i[4] (radix_no1_op_i[4]), .n7504(n7504), 
            .\radix_no1_op_i[7] (radix_no1_op_i[7]), .n7501(n7501), .\radix_no1_op_i[6] (radix_no1_op_i[6]), 
            .n7502(n7502), .\radix_no1_op_r[1] (radix_no1_op_r[1]), .\shift_8_dout_r[1] (shift_8_dout_r[1]), 
            .n7560(n7560), .\radix_no1_op_r[0] (radix_no1_op_r[0]), .\shift_8_dout_r[0] (shift_8_dout_r[0]), 
            .n7561(n7561), .\radix_no1_op_r[3] (radix_no1_op_r[3]), .\shift_8_dout_r[3] (shift_8_dout_r[3]), 
            .n7558(n7558), .\radix_no1_op_r[2] (radix_no1_op_r[2]), .\shift_8_dout_r[2] (shift_8_dout_r[2]), 
            .n7559(n7559), .\radix_no1_op_r[5] (radix_no1_op_r[5]), .\shift_8_dout_r[5] (shift_8_dout_r[5]), 
            .n7556(n7556), .\radix_no1_op_r[4] (radix_no1_op_r[4]), .\shift_8_dout_r[4] (shift_8_dout_r[4]), 
            .n7557(n7557), .\radix_no1_op_r[7] (radix_no1_op_r[7]), .\shift_8_dout_r[7] (shift_8_dout_r[7]), 
            .n7554(n7554), .\radix_no1_op_r[6] (radix_no1_op_r[6]), .\shift_8_dout_r[6] (shift_8_dout_r[6]), 
            .n7555(n7555), .\op_i_23__N_1130[8] (op_i_23__N_1130_adj_7330[8]), 
            .n31422(n31422), .\op_i_23__N_1130[9] (op_i_23__N_1130_adj_7330[9]), 
            .n31420(n31420), .\op_i_23__N_1130[13] (op_i_23__N_1130_adj_7330[13]), 
            .n31412(n31412), .\op_i_23__N_1130[10] (op_i_23__N_1130_adj_7330[10]), 
            .n31418(n31418), .\op_i_23__N_1130[11] (op_i_23__N_1130_adj_7330[11]), 
            .n31416(n31416), .\op_i_23__N_1130[14] (op_i_23__N_1130_adj_7330[14]), 
            .n31410(n31410), .\op_i_23__N_1130[15] (op_i_23__N_1130_adj_7330[15]), 
            .n31408(n31408), .\op_i_23__N_1130[12] (op_i_23__N_1130_adj_7330[12]), 
            .n31414(n31414), .\op_r_23__N_1082[14] (op_r_23__N_1082_adj_7327[14]), 
            .n31606(n31606), .\op_r_23__N_1082[15] (op_r_23__N_1082_adj_7327[15]), 
            .n31604(n31604), .\op_r_23__N_1082[12] (op_r_23__N_1082_adj_7327[12]), 
            .n31610(n31610), .\op_r_23__N_1082[13] (op_r_23__N_1082_adj_7327[13]), 
            .n31608(n31608), .\op_r_23__N_1082[10] (op_r_23__N_1082_adj_7327[10]), 
            .n31614(n31614), .\op_r_23__N_1082[11] (op_r_23__N_1082_adj_7327[11]), 
            .n31612(n31612), .\op_r_23__N_1082[8] (op_r_23__N_1082_adj_7327[8]), 
            .n31618(n31618), .\op_r_23__N_1082[9] (op_r_23__N_1082_adj_7327[9]), 
            .n31616(n31616), .n34625(n34625), .n34620(n34620), .n34619(n34619), 
            .n34614(n34614), .n34613(n34613), .n34608(n34608), .n34607(n34607), 
            .n34606(n34606), .n34605(n34605), .n34600(n34600), .n34599(n34599), 
            .n34598(n34598), .n34597(n34597), .n34592(n34592), .n34591(n34591), 
            .n34590(n34590), .n34589(n34589), .n34626(n34626), .n34631(n34631), 
            .n34632(n34632), .n34637(n34637), .n34638(n34638), .n34643(n34643), 
            .n34644(n34644), .n34647(n34647), .n34648(n34648), .n34653(n34653), 
            .n34654(n34654), .n34657(n34657), .n34658(n34658), .n34663(n34663), 
            .n34664(n34664), .n34681(n34681), .n34682(n34682), .n34687(n34687), 
            .n34688(n34688), .n34691(n34691), .n34692(n34692), .n34693(n34693), 
            .n34694(n34694), .n34695(n34695), .n34696(n34696), .n34697(n34697), 
            .n34698(n34698), .n34699(n34699), .n34700(n34700), .n34701(n34701), 
            .n34702(n34702), .valid(valid_adj_6771), .clk_c_enable_1373(clk_c_enable_1373), 
            .\op_i_23__N_1130[14]_adj_70 (op_i_23__N_1130_adj_7381[14]), .n31508(n31508), 
            .\op_i_23__N_1130[15]_adj_71 (op_i_23__N_1130_adj_7381[15]), .n31506(n31506), 
            .\op_r_23__N_1082[14]_adj_72 (op_r_23__N_1082_adj_7378[14]), .n31459(n31459), 
            .\op_r_23__N_1082[15]_adj_73 (op_r_23__N_1082_adj_7378[15]), .n31457(n31457), 
            .\op_i_23__N_1130[13]_adj_74 (op_i_23__N_1130_adj_7381[13]), .n31510(n31510), 
            .\op_r_23__N_1082[12]_adj_75 (op_r_23__N_1082_adj_7378[12]), .n31463(n31463), 
            .\op_r_23__N_1082[13]_adj_76 (op_r_23__N_1082_adj_7378[13]), .n31461(n31461), 
            .\op_i_23__N_1130[12]_adj_77 (op_i_23__N_1130_adj_7381[12]), .n31512(n31512), 
            .\op_r_23__N_1082[28] (op_r_23__N_1082_adj_7378[28]), .n31431(n31431), 
            .\op_r_23__N_1082[10]_adj_78 (op_r_23__N_1082_adj_7378[10]), .n31467(n31467), 
            .\op_r_23__N_1082[11]_adj_79 (op_r_23__N_1082_adj_7378[11]), .n31465(n31465), 
            .\op_i_23__N_1130[10]_adj_80 (op_i_23__N_1130_adj_7381[10]), .n31516(n31516), 
            .\op_i_23__N_1130[11]_adj_81 (op_i_23__N_1130_adj_7381[11]), .n31514(n31514), 
            .\op_r_23__N_1082[8]_adj_82 (op_r_23__N_1082_adj_7378[8]), .n31471(n31471), 
            .\op_r_23__N_1082[9]_adj_83 (op_r_23__N_1082_adj_7378[9]), .n31469(n31469), 
            .\op_i_23__N_1130[8]_adj_84 (op_i_23__N_1130_adj_7381[8]), .n31520(n31520), 
            .\op_i_23__N_1130[9]_adj_85 (op_i_23__N_1130_adj_7381[9]), .n31518(n31518), 
            .\op_i_23__N_1130[29] (op_i_23__N_1130_adj_7381[29]), .n31478(n31478), 
            .\op_i_23__N_1130[28] (op_i_23__N_1130_adj_7381[28]), .n31480(n31480)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(115[8] 128[2])
    LUT4 i863_3_lut_rep_379_3_lut_4_lut (.A(count_y[2]), .B(n34802), .C(n34771), 
         .D(count_y[3]), .Z(n34741)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i863_3_lut_rep_379_3_lut_4_lut.init = 16'hee10;
    LUT4 i1_2_lut_rep_409 (.A(count_y[0]), .B(n32925), .Z(n34771)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_409.init = 16'heeee;
    LUT4 i1_2_lut_rep_389_3_lut (.A(count_y[0]), .B(n32925), .C(count_y[3]), 
         .Z(n34751)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_389_3_lut.init = 16'hfefe;
    LUT4 i841_2_lut_rep_378_3_lut_3_lut (.A(count_y[0]), .B(n32925), .C(count_y[3]), 
         .Z(n34740)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i841_2_lut_rep_378_3_lut_3_lut.init = 16'h5454;
    LUT4 i15167_3_lut (.A(\result_i[30] [8]), .B(\result_i[31] [8]), .C(y_1_delay[0]), 
         .Z(n33551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15167_3_lut.init = 16'hcaca;
    LUT4 i15166_3_lut (.A(\result_i[28] [8]), .B(\result_i[29] [8]), .C(y_1_delay[0]), 
         .Z(n33550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15166_3_lut.init = 16'hcaca;
    LUT4 i15752_3_lut (.A(\result_r[22] [4]), .B(\result_r[23] [4]), .C(y_1_delay[0]), 
         .Z(n34136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15752_3_lut.init = 16'hcaca;
    LUT4 i15751_3_lut (.A(\result_r[20] [4]), .B(\result_r[21] [4]), .C(y_1_delay[0]), 
         .Z(n34135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15751_3_lut.init = 16'hcaca;
    LUT4 i15657_3_lut (.A(\result_r[18] [7]), .B(\result_r[19] [7]), .C(y_1_delay[0]), 
         .Z(n34041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15657_3_lut.init = 16'hcaca;
    LUT4 i15477_3_lut (.A(\result_r[30] [13]), .B(\result_r[31] [13]), .C(y_1_delay[0]), 
         .Z(n33861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15477_3_lut.init = 16'hcaca;
    LUT4 i15476_3_lut (.A(\result_r[28] [13]), .B(\result_r[29] [13]), .C(y_1_delay[0]), 
         .Z(n33860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15476_3_lut.init = 16'hcaca;
    LUT4 i15656_3_lut (.A(\result_r[16] [7]), .B(\result_r[17] [7]), .C(y_1_delay[0]), 
         .Z(n34040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15656_3_lut.init = 16'hcaca;
    LUT4 i15475_3_lut (.A(\result_r[26] [13]), .B(\result_r[27] [13]), .C(y_1_delay[0]), 
         .Z(n33859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15475_3_lut.init = 16'hcaca;
    LUT4 i15593_3_lut (.A(\result_r[14] [9]), .B(\result_r[15] [9]), .C(y_1_delay[0]), 
         .Z(n33977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15593_3_lut.init = 16'hcaca;
    LUT4 i6825_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[480])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6825_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6817_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[481])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6817_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15725_3_lut (.A(\result_r[30] [5]), .B(\result_r[31] [5]), .C(y_1_delay[0]), 
         .Z(n34109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15725_3_lut.init = 16'hcaca;
    LUT4 i15724_3_lut (.A(\result_r[28] [5]), .B(\result_r[29] [5]), .C(y_1_delay[0]), 
         .Z(n34108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15724_3_lut.init = 16'hcaca;
    LUT4 i6809_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[482])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6809_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i14945_3_lut (.A(\result_i[20] [15]), .B(\result_i[21] [15]), .C(y_1_delay[0]), 
         .Z(n33329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14945_3_lut.init = 16'hcaca;
    LUT4 i6801_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[483])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6801_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15474_3_lut (.A(\result_r[24] [13]), .B(\result_r[25] [13]), .C(y_1_delay[0]), 
         .Z(n33858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15474_3_lut.init = 16'hcaca;
    LUT4 i15750_3_lut (.A(\result_r[18] [4]), .B(\result_r[19] [4]), .C(y_1_delay[0]), 
         .Z(n34134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15750_3_lut.init = 16'hcaca;
    LUT4 i15749_3_lut (.A(\result_r[16] [4]), .B(\result_r[17] [4]), .C(y_1_delay[0]), 
         .Z(n34133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15749_3_lut.init = 16'hcaca;
    LUT4 i15655_3_lut (.A(\result_r[14] [7]), .B(\result_r[15] [7]), .C(y_1_delay[0]), 
         .Z(n34039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15655_3_lut.init = 16'hcaca;
    LUT4 i15473_3_lut (.A(\result_r[22] [13]), .B(\result_r[23] [13]), .C(y_1_delay[0]), 
         .Z(n33857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15473_3_lut.init = 16'hcaca;
    LUT4 i15592_3_lut (.A(\result_r[12] [9]), .B(\result_r[13] [9]), .C(y_1_delay[0]), 
         .Z(n33976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15592_3_lut.init = 16'hcaca;
    LUT4 i15472_3_lut (.A(\result_r[20] [13]), .B(\result_r[21] [13]), .C(y_1_delay[0]), 
         .Z(n33856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15472_3_lut.init = 16'hcaca;
    LUT4 i6793_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[484])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6793_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i6785_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[485])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6785_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15654_3_lut (.A(\result_r[12] [7]), .B(\result_r[13] [7]), .C(y_1_delay[0]), 
         .Z(n34038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15654_3_lut.init = 16'hcaca;
    LUT4 i15471_3_lut (.A(\result_r[18] [13]), .B(\result_r[19] [13]), .C(y_1_delay[0]), 
         .Z(n33855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15471_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_361_4_lut_4_lut_4_lut (.A(count_y[4]), .B(n34771), 
         .C(n34770), .D(count_y[3]), .Z(n34723)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_361_4_lut_4_lut_4_lut.init = 16'h5008;
    LUT4 i1_2_lut_rep_362_4_lut_4_lut_4_lut (.A(count_y[4]), .B(n34771), 
         .C(n34770), .D(count_y[3]), .Z(n34724)) /* synthesis lut_function=(!((B (C (D)+!C !(D))+!B (C (D)))+!A)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i1_2_lut_rep_362_4_lut_4_lut_4_lut.init = 16'h0aa2;
    LUT4 i15134_3_lut (.A(\result_i[26] [9]), .B(\result_i[27] [9]), .C(y_1_delay[0]), 
         .Z(n33518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15134_3_lut.init = 16'hcaca;
    LUT4 i15133_3_lut (.A(\result_i[24] [9]), .B(\result_i[25] [9]), .C(y_1_delay[0]), 
         .Z(n33517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15133_3_lut.init = 16'hcaca;
    LUT4 i15470_3_lut (.A(\result_r[16] [13]), .B(\result_r[17] [13]), .C(y_1_delay[0]), 
         .Z(n33854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15470_3_lut.init = 16'hcaca;
    LUT4 i12791_2_lut_rep_363_4_lut_4_lut_4_lut (.A(count_y[4]), .B(n34771), 
         .C(n34770), .D(count_y[3]), .Z(n34725)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i12791_2_lut_rep_363_4_lut_4_lut_4_lut.init = 16'hfaae;
    LUT4 i15165_3_lut (.A(\result_i[26] [8]), .B(\result_i[27] [8]), .C(y_1_delay[0]), 
         .Z(n33549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15165_3_lut.init = 16'hcaca;
    LUT4 i15164_3_lut (.A(\result_i[24] [8]), .B(\result_i[25] [8]), .C(y_1_delay[0]), 
         .Z(n33548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15164_3_lut.init = 16'hcaca;
    LUT4 i15748_3_lut (.A(\result_r[14] [4]), .B(\result_r[15] [4]), .C(y_1_delay[0]), 
         .Z(n34132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15748_3_lut.init = 16'hcaca;
    LUT4 i15747_3_lut (.A(\result_r[12] [4]), .B(\result_r[13] [4]), .C(y_1_delay[0]), 
         .Z(n34131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15747_3_lut.init = 16'hcaca;
    LUT4 i15653_3_lut (.A(\result_r[10] [7]), .B(\result_r[11] [7]), .C(y_1_delay[0]), 
         .Z(n34037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15653_3_lut.init = 16'hcaca;
    LUT4 i15132_3_lut (.A(\result_i[22] [9]), .B(\result_i[23] [9]), .C(y_1_delay[0]), 
         .Z(n33516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15132_3_lut.init = 16'hcaca;
    LUT4 i15469_3_lut (.A(\result_r[14] [13]), .B(\result_r[15] [13]), .C(y_1_delay[0]), 
         .Z(n33853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15469_3_lut.init = 16'hcaca;
    LUT4 i15468_3_lut (.A(\result_r[12] [13]), .B(\result_r[13] [13]), .C(y_1_delay[0]), 
         .Z(n33852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15468_3_lut.init = 16'hcaca;
    LUT4 i15131_3_lut (.A(\result_i[20] [9]), .B(\result_i[21] [9]), .C(y_1_delay[0]), 
         .Z(n33515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15131_3_lut.init = 16'hcaca;
    LUT4 i15467_3_lut (.A(\result_r[10] [13]), .B(\result_r[11] [13]), .C(y_1_delay[0]), 
         .Z(n33851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15467_3_lut.init = 16'hcaca;
    LUT4 i15466_3_lut (.A(\result_r[8] [13]), .B(\result_r[9] [13]), .C(y_1_delay[0]), 
         .Z(n33850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15466_3_lut.init = 16'hcaca;
    LUT4 i15130_3_lut (.A(\result_i[18] [9]), .B(\result_i[19] [9]), .C(y_1_delay[0]), 
         .Z(n33514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15130_3_lut.init = 16'hcaca;
    LUT4 i15465_3_lut (.A(\result_r[6] [13]), .B(\result_r[7] [13]), .C(y_1_delay[0]), 
         .Z(n33849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15465_3_lut.init = 16'hcaca;
    LUT4 i15464_3_lut (.A(\result_r[4] [13]), .B(\result_r[5] [13]), .C(y_1_delay[0]), 
         .Z(n33848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15464_3_lut.init = 16'hcaca;
    LUT4 i15129_3_lut (.A(\result_i[16] [9]), .B(\result_i[17] [9]), .C(y_1_delay[0]), 
         .Z(n33513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15129_3_lut.init = 16'hcaca;
    LUT4 i15746_3_lut (.A(\result_r[10] [4]), .B(\result_r[11] [4]), .C(y_1_delay[0]), 
         .Z(n34130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15746_3_lut.init = 16'hcaca;
    LUT4 i15745_3_lut (.A(\result_r[8] [4]), .B(\result_r[9] [4]), .C(y_1_delay[0]), 
         .Z(n34129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15745_3_lut.init = 16'hcaca;
    LUT4 i15652_3_lut (.A(\result_r[8] [7]), .B(\result_r[9] [7]), .C(y_1_delay[0]), 
         .Z(n34036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15652_3_lut.init = 16'hcaca;
    LUT4 i15463_3_lut (.A(\result_r[2] [13]), .B(\result_r[3] [13]), .C(y_1_delay[0]), 
         .Z(n33847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15463_3_lut.init = 16'hcaca;
    LUT4 i15128_3_lut (.A(\result_i[14] [9]), .B(\result_i[15] [9]), .C(y_1_delay[0]), 
         .Z(n33512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15128_3_lut.init = 16'hcaca;
    LUT4 i15127_3_lut (.A(\result_i[12] [9]), .B(\result_i[13] [9]), .C(y_1_delay[0]), 
         .Z(n33511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15127_3_lut.init = 16'hcaca;
    LUT4 i15462_3_lut (.A(\result_r[0] [13]), .B(\result_r[1] [13]), .C(y_1_delay[0]), 
         .Z(n33846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15462_3_lut.init = 16'hcaca;
    LUT4 i15163_3_lut (.A(\result_i[22] [8]), .B(\result_i[23] [8]), .C(y_1_delay[0]), 
         .Z(n33547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15163_3_lut.init = 16'hcaca;
    LUT4 i15126_3_lut (.A(\result_i[10] [9]), .B(\result_i[11] [9]), .C(y_1_delay[0]), 
         .Z(n33510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15126_3_lut.init = 16'hcaca;
    LUT4 i15162_3_lut (.A(\result_i[20] [8]), .B(\result_i[21] [8]), .C(y_1_delay[0]), 
         .Z(n33546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15162_3_lut.init = 16'hcaca;
    LUT4 i15651_3_lut (.A(\result_r[6] [7]), .B(\result_r[7] [7]), .C(y_1_delay[0]), 
         .Z(n34035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15651_3_lut.init = 16'hcaca;
    LUT4 i15161_3_lut (.A(\result_i[18] [8]), .B(\result_i[19] [8]), .C(y_1_delay[0]), 
         .Z(n33545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15161_3_lut.init = 16'hcaca;
    LUT4 i15125_3_lut (.A(\result_i[8] [9]), .B(\result_i[9] [9]), .C(y_1_delay[0]), 
         .Z(n33509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15125_3_lut.init = 16'hcaca;
    LUT4 i15160_3_lut (.A(\result_i[16] [8]), .B(\result_i[17] [8]), .C(y_1_delay[0]), 
         .Z(n33544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15160_3_lut.init = 16'hcaca;
    LUT4 i15260_3_lut (.A(\result_i[30] [5]), .B(\result_i[31] [5]), .C(y_1_delay[0]), 
         .Z(n33644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15260_3_lut.init = 16'hcaca;
    LUT4 i15259_3_lut (.A(\result_i[28] [5]), .B(\result_i[29] [5]), .C(y_1_delay[0]), 
         .Z(n33643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15259_3_lut.init = 16'hcaca;
    LUT4 i15258_3_lut (.A(\result_i[26] [5]), .B(\result_i[27] [5]), .C(y_1_delay[0]), 
         .Z(n33642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15258_3_lut.init = 16'hcaca;
    LUT4 i15257_3_lut (.A(\result_i[24] [5]), .B(\result_i[25] [5]), .C(y_1_delay[0]), 
         .Z(n33641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15257_3_lut.init = 16'hcaca;
    LUT4 i15256_3_lut (.A(\result_i[22] [5]), .B(\result_i[23] [5]), .C(y_1_delay[0]), 
         .Z(n33640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15256_3_lut.init = 16'hcaca;
    LUT4 i15255_3_lut (.A(\result_i[20] [5]), .B(\result_i[21] [5]), .C(y_1_delay[0]), 
         .Z(n33639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15255_3_lut.init = 16'hcaca;
    LUT4 i15254_3_lut (.A(\result_i[18] [5]), .B(\result_i[19] [5]), .C(y_1_delay[0]), 
         .Z(n33638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15254_3_lut.init = 16'hcaca;
    LUT4 i15253_3_lut (.A(\result_i[16] [5]), .B(\result_i[17] [5]), .C(y_1_delay[0]), 
         .Z(n33637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15253_3_lut.init = 16'hcaca;
    LUT4 i15252_3_lut (.A(\result_i[14] [5]), .B(\result_i[15] [5]), .C(y_1_delay[0]), 
         .Z(n33636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15252_3_lut.init = 16'hcaca;
    LUT4 i15251_3_lut (.A(\result_i[12] [5]), .B(\result_i[13] [5]), .C(y_1_delay[0]), 
         .Z(n33635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15251_3_lut.init = 16'hcaca;
    LUT4 i15632_3_lut (.A(\result_r[30] [8]), .B(\result_r[31] [8]), .C(y_1_delay[0]), 
         .Z(n34016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15632_3_lut.init = 16'hcaca;
    LUT4 i15631_3_lut (.A(\result_r[28] [8]), .B(\result_r[29] [8]), .C(y_1_delay[0]), 
         .Z(n34015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15631_3_lut.init = 16'hcaca;
    LUT4 i15250_3_lut (.A(\result_i[10] [5]), .B(\result_i[11] [5]), .C(y_1_delay[0]), 
         .Z(n33634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15250_3_lut.init = 16'hcaca;
    LUT4 i15249_3_lut (.A(\result_i[8] [5]), .B(\result_i[9] [5]), .C(y_1_delay[0]), 
         .Z(n33633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15249_3_lut.init = 16'hcaca;
    LUT4 i15248_3_lut (.A(\result_i[6] [5]), .B(\result_i[7] [5]), .C(y_1_delay[0]), 
         .Z(n33632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15248_3_lut.init = 16'hcaca;
    LUT4 i15247_3_lut (.A(\result_i[4] [5]), .B(\result_i[5] [5]), .C(y_1_delay[0]), 
         .Z(n33631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15247_3_lut.init = 16'hcaca;
    LUT4 i15630_3_lut (.A(\result_r[26] [8]), .B(\result_r[27] [8]), .C(y_1_delay[0]), 
         .Z(n34014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15630_3_lut.init = 16'hcaca;
    LUT4 i15629_3_lut (.A(\result_r[24] [8]), .B(\result_r[25] [8]), .C(y_1_delay[0]), 
         .Z(n34013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15629_3_lut.init = 16'hcaca;
    LUT4 i15628_3_lut (.A(\result_r[22] [8]), .B(\result_r[23] [8]), .C(y_1_delay[0]), 
         .Z(n34012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15628_3_lut.init = 16'hcaca;
    LUT4 i15627_3_lut (.A(\result_r[20] [8]), .B(\result_r[21] [8]), .C(y_1_delay[0]), 
         .Z(n34011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15627_3_lut.init = 16'hcaca;
    LUT4 i15626_3_lut (.A(\result_r[18] [8]), .B(\result_r[19] [8]), .C(y_1_delay[0]), 
         .Z(n34010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15626_3_lut.init = 16'hcaca;
    LUT4 i15625_3_lut (.A(\result_r[16] [8]), .B(\result_r[17] [8]), .C(y_1_delay[0]), 
         .Z(n34009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15625_3_lut.init = 16'hcaca;
    LUT4 i15624_3_lut (.A(\result_r[14] [8]), .B(\result_r[15] [8]), .C(y_1_delay[0]), 
         .Z(n34008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15624_3_lut.init = 16'hcaca;
    LUT4 i15623_3_lut (.A(\result_r[12] [8]), .B(\result_r[13] [8]), .C(y_1_delay[0]), 
         .Z(n34007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15623_3_lut.init = 16'hcaca;
    LUT4 i15622_3_lut (.A(\result_r[10] [8]), .B(\result_r[11] [8]), .C(y_1_delay[0]), 
         .Z(n34006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15622_3_lut.init = 16'hcaca;
    LUT4 i15621_3_lut (.A(\result_r[8] [8]), .B(\result_r[9] [8]), .C(y_1_delay[0]), 
         .Z(n34005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15621_3_lut.init = 16'hcaca;
    LUT4 i15620_3_lut (.A(\result_r[6] [8]), .B(\result_r[7] [8]), .C(y_1_delay[0]), 
         .Z(n34004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15620_3_lut.init = 16'hcaca;
    LUT4 i15619_3_lut (.A(\result_r[4] [8]), .B(\result_r[5] [8]), .C(y_1_delay[0]), 
         .Z(n34003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15619_3_lut.init = 16'hcaca;
    FD1P3AX dout_i_i0_i2 (.D(next_dout_i_15__N_1045[1]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_1));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i2.GSR = "ENABLED";
    LUT4 i15246_3_lut (.A(\result_i[2] [5]), .B(\result_i[3] [5]), .C(y_1_delay[0]), 
         .Z(n33630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15246_3_lut.init = 16'hcaca;
    LUT4 i15650_3_lut (.A(\result_r[4] [7]), .B(\result_r[5] [7]), .C(y_1_delay[0]), 
         .Z(n34034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15650_3_lut.init = 16'hcaca;
    LUT4 i15744_3_lut (.A(\result_r[6] [4]), .B(\result_r[7] [4]), .C(y_1_delay[0]), 
         .Z(n34128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15744_3_lut.init = 16'hcaca;
    LUT4 i15245_3_lut (.A(\result_i[0] [5]), .B(\result_i[1] [5]), .C(y_1_delay[0]), 
         .Z(n33629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15245_3_lut.init = 16'hcaca;
    LUT4 i15743_3_lut (.A(\result_r[4] [4]), .B(\result_r[5] [4]), .C(y_1_delay[0]), 
         .Z(n34127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15743_3_lut.init = 16'hcaca;
    LUT4 i15159_3_lut (.A(\result_i[14] [8]), .B(\result_i[15] [8]), .C(y_1_delay[0]), 
         .Z(n33543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15159_3_lut.init = 16'hcaca;
    LUT4 i15618_3_lut (.A(\result_r[2] [8]), .B(\result_r[3] [8]), .C(y_1_delay[0]), 
         .Z(n34002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15618_3_lut.init = 16'hcaca;
    LUT4 i15158_3_lut (.A(\result_i[12] [8]), .B(\result_i[13] [8]), .C(y_1_delay[0]), 
         .Z(n33542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15158_3_lut.init = 16'hcaca;
    LUT4 i15617_3_lut (.A(\result_r[0] [8]), .B(\result_r[1] [8]), .C(y_1_delay[0]), 
         .Z(n34001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15617_3_lut.init = 16'hcaca;
    LUT4 i15157_3_lut (.A(\result_i[10] [8]), .B(\result_i[11] [8]), .C(y_1_delay[0]), 
         .Z(n33541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15157_3_lut.init = 16'hcaca;
    LUT4 i15156_3_lut (.A(\result_i[8] [8]), .B(\result_i[9] [8]), .C(y_1_delay[0]), 
         .Z(n33540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15156_3_lut.init = 16'hcaca;
    LUT4 i15124_3_lut (.A(\result_i[6] [9]), .B(\result_i[7] [9]), .C(y_1_delay[0]), 
         .Z(n33508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15124_3_lut.init = 16'hcaca;
    LUT4 i15742_3_lut (.A(\result_r[2] [4]), .B(\result_r[3] [4]), .C(y_1_delay[0]), 
         .Z(n34126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15742_3_lut.init = 16'hcaca;
    LUT4 i15123_3_lut (.A(\result_i[4] [9]), .B(\result_i[5] [9]), .C(y_1_delay[0]), 
         .Z(n33507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15123_3_lut.init = 16'hcaca;
    LUT4 i15741_3_lut (.A(\result_r[0] [4]), .B(\result_r[1] [4]), .C(y_1_delay[0]), 
         .Z(n34125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15741_3_lut.init = 16'hcaca;
    LUT4 i15043_3_lut (.A(\result_i[30] [12]), .B(\result_i[31] [12]), .C(y_1_delay[0]), 
         .Z(n33427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15043_3_lut.init = 16'hcaca;
    LUT4 i15042_3_lut (.A(\result_i[28] [12]), .B(\result_i[29] [12]), .C(y_1_delay[0]), 
         .Z(n33426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15042_3_lut.init = 16'hcaca;
    LUT4 i15155_3_lut (.A(\result_i[6] [8]), .B(\result_i[7] [8]), .C(y_1_delay[0]), 
         .Z(n33539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15155_3_lut.init = 16'hcaca;
    LUT4 i15154_3_lut (.A(\result_i[4] [8]), .B(\result_i[5] [8]), .C(y_1_delay[0]), 
         .Z(n33538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15154_3_lut.init = 16'hcaca;
    LUT4 i15153_3_lut (.A(\result_i[2] [8]), .B(\result_i[3] [8]), .C(y_1_delay[0]), 
         .Z(n33537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15153_3_lut.init = 16'hcaca;
    LUT4 i15122_3_lut (.A(\result_i[2] [9]), .B(\result_i[3] [9]), .C(y_1_delay[0]), 
         .Z(n33506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15122_3_lut.init = 16'hcaca;
    LUT4 i15152_3_lut (.A(\result_i[0] [8]), .B(\result_i[1] [8]), .C(y_1_delay[0]), 
         .Z(n33536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15152_3_lut.init = 16'hcaca;
    LUT4 i15121_3_lut (.A(\result_i[0] [9]), .B(\result_i[1] [9]), .C(y_1_delay[0]), 
         .Z(n33505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15121_3_lut.init = 16'hcaca;
    LUT4 i15446_3_lut (.A(\result_r[30] [14]), .B(\result_r[31] [14]), .C(y_1_delay[0]), 
         .Z(n33830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15446_3_lut.init = 16'hcaca;
    LUT4 i15445_3_lut (.A(\result_r[28] [14]), .B(\result_r[29] [14]), .C(y_1_delay[0]), 
         .Z(n33829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15445_3_lut.init = 16'hcaca;
    L6MUX21 i14963 (.D0(n33343), .D1(n33344), .SD(y_1_delay[3]), .Z(n33347));
    L6MUX21 i14964 (.D0(n33345), .D1(n33346), .SD(y_1_delay[3]), .Z(n33348));
    L6MUX21 i15335 (.D0(n33715), .D1(n33716), .SD(y_1_delay[3]), .Z(n33719));
    L6MUX21 i15336 (.D0(n33717), .D1(n33718), .SD(y_1_delay[3]), .Z(n33720));
    L6MUX21 i15366 (.D0(n33746), .D1(n33747), .SD(y_1_delay[3]), .Z(n33750));
    L6MUX21 i15367 (.D0(n33748), .D1(n33749), .SD(y_1_delay[3]), .Z(n33751));
    L6MUX21 i15087 (.D0(n33467), .D1(n33468), .SD(y_1_delay[3]), .Z(n33471));
    L6MUX21 i15088 (.D0(n33469), .D1(n33470), .SD(y_1_delay[3]), .Z(n33472));
    LUT4 i15041_3_lut (.A(\result_i[26] [12]), .B(\result_i[27] [12]), .C(y_1_delay[0]), 
         .Z(n33425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15041_3_lut.init = 16'hcaca;
    LUT4 i15444_3_lut (.A(\result_r[26] [14]), .B(\result_r[27] [14]), .C(y_1_delay[0]), 
         .Z(n33828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15444_3_lut.init = 16'hcaca;
    L6MUX21 i14901 (.D0(n33281), .D1(n33282), .SD(y_1_delay[3]), .Z(n33285));
    L6MUX21 i14902 (.D0(n33283), .D1(n33284), .SD(y_1_delay[3]), .Z(n33286));
    L6MUX21 i15707 (.D0(n34087), .D1(n34088), .SD(y_1_delay[3]), .Z(n34091));
    L6MUX21 i15708 (.D0(n34089), .D1(n34090), .SD(y_1_delay[3]), .Z(n34092));
    L6MUX21 i14994 (.D0(n33374), .D1(n33375), .SD(y_1_delay[3]), .Z(n33378));
    L6MUX21 i14995 (.D0(n33376), .D1(n33377), .SD(y_1_delay[3]), .Z(n33379));
    L6MUX21 i15397 (.D0(n33777), .D1(n33778), .SD(y_1_delay[3]), .Z(n33781));
    L6MUX21 i15398 (.D0(n33779), .D1(n33780), .SD(y_1_delay[3]), .Z(n33782));
    L6MUX21 i15428 (.D0(n33808), .D1(n33809), .SD(y_1_delay[3]), .Z(n33812));
    L6MUX21 i15429 (.D0(n33810), .D1(n33811), .SD(y_1_delay[3]), .Z(n33813));
    L6MUX21 i15738 (.D0(n34118), .D1(n34119), .SD(y_1_delay[3]), .Z(n34122));
    L6MUX21 i15739 (.D0(n34120), .D1(n34121), .SD(y_1_delay[3]), .Z(n34123));
    L6MUX21 i15459 (.D0(n33839), .D1(n33840), .SD(y_1_delay[3]), .Z(n33843));
    L6MUX21 i15460 (.D0(n33841), .D1(n33842), .SD(y_1_delay[3]), .Z(n33844));
    L6MUX21 i14932 (.D0(n33312), .D1(n33313), .SD(y_1_delay[3]), .Z(n33316));
    L6MUX21 i15118 (.D0(n33498), .D1(n33499), .SD(y_1_delay[3]), .Z(n33502));
    L6MUX21 i15490 (.D0(n33870), .D1(n33871), .SD(y_1_delay[3]), .Z(n33874));
    L6MUX21 i15491 (.D0(n33872), .D1(n33873), .SD(y_1_delay[3]), .Z(n33875));
    L6MUX21 i14933 (.D0(n33314), .D1(n33315), .SD(y_1_delay[3]), .Z(n33317));
    L6MUX21 i15769 (.D0(n34149), .D1(n34150), .SD(y_1_delay[3]), .Z(n34153));
    L6MUX21 i15119 (.D0(n33500), .D1(n33501), .SD(y_1_delay[3]), .Z(n33503));
    L6MUX21 i15770 (.D0(n34151), .D1(n34152), .SD(y_1_delay[3]), .Z(n34154));
    L6MUX21 i15180 (.D0(n33560), .D1(n33561), .SD(y_1_delay[3]), .Z(n33564));
    L6MUX21 i15181 (.D0(n33562), .D1(n33563), .SD(y_1_delay[3]), .Z(n33565));
    L6MUX21 i15025 (.D0(n33405), .D1(n33406), .SD(y_1_delay[3]), .Z(n33409));
    L6MUX21 i15026 (.D0(n33407), .D1(n33408), .SD(y_1_delay[3]), .Z(n33410));
    LUT4 i15040_3_lut (.A(\result_i[24] [12]), .B(\result_i[25] [12]), .C(y_1_delay[0]), 
         .Z(n33424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15040_3_lut.init = 16'hcaca;
    LUT4 i15443_3_lut (.A(\result_r[24] [14]), .B(\result_r[25] [14]), .C(y_1_delay[0]), 
         .Z(n33827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15443_3_lut.init = 16'hcaca;
    LUT4 i15039_3_lut (.A(\result_i[22] [12]), .B(\result_i[23] [12]), .C(y_1_delay[0]), 
         .Z(n33423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15039_3_lut.init = 16'hcaca;
    L6MUX21 i15521 (.D0(n33901), .D1(n33902), .SD(y_1_delay[3]), .Z(n33905));
    L6MUX21 i15522 (.D0(n33903), .D1(n33904), .SD(y_1_delay[3]), .Z(n33906));
    L6MUX21 i15800 (.D0(n34180), .D1(n34181), .SD(y_1_delay[3]), .Z(n34184));
    L6MUX21 i15801 (.D0(n34182), .D1(n34183), .SD(y_1_delay[3]), .Z(n34185));
    L6MUX21 i15831 (.D0(n34211), .D1(n34212), .SD(y_1_delay[3]), .Z(n34215));
    L6MUX21 i15832 (.D0(n34213), .D1(n34214), .SD(y_1_delay[3]), .Z(n34216));
    L6MUX21 i15552 (.D0(n33932), .D1(n33933), .SD(y_1_delay[3]), .Z(n33936));
    L6MUX21 i15553 (.D0(n33934), .D1(n33935), .SD(y_1_delay[3]), .Z(n33937));
    L6MUX21 i15211 (.D0(n33591), .D1(n33592), .SD(y_1_delay[3]), .Z(n33595));
    L6MUX21 i15212 (.D0(n33593), .D1(n33594), .SD(y_1_delay[3]), .Z(n33596));
    L6MUX21 i15862 (.D0(n34242), .D1(n34243), .SD(y_1_delay[3]), .Z(n34246));
    L6MUX21 i15583 (.D0(n33963), .D1(n33964), .SD(y_1_delay[3]), .Z(n33967));
    L6MUX21 i15584 (.D0(n33965), .D1(n33966), .SD(y_1_delay[3]), .Z(n33968));
    L6MUX21 i15863 (.D0(n34244), .D1(n34245), .SD(y_1_delay[3]), .Z(n34247));
    L6MUX21 i15614 (.D0(n33994), .D1(n33995), .SD(y_1_delay[3]), .Z(n33998));
    L6MUX21 i15615 (.D0(n33996), .D1(n33997), .SD(y_1_delay[3]), .Z(n33999));
    L6MUX21 i15242 (.D0(n33622), .D1(n33623), .SD(y_1_delay[3]), .Z(n33626));
    L6MUX21 i15243 (.D0(n33624), .D1(n33625), .SD(y_1_delay[3]), .Z(n33627));
    L6MUX21 i15056 (.D0(n33436), .D1(n33437), .SD(y_1_delay[3]), .Z(n33440));
    L6MUX21 i15645 (.D0(n34025), .D1(n34026), .SD(y_1_delay[3]), .Z(n34029));
    L6MUX21 i15646 (.D0(n34027), .D1(n34028), .SD(y_1_delay[3]), .Z(n34030));
    L6MUX21 i15057 (.D0(n33438), .D1(n33439), .SD(y_1_delay[3]), .Z(n33441));
    L6MUX21 i15273 (.D0(n33653), .D1(n33654), .SD(y_1_delay[3]), .Z(n33657));
    L6MUX21 i15274 (.D0(n33655), .D1(n33656), .SD(y_1_delay[3]), .Z(n33658));
    L6MUX21 i15676 (.D0(n34056), .D1(n34057), .SD(y_1_delay[3]), .Z(n34060));
    L6MUX21 i15677 (.D0(n34058), .D1(n34059), .SD(y_1_delay[3]), .Z(n34061));
    LUT4 i15442_3_lut (.A(\result_r[22] [14]), .B(\result_r[23] [14]), .C(y_1_delay[0]), 
         .Z(n33826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15442_3_lut.init = 16'hcaca;
    LUT4 i15038_3_lut (.A(\result_i[20] [12]), .B(\result_i[21] [12]), .C(y_1_delay[0]), 
         .Z(n33422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15038_3_lut.init = 16'hcaca;
    L6MUX21 i15149 (.D0(n33529), .D1(n33530), .SD(y_1_delay[3]), .Z(n33533));
    LUT4 i15441_3_lut (.A(\result_r[20] [14]), .B(\result_r[21] [14]), .C(y_1_delay[0]), 
         .Z(n33825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15441_3_lut.init = 16'hcaca;
    L6MUX21 i15150 (.D0(n33531), .D1(n33532), .SD(y_1_delay[3]), .Z(n33534));
    L6MUX21 i15304 (.D0(n33684), .D1(n33685), .SD(y_1_delay[3]), .Z(n33688));
    L6MUX21 i15305 (.D0(n33686), .D1(n33687), .SD(y_1_delay[3]), .Z(n33689));
    L6MUX21 i14961 (.D0(n33339), .D1(n33340), .SD(y_1_delay[2]), .Z(n33345));
    L6MUX21 i14962 (.D0(n33341), .D1(n33342), .SD(y_1_delay[2]), .Z(n33346));
    L6MUX21 i15083 (.D0(n33459), .D1(n33460), .SD(y_1_delay[2]), .Z(n33467));
    L6MUX21 i15084 (.D0(n33461), .D1(n33462), .SD(y_1_delay[2]), .Z(n33468));
    L6MUX21 i15085 (.D0(n33463), .D1(n33464), .SD(y_1_delay[2]), .Z(n33469));
    L6MUX21 i15331 (.D0(n33707), .D1(n33708), .SD(y_1_delay[2]), .Z(n33715));
    L6MUX21 i15332 (.D0(n33709), .D1(n33710), .SD(y_1_delay[2]), .Z(n33716));
    L6MUX21 i15333 (.D0(n33711), .D1(n33712), .SD(y_1_delay[2]), .Z(n33717));
    L6MUX21 i15334 (.D0(n33713), .D1(n33714), .SD(y_1_delay[2]), .Z(n33718));
    L6MUX21 i15086 (.D0(n33465), .D1(n33466), .SD(y_1_delay[2]), .Z(n33470));
    L6MUX21 i15362 (.D0(n33738), .D1(n33739), .SD(y_1_delay[2]), .Z(n33746));
    L6MUX21 i15363 (.D0(n33740), .D1(n33741), .SD(y_1_delay[2]), .Z(n33747));
    L6MUX21 i15364 (.D0(n33742), .D1(n33743), .SD(y_1_delay[2]), .Z(n33748));
    L6MUX21 i15365 (.D0(n33744), .D1(n33745), .SD(y_1_delay[2]), .Z(n33749));
    L6MUX21 i15703 (.D0(n34079), .D1(n34080), .SD(y_1_delay[2]), .Z(n34087));
    L6MUX21 i15704 (.D0(n34081), .D1(n34082), .SD(y_1_delay[2]), .Z(n34088));
    L6MUX21 i15705 (.D0(n34083), .D1(n34084), .SD(y_1_delay[2]), .Z(n34089));
    L6MUX21 i15706 (.D0(n34085), .D1(n34086), .SD(y_1_delay[2]), .Z(n34090));
    LUT4 i15037_3_lut (.A(\result_i[18] [12]), .B(\result_i[19] [12]), .C(y_1_delay[0]), 
         .Z(n33421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15037_3_lut.init = 16'hcaca;
    L6MUX21 i14897 (.D0(n33273), .D1(n33274), .SD(y_1_delay[2]), .Z(n33281));
    L6MUX21 i14898 (.D0(n33275), .D1(n33276), .SD(y_1_delay[2]), .Z(n33282));
    L6MUX21 i14899 (.D0(n33277), .D1(n33278), .SD(y_1_delay[2]), .Z(n33283));
    L6MUX21 i14900 (.D0(n33279), .D1(n33280), .SD(y_1_delay[2]), .Z(n33284));
    L6MUX21 i15393 (.D0(n33769), .D1(n33770), .SD(y_1_delay[2]), .Z(n33777));
    L6MUX21 i14990 (.D0(n33366), .D1(n33367), .SD(y_1_delay[2]), .Z(n33374));
    L6MUX21 i14991 (.D0(n33368), .D1(n33369), .SD(y_1_delay[2]), .Z(n33375));
    L6MUX21 i14992 (.D0(n33370), .D1(n33371), .SD(y_1_delay[2]), .Z(n33376));
    L6MUX21 i14993 (.D0(n33372), .D1(n33373), .SD(y_1_delay[2]), .Z(n33377));
    L6MUX21 i15394 (.D0(n33771), .D1(n33772), .SD(y_1_delay[2]), .Z(n33778));
    L6MUX21 i15395 (.D0(n33773), .D1(n33774), .SD(y_1_delay[2]), .Z(n33779));
    L6MUX21 i15396 (.D0(n33775), .D1(n33776), .SD(y_1_delay[2]), .Z(n33780));
    L6MUX21 i14928 (.D0(n33304), .D1(n33305), .SD(y_1_delay[2]), .Z(n33312));
    L6MUX21 i14929 (.D0(n33306), .D1(n33307), .SD(y_1_delay[2]), .Z(n33313));
    L6MUX21 i14930 (.D0(n33308), .D1(n33309), .SD(y_1_delay[2]), .Z(n33314));
    L6MUX21 i14959 (.D0(n33335), .D1(n33336), .SD(y_1_delay[2]), .Z(n33343));
    L6MUX21 i14960 (.D0(n33337), .D1(n33338), .SD(y_1_delay[2]), .Z(n33344));
    L6MUX21 i15424 (.D0(n33800), .D1(n33801), .SD(y_1_delay[2]), .Z(n33808));
    L6MUX21 i15425 (.D0(n33802), .D1(n33803), .SD(y_1_delay[2]), .Z(n33809));
    L6MUX21 i15426 (.D0(n33804), .D1(n33805), .SD(y_1_delay[2]), .Z(n33810));
    L6MUX21 i15427 (.D0(n33806), .D1(n33807), .SD(y_1_delay[2]), .Z(n33811));
    L6MUX21 i15021 (.D0(n33397), .D1(n33398), .SD(y_1_delay[2]), .Z(n33405));
    L6MUX21 i15734 (.D0(n34110), .D1(n34111), .SD(y_1_delay[2]), .Z(n34118));
    L6MUX21 i15735 (.D0(n34112), .D1(n34113), .SD(y_1_delay[2]), .Z(n34119));
    L6MUX21 i15736 (.D0(n34114), .D1(n34115), .SD(y_1_delay[2]), .Z(n34120));
    L6MUX21 i15737 (.D0(n34116), .D1(n34117), .SD(y_1_delay[2]), .Z(n34121));
    L6MUX21 i14931 (.D0(n33310), .D1(n33311), .SD(y_1_delay[2]), .Z(n33315));
    L6MUX21 i15022 (.D0(n33399), .D1(n33400), .SD(y_1_delay[2]), .Z(n33406));
    L6MUX21 i15455 (.D0(n33831), .D1(n33832), .SD(y_1_delay[2]), .Z(n33839));
    L6MUX21 i15456 (.D0(n33833), .D1(n33834), .SD(y_1_delay[2]), .Z(n33840));
    L6MUX21 i15457 (.D0(n33835), .D1(n33836), .SD(y_1_delay[2]), .Z(n33841));
    L6MUX21 i15458 (.D0(n33837), .D1(n33838), .SD(y_1_delay[2]), .Z(n33842));
    L6MUX21 i15114 (.D0(n33490), .D1(n33491), .SD(y_1_delay[2]), .Z(n33498));
    L6MUX21 i15023 (.D0(n33401), .D1(n33402), .SD(y_1_delay[2]), .Z(n33407));
    L6MUX21 i15115 (.D0(n33492), .D1(n33493), .SD(y_1_delay[2]), .Z(n33499));
    L6MUX21 i15116 (.D0(n33494), .D1(n33495), .SD(y_1_delay[2]), .Z(n33500));
    L6MUX21 i15117 (.D0(n33496), .D1(n33497), .SD(y_1_delay[2]), .Z(n33501));
    L6MUX21 i15486 (.D0(n33862), .D1(n33863), .SD(y_1_delay[2]), .Z(n33870));
    L6MUX21 i15487 (.D0(n33864), .D1(n33865), .SD(y_1_delay[2]), .Z(n33871));
    L6MUX21 i15488 (.D0(n33866), .D1(n33867), .SD(y_1_delay[2]), .Z(n33872));
    L6MUX21 i15489 (.D0(n33868), .D1(n33869), .SD(y_1_delay[2]), .Z(n33873));
    L6MUX21 i15176 (.D0(n33552), .D1(n33553), .SD(y_1_delay[2]), .Z(n33560));
    L6MUX21 i15765 (.D0(n34141), .D1(n34142), .SD(y_1_delay[2]), .Z(n34149));
    L6MUX21 i15766 (.D0(n34143), .D1(n34144), .SD(y_1_delay[2]), .Z(n34150));
    L6MUX21 i15767 (.D0(n34145), .D1(n34146), .SD(y_1_delay[2]), .Z(n34151));
    L6MUX21 i15177 (.D0(n33554), .D1(n33555), .SD(y_1_delay[2]), .Z(n33561));
    L6MUX21 i15768 (.D0(n34147), .D1(n34148), .SD(y_1_delay[2]), .Z(n34152));
    L6MUX21 i15024 (.D0(n33403), .D1(n33404), .SD(y_1_delay[2]), .Z(n33408));
    L6MUX21 i15178 (.D0(n33556), .D1(n33557), .SD(y_1_delay[2]), .Z(n33562));
    L6MUX21 i15179 (.D0(n33558), .D1(n33559), .SD(y_1_delay[2]), .Z(n33563));
    L6MUX21 i15517 (.D0(n33893), .D1(n33894), .SD(y_1_delay[2]), .Z(n33901));
    L6MUX21 i15518 (.D0(n33895), .D1(n33896), .SD(y_1_delay[2]), .Z(n33902));
    L6MUX21 i15519 (.D0(n33897), .D1(n33898), .SD(y_1_delay[2]), .Z(n33903));
    L6MUX21 i15520 (.D0(n33899), .D1(n33900), .SD(y_1_delay[2]), .Z(n33904));
    L6MUX21 i15796 (.D0(n34172), .D1(n34173), .SD(y_1_delay[2]), .Z(n34180));
    L6MUX21 i15797 (.D0(n34174), .D1(n34175), .SD(y_1_delay[2]), .Z(n34181));
    L6MUX21 i15798 (.D0(n34176), .D1(n34177), .SD(y_1_delay[2]), .Z(n34182));
    L6MUX21 i15799 (.D0(n34178), .D1(n34179), .SD(y_1_delay[2]), .Z(n34183));
    L6MUX21 i15827 (.D0(n34203), .D1(n34204), .SD(y_1_delay[2]), .Z(n34211));
    L6MUX21 i15828 (.D0(n34205), .D1(n34206), .SD(y_1_delay[2]), .Z(n34212));
    L6MUX21 i15829 (.D0(n34207), .D1(n34208), .SD(y_1_delay[2]), .Z(n34213));
    L6MUX21 i15830 (.D0(n34209), .D1(n34210), .SD(y_1_delay[2]), .Z(n34214));
    L6MUX21 i15548 (.D0(n33924), .D1(n33925), .SD(y_1_delay[2]), .Z(n33932));
    L6MUX21 i15549 (.D0(n33926), .D1(n33927), .SD(y_1_delay[2]), .Z(n33933));
    L6MUX21 i15550 (.D0(n33928), .D1(n33929), .SD(y_1_delay[2]), .Z(n33934));
    L6MUX21 i15551 (.D0(n33930), .D1(n33931), .SD(y_1_delay[2]), .Z(n33935));
    L6MUX21 i15207 (.D0(n33583), .D1(n33584), .SD(y_1_delay[2]), .Z(n33591));
    L6MUX21 i15208 (.D0(n33585), .D1(n33586), .SD(y_1_delay[2]), .Z(n33592));
    L6MUX21 i15209 (.D0(n33587), .D1(n33588), .SD(y_1_delay[2]), .Z(n33593));
    L6MUX21 i15210 (.D0(n33589), .D1(n33590), .SD(y_1_delay[2]), .Z(n33594));
    L6MUX21 i15858 (.D0(n34234), .D1(n34235), .SD(y_1_delay[2]), .Z(n34242));
    L6MUX21 i15859 (.D0(n34236), .D1(n34237), .SD(y_1_delay[2]), .Z(n34243));
    L6MUX21 i15860 (.D0(n34238), .D1(n34239), .SD(y_1_delay[2]), .Z(n34244));
    L6MUX21 i15579 (.D0(n33955), .D1(n33956), .SD(y_1_delay[2]), .Z(n33963));
    L6MUX21 i15580 (.D0(n33957), .D1(n33958), .SD(y_1_delay[2]), .Z(n33964));
    L6MUX21 i15861 (.D0(n34240), .D1(n34241), .SD(y_1_delay[2]), .Z(n34245));
    L6MUX21 i15581 (.D0(n33959), .D1(n33960), .SD(y_1_delay[2]), .Z(n33965));
    L6MUX21 i15582 (.D0(n33961), .D1(n33962), .SD(y_1_delay[2]), .Z(n33966));
    L6MUX21 i15610 (.D0(n33986), .D1(n33987), .SD(y_1_delay[2]), .Z(n33994));
    L6MUX21 i15611 (.D0(n33988), .D1(n33989), .SD(y_1_delay[2]), .Z(n33995));
    L6MUX21 i15238 (.D0(n33614), .D1(n33615), .SD(y_1_delay[2]), .Z(n33622));
    L6MUX21 i15612 (.D0(n33990), .D1(n33991), .SD(y_1_delay[2]), .Z(n33996));
    L6MUX21 i15613 (.D0(n33992), .D1(n33993), .SD(y_1_delay[2]), .Z(n33997));
    L6MUX21 i15239 (.D0(n33616), .D1(n33617), .SD(y_1_delay[2]), .Z(n33623));
    L6MUX21 i15240 (.D0(n33618), .D1(n33619), .SD(y_1_delay[2]), .Z(n33624));
    L6MUX21 i15241 (.D0(n33620), .D1(n33621), .SD(y_1_delay[2]), .Z(n33625));
    L6MUX21 i15052 (.D0(n33428), .D1(n33429), .SD(y_1_delay[2]), .Z(n33436));
    L6MUX21 i15053 (.D0(n33430), .D1(n33431), .SD(y_1_delay[2]), .Z(n33437));
    L6MUX21 i15054 (.D0(n33432), .D1(n33433), .SD(y_1_delay[2]), .Z(n33438));
    L6MUX21 i15055 (.D0(n33434), .D1(n33435), .SD(y_1_delay[2]), .Z(n33439));
    L6MUX21 i15641 (.D0(n34017), .D1(n34018), .SD(y_1_delay[2]), .Z(n34025));
    L6MUX21 i15642 (.D0(n34019), .D1(n34020), .SD(y_1_delay[2]), .Z(n34026));
    L6MUX21 i15643 (.D0(n34021), .D1(n34022), .SD(y_1_delay[2]), .Z(n34027));
    L6MUX21 i15644 (.D0(n34023), .D1(n34024), .SD(y_1_delay[2]), .Z(n34028));
    L6MUX21 i15269 (.D0(n33645), .D1(n33646), .SD(y_1_delay[2]), .Z(n33653));
    L6MUX21 i15270 (.D0(n33647), .D1(n33648), .SD(y_1_delay[2]), .Z(n33654));
    L6MUX21 i15271 (.D0(n33649), .D1(n33650), .SD(y_1_delay[2]), .Z(n33655));
    L6MUX21 i15272 (.D0(n33651), .D1(n33652), .SD(y_1_delay[2]), .Z(n33656));
    L6MUX21 i15145 (.D0(n33521), .D1(n33522), .SD(y_1_delay[2]), .Z(n33529));
    L6MUX21 i15146 (.D0(n33523), .D1(n33524), .SD(y_1_delay[2]), .Z(n33530));
    L6MUX21 i15147 (.D0(n33525), .D1(n33526), .SD(y_1_delay[2]), .Z(n33531));
    L6MUX21 i15672 (.D0(n34048), .D1(n34049), .SD(y_1_delay[2]), .Z(n34056));
    L6MUX21 i15673 (.D0(n34050), .D1(n34051), .SD(y_1_delay[2]), .Z(n34057));
    L6MUX21 i15674 (.D0(n34052), .D1(n34053), .SD(y_1_delay[2]), .Z(n34058));
    L6MUX21 i15675 (.D0(n34054), .D1(n34055), .SD(y_1_delay[2]), .Z(n34059));
    L6MUX21 i15148 (.D0(n33527), .D1(n33528), .SD(y_1_delay[2]), .Z(n33532));
    L6MUX21 i15300 (.D0(n33676), .D1(n33677), .SD(y_1_delay[2]), .Z(n33684));
    L6MUX21 i15301 (.D0(n33678), .D1(n33679), .SD(y_1_delay[2]), .Z(n33685));
    L6MUX21 i15302 (.D0(n33680), .D1(n33681), .SD(y_1_delay[2]), .Z(n33686));
    L6MUX21 i15303 (.D0(n33682), .D1(n33683), .SD(y_1_delay[2]), .Z(n33687));
    PFUMX i15075 (.BLUT(n33443), .ALUT(n33444), .C0(y_1_delay[1]), .Z(n33459));
    PFUMX i15076 (.BLUT(n33445), .ALUT(n33446), .C0(y_1_delay[1]), .Z(n33460));
    PFUMX i14951 (.BLUT(n33319), .ALUT(n33320), .C0(y_1_delay[1]), .Z(n33335));
    PFUMX i15695 (.BLUT(n34063), .ALUT(n34064), .C0(y_1_delay[1]), .Z(n34079));
    PFUMX i15696 (.BLUT(n34065), .ALUT(n34066), .C0(y_1_delay[1]), .Z(n34080));
    PFUMX i15077 (.BLUT(n33447), .ALUT(n33448), .C0(y_1_delay[1]), .Z(n33461));
    PFUMX i15078 (.BLUT(n33449), .ALUT(n33450), .C0(y_1_delay[1]), .Z(n33462));
    PFUMX i15323 (.BLUT(n33691), .ALUT(n33692), .C0(y_1_delay[1]), .Z(n33707));
    PFUMX i15697 (.BLUT(n34067), .ALUT(n34068), .C0(y_1_delay[1]), .Z(n34081));
    PFUMX i15079 (.BLUT(n33451), .ALUT(n33452), .C0(y_1_delay[1]), .Z(n33463));
    PFUMX i15698 (.BLUT(n34069), .ALUT(n34070), .C0(y_1_delay[1]), .Z(n34082));
    PFUMX i15080 (.BLUT(n33453), .ALUT(n33454), .C0(y_1_delay[1]), .Z(n33464));
    PFUMX i15324 (.BLUT(n33693), .ALUT(n33694), .C0(y_1_delay[1]), .Z(n33708));
    PFUMX i15081 (.BLUT(n33455), .ALUT(n33456), .C0(y_1_delay[1]), .Z(n33465));
    PFUMX i15325 (.BLUT(n33695), .ALUT(n33696), .C0(y_1_delay[1]), .Z(n33709));
    PFUMX i15082 (.BLUT(n33457), .ALUT(n33458), .C0(y_1_delay[1]), .Z(n33466));
    PFUMX i15699 (.BLUT(n34071), .ALUT(n34072), .C0(y_1_delay[1]), .Z(n34083));
    PFUMX i15326 (.BLUT(n33697), .ALUT(n33698), .C0(y_1_delay[1]), .Z(n33710));
    PFUMX i15327 (.BLUT(n33699), .ALUT(n33700), .C0(y_1_delay[1]), .Z(n33711));
    PFUMX i15328 (.BLUT(n33701), .ALUT(n33702), .C0(y_1_delay[1]), .Z(n33712));
    PFUMX i15329 (.BLUT(n33703), .ALUT(n33704), .C0(y_1_delay[1]), .Z(n33713));
    PFUMX i15330 (.BLUT(n33705), .ALUT(n33706), .C0(y_1_delay[1]), .Z(n33714));
    PFUMX i15354 (.BLUT(n33722), .ALUT(n33723), .C0(y_1_delay[1]), .Z(n33738));
    PFUMX i15355 (.BLUT(n33724), .ALUT(n33725), .C0(y_1_delay[1]), .Z(n33739));
    PFUMX i15356 (.BLUT(n33726), .ALUT(n33727), .C0(y_1_delay[1]), .Z(n33740));
    PFUMX i15357 (.BLUT(n33728), .ALUT(n33729), .C0(y_1_delay[1]), .Z(n33741));
    PFUMX i15358 (.BLUT(n33730), .ALUT(n33731), .C0(y_1_delay[1]), .Z(n33742));
    PFUMX i15359 (.BLUT(n33732), .ALUT(n33733), .C0(y_1_delay[1]), .Z(n33743));
    PFUMX i15360 (.BLUT(n33734), .ALUT(n33735), .C0(y_1_delay[1]), .Z(n33744));
    PFUMX i15361 (.BLUT(n33736), .ALUT(n33737), .C0(y_1_delay[1]), .Z(n33745));
    PFUMX i15700 (.BLUT(n34073), .ALUT(n34074), .C0(y_1_delay[1]), .Z(n34084));
    PFUMX i15701 (.BLUT(n34075), .ALUT(n34076), .C0(y_1_delay[1]), .Z(n34085));
    PFUMX i15702 (.BLUT(n34077), .ALUT(n34078), .C0(y_1_delay[1]), .Z(n34086));
    PFUMX i14889 (.BLUT(n33257), .ALUT(n33258), .C0(y_1_delay[1]), .Z(n33273));
    PFUMX i14890 (.BLUT(n33259), .ALUT(n33260), .C0(y_1_delay[1]), .Z(n33274));
    PFUMX i14891 (.BLUT(n33261), .ALUT(n33262), .C0(y_1_delay[1]), .Z(n33275));
    PFUMX i14892 (.BLUT(n33263), .ALUT(n33264), .C0(y_1_delay[1]), .Z(n33276));
    PFUMX i14893 (.BLUT(n33265), .ALUT(n33266), .C0(y_1_delay[1]), .Z(n33277));
    PFUMX i14894 (.BLUT(n33267), .ALUT(n33268), .C0(y_1_delay[1]), .Z(n33278));
    PFUMX i14895 (.BLUT(n33269), .ALUT(n33270), .C0(y_1_delay[1]), .Z(n33279));
    PFUMX i14896 (.BLUT(n33271), .ALUT(n33272), .C0(y_1_delay[1]), .Z(n33280));
    PFUMX i15385 (.BLUT(n33753), .ALUT(n33754), .C0(y_1_delay[1]), .Z(n33769));
    PFUMX i15386 (.BLUT(n33755), .ALUT(n33756), .C0(y_1_delay[1]), .Z(n33770));
    PFUMX i15387 (.BLUT(n33757), .ALUT(n33758), .C0(y_1_delay[1]), .Z(n33771));
    PFUMX i15388 (.BLUT(n33759), .ALUT(n33760), .C0(y_1_delay[1]), .Z(n33772));
    PFUMX i15389 (.BLUT(n33761), .ALUT(n33762), .C0(y_1_delay[1]), .Z(n33773));
    PFUMX i15390 (.BLUT(n33763), .ALUT(n33764), .C0(y_1_delay[1]), .Z(n33774));
    PFUMX i15391 (.BLUT(n33765), .ALUT(n33766), .C0(y_1_delay[1]), .Z(n33775));
    PFUMX i15392 (.BLUT(n33767), .ALUT(n33768), .C0(y_1_delay[1]), .Z(n33776));
    PFUMX i14952 (.BLUT(n33321), .ALUT(n33322), .C0(y_1_delay[1]), .Z(n33336));
    PFUMX i14982 (.BLUT(n33350), .ALUT(n33351), .C0(y_1_delay[1]), .Z(n33366));
    PFUMX i14983 (.BLUT(n33352), .ALUT(n33353), .C0(y_1_delay[1]), .Z(n33367));
    PFUMX i14984 (.BLUT(n33354), .ALUT(n33355), .C0(y_1_delay[1]), .Z(n33368));
    PFUMX i14985 (.BLUT(n33356), .ALUT(n33357), .C0(y_1_delay[1]), .Z(n33369));
    PFUMX i14920 (.BLUT(n33288), .ALUT(n33289), .C0(y_1_delay[1]), .Z(n33304));
    PFUMX i14986 (.BLUT(n33358), .ALUT(n33359), .C0(y_1_delay[1]), .Z(n33370));
    PFUMX i14921 (.BLUT(n33290), .ALUT(n33291), .C0(y_1_delay[1]), .Z(n33305));
    PFUMX i14922 (.BLUT(n33292), .ALUT(n33293), .C0(y_1_delay[1]), .Z(n33306));
    PFUMX i14923 (.BLUT(n33294), .ALUT(n33295), .C0(y_1_delay[1]), .Z(n33307));
    PFUMX i14987 (.BLUT(n33360), .ALUT(n33361), .C0(y_1_delay[1]), .Z(n33371));
    PFUMX i14924 (.BLUT(n33296), .ALUT(n33297), .C0(y_1_delay[1]), .Z(n33308));
    PFUMX i14988 (.BLUT(n33362), .ALUT(n33363), .C0(y_1_delay[1]), .Z(n33372));
    PFUMX i14989 (.BLUT(n33364), .ALUT(n33365), .C0(y_1_delay[1]), .Z(n33373));
    PFUMX i14925 (.BLUT(n33298), .ALUT(n33299), .C0(y_1_delay[1]), .Z(n33309));
    PFUMX i14926 (.BLUT(n33300), .ALUT(n33301), .C0(y_1_delay[1]), .Z(n33310));
    PFUMX i15726 (.BLUT(n34094), .ALUT(n34095), .C0(y_1_delay[1]), .Z(n34110));
    PFUMX i14927 (.BLUT(n33302), .ALUT(n33303), .C0(y_1_delay[1]), .Z(n33311));
    PFUMX i15727 (.BLUT(n34096), .ALUT(n34097), .C0(y_1_delay[1]), .Z(n34111));
    PFUMX i15728 (.BLUT(n34098), .ALUT(n34099), .C0(y_1_delay[1]), .Z(n34112));
    PFUMX i14953 (.BLUT(n33323), .ALUT(n33324), .C0(y_1_delay[1]), .Z(n33337));
    PFUMX i15729 (.BLUT(n34100), .ALUT(n34101), .C0(y_1_delay[1]), .Z(n34113));
    LUT4 i15440_3_lut (.A(\result_r[18] [14]), .B(\result_r[19] [14]), .C(y_1_delay[0]), 
         .Z(n33824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15440_3_lut.init = 16'hcaca;
    LUT4 i2606_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[496])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2606_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2598_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[497])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2598_3_lut_4_lut.init = 16'hf1e0;
    radix2_U1 radix_no3 (.shift_4_dout_i({shift_4_dout_i}), .n12300(n12300), 
            .n12301(n12301), .n12302(n12302), .n12303(n12303), .n12304(n12304), 
            .n12305(n12305), .n12306(n12306), .n12307(n12307), .n12308(n12308), 
            .n12309(n12309), .n119(n119_adj_6625), .GND_net(GND_net), 
            .VCC_net(VCC_net), .\op_r_23__N_1268[0] (op_r_23__N_1268_adj_7375[0]), 
            .\op_r_23__N_1268[1] (op_r_23__N_1268_adj_7375[1]), .\op_r_23__N_1268[2] (op_r_23__N_1268_adj_7375[2]), 
            .\op_r_23__N_1268[3] (op_r_23__N_1268_adj_7375[3]), .\op_r_23__N_1268[4] (op_r_23__N_1268_adj_7375[4]), 
            .\op_r_23__N_1268[5] (op_r_23__N_1268_adj_7375[5]), .\op_r_23__N_1268[6] (op_r_23__N_1268_adj_7375[6]), 
            .\op_r_23__N_1268[7] (op_r_23__N_1268_adj_7375[7]), .\op_r_23__N_1268[8] (op_r_23__N_1268_adj_7375[8]), 
            .\op_r_23__N_1268[9] (op_r_23__N_1268_adj_7375[9]), .\op_r_23__N_1268[10] (op_r_23__N_1268_adj_7375[10]), 
            .\op_r_23__N_1268[11] (op_r_23__N_1268_adj_7375[11]), .\op_r_23__N_1268[12] (op_r_23__N_1268_adj_7375[12]), 
            .\op_r_23__N_1268[13] (op_r_23__N_1268_adj_7375[13]), .\op_r_23__N_1268[14] (op_r_23__N_1268_adj_7375[14]), 
            .\op_r_23__N_1268[15] (op_r_23__N_1268_adj_7375[15]), .\op_r_23__N_1268[16] (op_r_23__N_1268_adj_7375[16]), 
            .\op_r_23__N_1268[17] (op_r_23__N_1268_adj_7375[17]), .\op_r_23__N_1226[0] (op_r_23__N_1226_adj_7377[0]), 
            .\op_r_23__N_1226[1] (op_r_23__N_1226_adj_7377[1]), .\op_r_23__N_1226[2] (op_r_23__N_1226_adj_7377[2]), 
            .\op_r_23__N_1226[3] (op_r_23__N_1226_adj_7377[3]), .\op_r_23__N_1226[4] (op_r_23__N_1226_adj_7377[4]), 
            .\op_r_23__N_1226[5] (op_r_23__N_1226_adj_7377[5]), .\op_r_23__N_1226[6] (op_r_23__N_1226_adj_7377[6]), 
            .\op_r_23__N_1226[7] (op_r_23__N_1226_adj_7377[7]), .\op_r_23__N_1226[8] (op_r_23__N_1226_adj_7377[8]), 
            .\op_r_23__N_1226[9] (op_r_23__N_1226_adj_7377[9]), .\op_r_23__N_1226[10] (op_r_23__N_1226_adj_7377[10]), 
            .\op_r_23__N_1226[11] (op_r_23__N_1226_adj_7377[11]), .\op_r_23__N_1226[12] (op_r_23__N_1226_adj_7377[12]), 
            .\op_r_23__N_1226[13] (op_r_23__N_1226_adj_7377[13]), .\op_r_23__N_1226[14] (op_r_23__N_1226_adj_7377[14]), 
            .\op_r_23__N_1226[15] (op_r_23__N_1226_adj_7377[15]), .\op_r_23__N_1226[16] (op_r_23__N_1226_adj_7377[16]), 
            .\op_r_23__N_1226[17] (op_r_23__N_1226_adj_7377[17]), .\op_r_23__N_1226[18] (op_r_23__N_1226_adj_7377[18]), 
            .\op_r_23__N_1226[19] (op_r_23__N_1226_adj_7377[19]), .\op_r_23__N_1226[20] (op_r_23__N_1226_adj_7377[20]), 
            .\op_r_23__N_1226[21] (op_r_23__N_1226_adj_7377[21]), .\op_r_23__N_1226[22] (op_r_23__N_1226_adj_7377[22]), 
            .\op_r_23__N_1226[23] (op_r_23__N_1226_adj_7377[23]), .\op_r_23__N_1226[24] (op_r_23__N_1226_adj_7377[24]), 
            .\op_r_23__N_1226[25] (op_r_23__N_1226_adj_7377[25]), .\op_r_23__N_1226[26] (op_r_23__N_1226_adj_7377[26]), 
            .\op_r_23__N_1226[27] (op_r_23__N_1226_adj_7377[27]), .\op_r_23__N_1226[28] (op_r_23__N_1226_adj_7377[28]), 
            .\op_r_23__N_1226[29] (op_r_23__N_1226_adj_7377[29]), .\op_r_23__N_1226[30] (op_r_23__N_1226_adj_7377[30]), 
            .\op_r_23__N_1226[31] (op_r_23__N_1226_adj_7377[31]), .\op_r_23__N_1268[18] (op_r_23__N_1268_adj_7375[18]), 
            .\op_r_23__N_1268[19] (op_r_23__N_1268_adj_7375[19]), .\op_r_23__N_1268[20] (op_r_23__N_1268_adj_7375[20]), 
            .\op_r_23__N_1268[21] (op_r_23__N_1268_adj_7375[21]), .\op_r_23__N_1268[22] (op_r_23__N_1268_adj_7375[22]), 
            .\op_r_23__N_1268[23] (op_r_23__N_1268_adj_7375[23]), .\op_r_23__N_1268[24] (op_r_23__N_1268_adj_7375[24]), 
            .\op_r_23__N_1268[25] (op_r_23__N_1268_adj_7375[25]), .\op_r_23__N_1268[26] (op_r_23__N_1268_adj_7375[26]), 
            .\op_r_23__N_1268[27] (op_r_23__N_1268_adj_7375[27]), .\op_r_23__N_1268[28] (op_r_23__N_1268_adj_7375[28]), 
            .\op_r_23__N_1268[29] (op_r_23__N_1268_adj_7375[29]), .\op_r_23__N_1268[30] (op_r_23__N_1268_adj_7375[30]), 
            .\op_r_23__N_1268[31] (op_r_23__N_1268_adj_7375[31]), .n8849(n8849), 
            .n8848(n8848), .n8847(n8847), .n8846(n8846), .n8845(n8845), 
            .n8844(n8844), .n8843(n8843), .n8842(n8842), .n8841(n8841), 
            .n8840(n8840), .n8839(n8839), .n8838(n8838), .n8837(n8837), 
            .n8836(n8836), .n8835(n8835), .n8834(n8834), .n8833(n8833), 
            .n8832(n8832), .n8831(n8831), .n8830(n8830), .n8829(n8829), 
            .n8828(n8828), .n8827(n8827), .n8826(n8826), .n8825(n8825), 
            .n8824(n8824), .n34777(n34777), .\rom4_w_r[1] (rom4_w_r[1]), 
            .\rom4_w_r[5] (rom4_w_r[5]), .\rom4_w_r[8] (rom4_w_r[8]), .n12240(n12240), 
            .n12241(n12241), .n12242(n12242), .n12243(n12243), .n12244(n12244), 
            .n12245(n12245), .n12246(n12246), .n12247(n12247), .n12248(n12248), 
            .n12249(n12249), .n12250(n12250), .n12251(n12251), .n12252(n12252), 
            .n12253(n12253), .n12254(n12254), .n12255(n12255), .n12256(n12256), 
            .n12257(n12257), .\rom4_w_i[12] (rom4_w_i[12]), .n319(n319_adj_6714), 
            .n10718(n10718), .n10719(n10719), .n10720(n10720), .n10721(n10721), 
            .n10722(n10722), .n10723(n10723), .n10724(n10724), .n10725(n10725), 
            .n10726(n10726), .n10727(n10727), .n10728(n10728), .n10729(n10729), 
            .n10730(n10730), .n10731(n10731), .n10732(n10732), .n10733(n10733), 
            .n10734(n10734), .n10735(n10735), .n12258(n12258), .n12259(n12259), 
            .n12260(n12260), .n12261(n12261), .n12262(n12262), .n12263(n12263), 
            .n12264(n12264), .op_i_23__N_1154({op_i_23__N_1154_adj_7371}), 
            .n34841(n34841), .n30179(n30179), .\delay_i_23__N_1202[18] (delay_i_23__N_1202_adj_7428[18]), 
            .\dout_i_23__N_5777[18] (dout_i_23__N_5777[18]), .\delay_i_23__N_1202[2] (delay_i_23__N_1202_adj_7428[2]), 
            .\dout_i_23__N_5777[2] (dout_i_23__N_5777[2]), .\delay_i_23__N_1202[1] (delay_i_23__N_1202_adj_7428[1]), 
            .\dout_i_23__N_5777[1] (dout_i_23__N_5777[1]), .\delay_i_23__N_1202[0] (delay_i_23__N_1202_adj_7428[0]), 
            .\dout_i_23__N_5777[0] (dout_i_23__N_5777[0]), .\rom4_state[0] (rom4_state[0]), 
            .n34799(n34799), .op_r_23__N_1106({op_r_23__N_1106_adj_7370}), 
            .n34610(n34610), .n34609(n34609), .n34576(n34576), .n34575(n34575), 
            .n34690(n34690), .n34612(n34612), .valid(valid_adj_7001), 
            .clk_c_enable_1396(clk_c_enable_1396), .n34621(n34621), .n34665(n34665), 
            .n34593(n34593), .n34578(n34578), .\delay_r_23__N_1178[0] (delay_r_23__N_1178_adj_7427[0]), 
            .\dout_r_23__N_5681[0] (dout_r_23__N_5681[0]), .n34624(n34624), 
            .n34579(n34579), .n34587(n34587), .n34588(n34588), .n34666(n34666), 
            .n34594(n34594), .n34622(n34622), .n34577(n34577), .n34623(n34623), 
            .n34611(n34611), .n34689(n34689), .n34633(n34633), .n34580(n34580), 
            .n34634(n34634), .n34581(n34581), .n34635(n34635), .n34582(n34582), 
            .n34636(n34636), .n34583(n34583), .n34645(n34645), .n34584(n34584), 
            .n34646(n34646), .n34585(n34585), .n34655(n34655), .n34586(n34586), 
            .n34656(n34656), .n34667(n34667), .n34595(n34595), .n34668(n34668), 
            .n34596(n34596), .n34673(n34673), .n34601(n34601), .n34674(n34674), 
            .n34602(n34602), .n34679(n34679), .n34603(n34603), .n34604(n34604), 
            .n34680(n34680)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(149[8] 162[2])
    LUT4 i2590_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[498])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2590_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2582_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[499])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2582_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2574_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[500])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2574_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2566_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[501])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2566_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2558_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[502])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2558_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15439_3_lut (.A(\result_r[16] [14]), .B(\result_r[17] [14]), .C(y_1_delay[0]), 
         .Z(n33823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15439_3_lut.init = 16'hcaca;
    LUT4 i15036_3_lut (.A(\result_i[16] [12]), .B(\result_i[17] [12]), .C(y_1_delay[0]), 
         .Z(n33420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15036_3_lut.init = 16'hcaca;
    LUT4 i15438_3_lut (.A(\result_r[14] [14]), .B(\result_r[15] [14]), .C(y_1_delay[0]), 
         .Z(n33822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15438_3_lut.init = 16'hcaca;
    PFUMX i15203 (.BLUT(n33575), .ALUT(n33576), .C0(y_1_delay[1]), .Z(n33587));
    LUT4 i2550_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[503])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2550_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15437_3_lut (.A(\result_r[12] [14]), .B(\result_r[13] [14]), .C(y_1_delay[0]), 
         .Z(n33821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15437_3_lut.init = 16'hcaca;
    LUT4 i15035_3_lut (.A(\result_i[14] [12]), .B(\result_i[15] [12]), .C(y_1_delay[0]), 
         .Z(n33419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15035_3_lut.init = 16'hcaca;
    LUT4 i2542_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[504])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2542_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15436_3_lut (.A(\result_r[10] [14]), .B(\result_r[11] [14]), .C(y_1_delay[0]), 
         .Z(n33820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15436_3_lut.init = 16'hcaca;
    LUT4 i15034_3_lut (.A(\result_i[12] [12]), .B(\result_i[13] [12]), .C(y_1_delay[0]), 
         .Z(n33418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15034_3_lut.init = 16'hcaca;
    LUT4 i15435_3_lut (.A(\result_r[8] [14]), .B(\result_r[9] [14]), .C(y_1_delay[0]), 
         .Z(n33819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15435_3_lut.init = 16'hcaca;
    FD1P3AX dout_i_i0_i3 (.D(next_dout_i_15__N_1045[2]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_2));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i3.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i4 (.D(next_dout_i_15__N_1045[3]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_3));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i4.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i5 (.D(next_dout_i_15__N_1045[4]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_4));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i5.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i6 (.D(next_dout_i_15__N_1045[5]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_5));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i6.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i7 (.D(next_dout_i_15__N_1045[6]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_6));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i7.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i8 (.D(next_dout_i_15__N_1045[7]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_7));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i8.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i9 (.D(next_dout_i_15__N_1045[8]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_8));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i9.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i10 (.D(next_dout_i_15__N_1045[9]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_9));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i10.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i11 (.D(next_dout_i_15__N_1045[10]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_10));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i11.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i12 (.D(next_dout_i_15__N_1045[11]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_11));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i12.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i13 (.D(next_dout_i_15__N_1045[12]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_12));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i13.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i14 (.D(next_dout_i_15__N_1045[13]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_13));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i14.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i15 (.D(next_dout_i_15__N_1045[14]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_14));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i15.GSR = "ENABLED";
    FD1P3AX dout_i_i0_i16 (.D(next_dout_i_15__N_1045[15]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_i_c_15));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_i_i0_i16.GSR = "ENABLED";
    FD1P3AX result_r_31___i2 (.D(result_r_ns_0__15__N_3[1]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i2.GSR = "ENABLED";
    LUT4 i15601_3_lut (.A(\result_r[30] [9]), .B(\result_r[31] [9]), .C(y_1_delay[0]), 
         .Z(n33985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15601_3_lut.init = 16'hcaca;
    LUT4 i15600_3_lut (.A(\result_r[28] [9]), .B(\result_r[29] [9]), .C(y_1_delay[0]), 
         .Z(n33984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15600_3_lut.init = 16'hcaca;
    LUT4 i15434_3_lut (.A(\result_r[6] [14]), .B(\result_r[7] [14]), .C(y_1_delay[0]), 
         .Z(n33818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15434_3_lut.init = 16'hcaca;
    LUT4 i15433_3_lut (.A(\result_r[4] [14]), .B(\result_r[5] [14]), .C(y_1_delay[0]), 
         .Z(n33817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15433_3_lut.init = 16'hcaca;
    LUT4 i15105_3_lut (.A(\result_i[30] [10]), .B(\result_i[31] [10]), .C(y_1_delay[0]), 
         .Z(n33489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15105_3_lut.init = 16'hcaca;
    LUT4 i15104_3_lut (.A(\result_i[28] [10]), .B(\result_i[29] [10]), .C(y_1_delay[0]), 
         .Z(n33488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15104_3_lut.init = 16'hcaca;
    FD1P3AX result_r_31___i3 (.D(result_r_ns_0__15__N_3[2]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i3.GSR = "ENABLED";
    FD1P3AX result_r_31___i4 (.D(result_r_ns_0__15__N_3[3]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i4.GSR = "ENABLED";
    FD1P3AX result_r_31___i5 (.D(result_r_ns_0__15__N_3[4]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i5.GSR = "ENABLED";
    FD1P3AX result_r_31___i6 (.D(result_r_ns_0__15__N_3[5]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i6.GSR = "ENABLED";
    FD1P3AX result_r_31___i7 (.D(result_r_ns_0__15__N_3[6]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i7.GSR = "ENABLED";
    FD1P3AX result_r_31___i8 (.D(result_r_ns_0__15__N_3[7]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i8.GSR = "ENABLED";
    FD1P3AX result_r_31___i9 (.D(result_r_ns_0__15__N_3[8]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i9.GSR = "ENABLED";
    FD1P3AX result_r_31___i10 (.D(result_r_ns_0__15__N_3[9]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i10.GSR = "ENABLED";
    FD1P3AX result_r_31___i11 (.D(result_r_ns_0__15__N_3[10]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i11.GSR = "ENABLED";
    FD1P3AX result_r_31___i12 (.D(result_r_ns_0__15__N_3[11]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i12.GSR = "ENABLED";
    FD1P3AX result_r_31___i13 (.D(result_r_ns_0__15__N_3[12]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i13.GSR = "ENABLED";
    FD1P3AX result_r_31___i14 (.D(result_r_ns_0__15__N_3[13]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i14.GSR = "ENABLED";
    FD1P3AX result_r_31___i15 (.D(result_r_ns_0__15__N_3[14]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i15.GSR = "ENABLED";
    FD1P3AX result_r_31___i16 (.D(result_r_ns_0__15__N_3[15]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[31] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i16.GSR = "ENABLED";
    FD1P3AX result_r_31___i17 (.D(result_r_ns_0__15__N_3[16]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i17.GSR = "ENABLED";
    FD1P3AX result_r_31___i18 (.D(result_r_ns_0__15__N_3[17]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i18.GSR = "ENABLED";
    FD1P3AX result_r_31___i19 (.D(result_r_ns_0__15__N_3[18]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i19.GSR = "ENABLED";
    FD1P3AX result_r_31___i20 (.D(result_r_ns_0__15__N_3[19]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i20.GSR = "ENABLED";
    FD1P3AX result_r_31___i21 (.D(result_r_ns_0__15__N_3[20]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i21.GSR = "ENABLED";
    FD1P3AX result_r_31___i22 (.D(result_r_ns_0__15__N_3[21]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i22.GSR = "ENABLED";
    FD1P3AX result_r_31___i23 (.D(result_r_ns_0__15__N_3[22]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i23.GSR = "ENABLED";
    FD1P3AX result_r_31___i24 (.D(result_r_ns_0__15__N_3[23]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i24.GSR = "ENABLED";
    FD1P3AX result_r_31___i25 (.D(result_r_ns_0__15__N_3[24]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i25.GSR = "ENABLED";
    FD1P3AX result_r_31___i26 (.D(result_r_ns_0__15__N_3[25]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i26.GSR = "ENABLED";
    FD1P3AX result_r_31___i27 (.D(result_r_ns_0__15__N_3[26]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i27.GSR = "ENABLED";
    FD1P3AX result_r_31___i28 (.D(result_r_ns_0__15__N_3[27]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i28.GSR = "ENABLED";
    FD1P3AX result_r_31___i29 (.D(result_r_ns_0__15__N_3[28]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i29.GSR = "ENABLED";
    FD1P3AX result_r_31___i30 (.D(result_r_ns_0__15__N_3[29]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i30.GSR = "ENABLED";
    FD1P3AX result_r_31___i31 (.D(result_r_ns_0__15__N_3[30]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i31.GSR = "ENABLED";
    FD1P3AX result_r_31___i32 (.D(result_r_ns_0__15__N_3[31]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[30] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i32.GSR = "ENABLED";
    FD1P3AX result_r_31___i33 (.D(result_r_ns_0__15__N_3[32]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i33.GSR = "ENABLED";
    FD1P3AX result_r_31___i34 (.D(result_r_ns_0__15__N_3[33]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i34.GSR = "ENABLED";
    FD1P3AX result_r_31___i35 (.D(result_r_ns_0__15__N_3[34]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i35.GSR = "ENABLED";
    FD1P3AX result_r_31___i36 (.D(result_r_ns_0__15__N_3[35]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i36.GSR = "ENABLED";
    FD1P3AX result_r_31___i37 (.D(result_r_ns_0__15__N_3[36]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i37.GSR = "ENABLED";
    FD1P3AX result_r_31___i38 (.D(result_r_ns_0__15__N_3[37]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i38.GSR = "ENABLED";
    FD1P3AX result_r_31___i39 (.D(result_r_ns_0__15__N_3[38]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i39.GSR = "ENABLED";
    FD1P3AX result_r_31___i40 (.D(result_r_ns_0__15__N_3[39]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i40.GSR = "ENABLED";
    FD1P3AX result_r_31___i41 (.D(result_r_ns_0__15__N_3[40]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i41.GSR = "ENABLED";
    FD1P3AX result_r_31___i42 (.D(result_r_ns_0__15__N_3[41]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i42.GSR = "ENABLED";
    FD1P3AX result_r_31___i43 (.D(result_r_ns_0__15__N_3[42]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i43.GSR = "ENABLED";
    FD1P3AX result_r_31___i44 (.D(result_r_ns_0__15__N_3[43]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i44.GSR = "ENABLED";
    FD1P3AX result_r_31___i45 (.D(result_r_ns_0__15__N_3[44]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i45.GSR = "ENABLED";
    FD1P3AX result_r_31___i46 (.D(result_r_ns_0__15__N_3[45]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i46.GSR = "ENABLED";
    FD1P3AX result_r_31___i47 (.D(result_r_ns_0__15__N_3[46]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i47.GSR = "ENABLED";
    FD1P3AX result_r_31___i48 (.D(result_r_ns_0__15__N_3[47]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[29] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i48.GSR = "ENABLED";
    FD1P3AX result_r_31___i49 (.D(result_r_ns_0__15__N_3[48]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i49.GSR = "ENABLED";
    FD1P3AX result_r_31___i50 (.D(result_r_ns_0__15__N_3[49]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i50.GSR = "ENABLED";
    FD1P3AX result_r_31___i51 (.D(result_r_ns_0__15__N_3[50]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i51.GSR = "ENABLED";
    FD1P3AX result_r_31___i52 (.D(result_r_ns_0__15__N_3[51]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i52.GSR = "ENABLED";
    FD1P3AX result_r_31___i53 (.D(result_r_ns_0__15__N_3[52]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i53.GSR = "ENABLED";
    FD1P3AX result_r_31___i54 (.D(result_r_ns_0__15__N_3[53]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i54.GSR = "ENABLED";
    FD1P3AX result_r_31___i55 (.D(result_r_ns_0__15__N_3[54]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i55.GSR = "ENABLED";
    FD1P3AX result_r_31___i56 (.D(result_r_ns_0__15__N_3[55]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i56.GSR = "ENABLED";
    FD1P3AX result_r_31___i57 (.D(result_r_ns_0__15__N_3[56]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i57.GSR = "ENABLED";
    FD1P3AX result_r_31___i58 (.D(result_r_ns_0__15__N_3[57]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i58.GSR = "ENABLED";
    FD1P3AX result_r_31___i59 (.D(result_r_ns_0__15__N_3[58]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i59.GSR = "ENABLED";
    FD1P3AX result_r_31___i60 (.D(result_r_ns_0__15__N_3[59]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i60.GSR = "ENABLED";
    FD1P3AX result_r_31___i61 (.D(result_r_ns_0__15__N_3[60]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i61.GSR = "ENABLED";
    FD1P3AX result_r_31___i62 (.D(result_r_ns_0__15__N_3[61]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i62.GSR = "ENABLED";
    FD1P3AX result_r_31___i63 (.D(result_r_ns_0__15__N_3[62]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i63.GSR = "ENABLED";
    FD1P3AX result_r_31___i64 (.D(result_r_ns_0__15__N_3[63]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[28] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i64.GSR = "ENABLED";
    FD1P3AX result_r_31___i65 (.D(result_r_ns_0__15__N_3[64]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i65.GSR = "ENABLED";
    FD1P3AX result_r_31___i66 (.D(result_r_ns_0__15__N_3[65]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i66.GSR = "ENABLED";
    FD1P3AX result_r_31___i67 (.D(result_r_ns_0__15__N_3[66]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i67.GSR = "ENABLED";
    FD1P3AX result_r_31___i68 (.D(result_r_ns_0__15__N_3[67]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i68.GSR = "ENABLED";
    FD1P3AX result_r_31___i69 (.D(result_r_ns_0__15__N_3[68]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i69.GSR = "ENABLED";
    FD1P3AX result_r_31___i70 (.D(result_r_ns_0__15__N_3[69]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i70.GSR = "ENABLED";
    FD1P3AX result_r_31___i71 (.D(result_r_ns_0__15__N_3[70]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i71.GSR = "ENABLED";
    FD1P3AX result_r_31___i72 (.D(result_r_ns_0__15__N_3[71]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i72.GSR = "ENABLED";
    FD1P3AX result_r_31___i73 (.D(result_r_ns_0__15__N_3[72]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i73.GSR = "ENABLED";
    FD1P3AX result_r_31___i74 (.D(result_r_ns_0__15__N_3[73]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i74.GSR = "ENABLED";
    FD1P3AX result_r_31___i75 (.D(result_r_ns_0__15__N_3[74]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i75.GSR = "ENABLED";
    FD1P3AX result_r_31___i76 (.D(result_r_ns_0__15__N_3[75]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i76.GSR = "ENABLED";
    FD1P3AX result_r_31___i77 (.D(result_r_ns_0__15__N_3[76]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i77.GSR = "ENABLED";
    FD1P3AX result_r_31___i78 (.D(result_r_ns_0__15__N_3[77]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i78.GSR = "ENABLED";
    FD1P3AX result_r_31___i79 (.D(result_r_ns_0__15__N_3[78]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i79.GSR = "ENABLED";
    FD1P3AX result_r_31___i80 (.D(result_r_ns_0__15__N_3[79]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[27] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i80.GSR = "ENABLED";
    FD1P3AX result_r_31___i81 (.D(result_r_ns_0__15__N_3[80]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i81.GSR = "ENABLED";
    FD1P3AX result_r_31___i82 (.D(result_r_ns_0__15__N_3[81]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i82.GSR = "ENABLED";
    FD1P3AX result_r_31___i83 (.D(result_r_ns_0__15__N_3[82]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i83.GSR = "ENABLED";
    FD1P3AX result_r_31___i84 (.D(result_r_ns_0__15__N_3[83]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i84.GSR = "ENABLED";
    FD1P3AX result_r_31___i85 (.D(result_r_ns_0__15__N_3[84]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i85.GSR = "ENABLED";
    FD1P3AX result_r_31___i86 (.D(result_r_ns_0__15__N_3[85]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i86.GSR = "ENABLED";
    FD1P3AX result_r_31___i87 (.D(result_r_ns_0__15__N_3[86]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i87.GSR = "ENABLED";
    FD1P3AX result_r_31___i88 (.D(result_r_ns_0__15__N_3[87]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i88.GSR = "ENABLED";
    FD1P3AX result_r_31___i89 (.D(result_r_ns_0__15__N_3[88]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i89.GSR = "ENABLED";
    FD1P3AX result_r_31___i90 (.D(result_r_ns_0__15__N_3[89]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i90.GSR = "ENABLED";
    FD1P3AX result_r_31___i91 (.D(result_r_ns_0__15__N_3[90]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i91.GSR = "ENABLED";
    FD1P3AX result_r_31___i92 (.D(result_r_ns_0__15__N_3[91]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i92.GSR = "ENABLED";
    FD1P3AX result_r_31___i93 (.D(result_r_ns_0__15__N_3[92]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i93.GSR = "ENABLED";
    FD1P3AX result_r_31___i94 (.D(result_r_ns_0__15__N_3[93]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i94.GSR = "ENABLED";
    FD1P3AX result_r_31___i95 (.D(result_r_ns_0__15__N_3[94]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i95.GSR = "ENABLED";
    FD1P3AX result_r_31___i96 (.D(result_r_ns_0__15__N_3[95]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[26] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i96.GSR = "ENABLED";
    FD1P3AX result_r_31___i97 (.D(result_r_ns_0__15__N_3[96]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i97.GSR = "ENABLED";
    FD1P3AX result_r_31___i98 (.D(result_r_ns_0__15__N_3[97]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i98.GSR = "ENABLED";
    FD1P3AX result_r_31___i99 (.D(result_r_ns_0__15__N_3[98]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i99.GSR = "ENABLED";
    FD1P3AX result_r_31___i100 (.D(result_r_ns_0__15__N_3[99]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i100.GSR = "ENABLED";
    FD1P3AX result_r_31___i101 (.D(result_r_ns_0__15__N_3[100]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i101.GSR = "ENABLED";
    FD1P3AX result_r_31___i102 (.D(result_r_ns_0__15__N_3[101]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i102.GSR = "ENABLED";
    FD1P3AX result_r_31___i103 (.D(result_r_ns_0__15__N_3[102]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i103.GSR = "ENABLED";
    FD1P3AX result_r_31___i104 (.D(result_r_ns_0__15__N_3[103]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i104.GSR = "ENABLED";
    FD1P3AX result_r_31___i105 (.D(result_r_ns_0__15__N_3[104]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i105.GSR = "ENABLED";
    FD1P3AX result_r_31___i106 (.D(result_r_ns_0__15__N_3[105]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i106.GSR = "ENABLED";
    FD1P3AX result_r_31___i107 (.D(result_r_ns_0__15__N_3[106]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i107.GSR = "ENABLED";
    FD1P3AX result_r_31___i108 (.D(result_r_ns_0__15__N_3[107]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i108.GSR = "ENABLED";
    FD1P3AX result_r_31___i109 (.D(result_r_ns_0__15__N_3[108]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i109.GSR = "ENABLED";
    FD1P3AX result_r_31___i110 (.D(result_r_ns_0__15__N_3[109]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i110.GSR = "ENABLED";
    FD1P3AX result_r_31___i111 (.D(result_r_ns_0__15__N_3[110]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i111.GSR = "ENABLED";
    FD1P3AX result_r_31___i112 (.D(result_r_ns_0__15__N_3[111]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[25] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i112.GSR = "ENABLED";
    FD1P3AX result_r_31___i113 (.D(result_r_ns_0__15__N_3[112]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i113.GSR = "ENABLED";
    FD1P3AX result_r_31___i114 (.D(result_r_ns_0__15__N_3[113]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i114.GSR = "ENABLED";
    FD1P3AX result_r_31___i115 (.D(result_r_ns_0__15__N_3[114]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i115.GSR = "ENABLED";
    FD1P3AX result_r_31___i116 (.D(result_r_ns_0__15__N_3[115]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i116.GSR = "ENABLED";
    FD1P3AX result_r_31___i117 (.D(result_r_ns_0__15__N_3[116]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i117.GSR = "ENABLED";
    FD1P3AX result_r_31___i118 (.D(result_r_ns_0__15__N_3[117]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i118.GSR = "ENABLED";
    FD1P3AX result_r_31___i119 (.D(result_r_ns_0__15__N_3[118]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i119.GSR = "ENABLED";
    FD1P3AX result_r_31___i120 (.D(result_r_ns_0__15__N_3[119]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i120.GSR = "ENABLED";
    FD1P3AX result_r_31___i121 (.D(result_r_ns_0__15__N_3[120]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i121.GSR = "ENABLED";
    FD1P3AX result_r_31___i122 (.D(result_r_ns_0__15__N_3[121]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i122.GSR = "ENABLED";
    FD1P3AX result_r_31___i123 (.D(result_r_ns_0__15__N_3[122]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i123.GSR = "ENABLED";
    FD1P3AX result_r_31___i124 (.D(result_r_ns_0__15__N_3[123]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i124.GSR = "ENABLED";
    FD1P3AX result_r_31___i125 (.D(result_r_ns_0__15__N_3[124]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i125.GSR = "ENABLED";
    FD1P3AX result_r_31___i126 (.D(result_r_ns_0__15__N_3[125]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i126.GSR = "ENABLED";
    FD1P3AX result_r_31___i127 (.D(result_r_ns_0__15__N_3[126]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i127.GSR = "ENABLED";
    FD1P3AX result_r_31___i128 (.D(result_r_ns_0__15__N_3[127]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[24] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i128.GSR = "ENABLED";
    FD1P3AX result_r_31___i129 (.D(result_r_ns_0__15__N_3[128]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i129.GSR = "ENABLED";
    FD1P3AX result_r_31___i130 (.D(result_r_ns_0__15__N_3[129]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i130.GSR = "ENABLED";
    FD1P3AX result_r_31___i131 (.D(result_r_ns_0__15__N_3[130]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i131.GSR = "ENABLED";
    FD1P3AX result_r_31___i132 (.D(result_r_ns_0__15__N_3[131]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i132.GSR = "ENABLED";
    FD1P3AX result_r_31___i133 (.D(result_r_ns_0__15__N_3[132]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i133.GSR = "ENABLED";
    FD1P3AX result_r_31___i134 (.D(result_r_ns_0__15__N_3[133]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i134.GSR = "ENABLED";
    FD1P3AX result_r_31___i135 (.D(result_r_ns_0__15__N_3[134]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i135.GSR = "ENABLED";
    FD1P3AX result_r_31___i136 (.D(result_r_ns_0__15__N_3[135]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i136.GSR = "ENABLED";
    FD1P3AX result_r_31___i137 (.D(result_r_ns_0__15__N_3[136]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i137.GSR = "ENABLED";
    FD1P3AX result_r_31___i138 (.D(result_r_ns_0__15__N_3[137]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i138.GSR = "ENABLED";
    FD1P3AX result_r_31___i139 (.D(result_r_ns_0__15__N_3[138]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i139.GSR = "ENABLED";
    FD1P3AX result_r_31___i140 (.D(result_r_ns_0__15__N_3[139]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i140.GSR = "ENABLED";
    FD1P3AX result_r_31___i141 (.D(result_r_ns_0__15__N_3[140]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i141.GSR = "ENABLED";
    FD1P3AX result_r_31___i142 (.D(result_r_ns_0__15__N_3[141]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i142.GSR = "ENABLED";
    FD1P3AX result_r_31___i143 (.D(result_r_ns_0__15__N_3[142]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i143.GSR = "ENABLED";
    FD1P3AX result_r_31___i144 (.D(result_r_ns_0__15__N_3[143]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[23] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i144.GSR = "ENABLED";
    FD1P3AX result_r_31___i145 (.D(result_r_ns_0__15__N_3[144]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i145.GSR = "ENABLED";
    FD1P3AX result_r_31___i146 (.D(result_r_ns_0__15__N_3[145]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i146.GSR = "ENABLED";
    FD1P3AX result_r_31___i147 (.D(result_r_ns_0__15__N_3[146]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i147.GSR = "ENABLED";
    FD1P3AX result_r_31___i148 (.D(result_r_ns_0__15__N_3[147]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i148.GSR = "ENABLED";
    FD1P3AX result_r_31___i149 (.D(result_r_ns_0__15__N_3[148]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i149.GSR = "ENABLED";
    FD1P3AX result_r_31___i150 (.D(result_r_ns_0__15__N_3[149]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i150.GSR = "ENABLED";
    FD1P3AX result_r_31___i151 (.D(result_r_ns_0__15__N_3[150]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i151.GSR = "ENABLED";
    FD1P3AX result_r_31___i152 (.D(result_r_ns_0__15__N_3[151]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i152.GSR = "ENABLED";
    FD1P3AX result_r_31___i153 (.D(result_r_ns_0__15__N_3[152]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i153.GSR = "ENABLED";
    FD1P3AX result_r_31___i154 (.D(result_r_ns_0__15__N_3[153]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i154.GSR = "ENABLED";
    FD1P3AX result_r_31___i155 (.D(result_r_ns_0__15__N_3[154]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i155.GSR = "ENABLED";
    FD1P3AX result_r_31___i156 (.D(result_r_ns_0__15__N_3[155]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i156.GSR = "ENABLED";
    FD1P3AX result_r_31___i157 (.D(result_r_ns_0__15__N_3[156]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i157.GSR = "ENABLED";
    FD1P3AX result_r_31___i158 (.D(result_r_ns_0__15__N_3[157]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i158.GSR = "ENABLED";
    FD1P3AX result_r_31___i159 (.D(result_r_ns_0__15__N_3[158]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i159.GSR = "ENABLED";
    FD1P3AX result_r_31___i160 (.D(result_r_ns_0__15__N_3[159]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[22] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i160.GSR = "ENABLED";
    FD1P3AX result_r_31___i161 (.D(result_r_ns_0__15__N_3[160]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i161.GSR = "ENABLED";
    FD1P3AX result_r_31___i162 (.D(result_r_ns_0__15__N_3[161]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i162.GSR = "ENABLED";
    FD1P3AX result_r_31___i163 (.D(result_r_ns_0__15__N_3[162]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i163.GSR = "ENABLED";
    FD1P3AX result_r_31___i164 (.D(result_r_ns_0__15__N_3[163]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i164.GSR = "ENABLED";
    FD1P3AX result_r_31___i165 (.D(result_r_ns_0__15__N_3[164]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i165.GSR = "ENABLED";
    FD1P3AX result_r_31___i166 (.D(result_r_ns_0__15__N_3[165]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i166.GSR = "ENABLED";
    FD1P3AX result_r_31___i167 (.D(result_r_ns_0__15__N_3[166]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i167.GSR = "ENABLED";
    FD1P3AX result_r_31___i168 (.D(result_r_ns_0__15__N_3[167]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i168.GSR = "ENABLED";
    FD1P3AX result_r_31___i169 (.D(result_r_ns_0__15__N_3[168]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i169.GSR = "ENABLED";
    FD1P3AX result_r_31___i170 (.D(result_r_ns_0__15__N_3[169]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i170.GSR = "ENABLED";
    FD1P3AX result_r_31___i171 (.D(result_r_ns_0__15__N_3[170]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i171.GSR = "ENABLED";
    FD1P3AX result_r_31___i172 (.D(result_r_ns_0__15__N_3[171]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i172.GSR = "ENABLED";
    FD1P3AX result_r_31___i173 (.D(result_r_ns_0__15__N_3[172]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i173.GSR = "ENABLED";
    FD1P3AX result_r_31___i174 (.D(result_r_ns_0__15__N_3[173]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i174.GSR = "ENABLED";
    FD1P3AX result_r_31___i175 (.D(result_r_ns_0__15__N_3[174]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i175.GSR = "ENABLED";
    FD1P3AX result_r_31___i176 (.D(result_r_ns_0__15__N_3[175]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[21] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i176.GSR = "ENABLED";
    FD1P3AX result_r_31___i177 (.D(result_r_ns_0__15__N_3[176]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i177.GSR = "ENABLED";
    FD1P3AX result_r_31___i178 (.D(result_r_ns_0__15__N_3[177]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i178.GSR = "ENABLED";
    FD1P3AX result_r_31___i179 (.D(result_r_ns_0__15__N_3[178]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i179.GSR = "ENABLED";
    FD1P3AX result_r_31___i180 (.D(result_r_ns_0__15__N_3[179]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i180.GSR = "ENABLED";
    FD1P3AX result_r_31___i181 (.D(result_r_ns_0__15__N_3[180]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i181.GSR = "ENABLED";
    FD1P3AX result_r_31___i182 (.D(result_r_ns_0__15__N_3[181]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i182.GSR = "ENABLED";
    FD1P3AX result_r_31___i183 (.D(result_r_ns_0__15__N_3[182]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i183.GSR = "ENABLED";
    FD1P3AX result_r_31___i184 (.D(result_r_ns_0__15__N_3[183]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i184.GSR = "ENABLED";
    FD1P3AX result_r_31___i185 (.D(result_r_ns_0__15__N_3[184]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i185.GSR = "ENABLED";
    FD1P3AX result_r_31___i186 (.D(result_r_ns_0__15__N_3[185]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i186.GSR = "ENABLED";
    FD1P3AX result_r_31___i187 (.D(result_r_ns_0__15__N_3[186]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i187.GSR = "ENABLED";
    FD1P3AX result_r_31___i188 (.D(result_r_ns_0__15__N_3[187]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i188.GSR = "ENABLED";
    FD1P3AX result_r_31___i189 (.D(result_r_ns_0__15__N_3[188]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i189.GSR = "ENABLED";
    FD1P3AX result_r_31___i190 (.D(result_r_ns_0__15__N_3[189]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i190.GSR = "ENABLED";
    FD1P3AX result_r_31___i191 (.D(result_r_ns_0__15__N_3[190]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i191.GSR = "ENABLED";
    FD1P3AX result_r_31___i192 (.D(result_r_ns_0__15__N_3[191]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[20] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i192.GSR = "ENABLED";
    FD1P3AX result_r_31___i193 (.D(result_r_ns_0__15__N_3[192]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i193.GSR = "ENABLED";
    FD1P3AX result_r_31___i194 (.D(result_r_ns_0__15__N_3[193]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i194.GSR = "ENABLED";
    FD1P3AX result_r_31___i195 (.D(result_r_ns_0__15__N_3[194]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i195.GSR = "ENABLED";
    FD1P3AX result_r_31___i196 (.D(result_r_ns_0__15__N_3[195]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i196.GSR = "ENABLED";
    FD1P3AX result_r_31___i197 (.D(result_r_ns_0__15__N_3[196]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i197.GSR = "ENABLED";
    FD1P3AX result_r_31___i198 (.D(result_r_ns_0__15__N_3[197]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i198.GSR = "ENABLED";
    FD1P3AX result_r_31___i199 (.D(result_r_ns_0__15__N_3[198]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i199.GSR = "ENABLED";
    FD1P3AX result_r_31___i200 (.D(result_r_ns_0__15__N_3[199]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i200.GSR = "ENABLED";
    FD1P3AX result_r_31___i201 (.D(result_r_ns_0__15__N_3[200]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i201.GSR = "ENABLED";
    FD1P3AX result_r_31___i202 (.D(result_r_ns_0__15__N_3[201]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i202.GSR = "ENABLED";
    FD1P3AX result_r_31___i203 (.D(result_r_ns_0__15__N_3[202]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i203.GSR = "ENABLED";
    FD1P3AX result_r_31___i204 (.D(result_r_ns_0__15__N_3[203]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i204.GSR = "ENABLED";
    FD1P3AX result_r_31___i205 (.D(result_r_ns_0__15__N_3[204]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i205.GSR = "ENABLED";
    FD1P3AX result_r_31___i206 (.D(result_r_ns_0__15__N_3[205]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i206.GSR = "ENABLED";
    FD1P3AX result_r_31___i207 (.D(result_r_ns_0__15__N_3[206]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i207.GSR = "ENABLED";
    FD1P3AX result_r_31___i208 (.D(result_r_ns_0__15__N_3[207]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[19] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i208.GSR = "ENABLED";
    FD1P3AX result_r_31___i209 (.D(result_r_ns_0__15__N_3[208]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i209.GSR = "ENABLED";
    FD1P3AX result_r_31___i210 (.D(result_r_ns_0__15__N_3[209]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i210.GSR = "ENABLED";
    FD1P3AX result_r_31___i211 (.D(result_r_ns_0__15__N_3[210]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i211.GSR = "ENABLED";
    FD1P3AX result_r_31___i212 (.D(result_r_ns_0__15__N_3[211]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i212.GSR = "ENABLED";
    FD1P3AX result_r_31___i213 (.D(result_r_ns_0__15__N_3[212]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i213.GSR = "ENABLED";
    FD1P3AX result_r_31___i214 (.D(result_r_ns_0__15__N_3[213]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i214.GSR = "ENABLED";
    FD1P3AX result_r_31___i215 (.D(result_r_ns_0__15__N_3[214]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i215.GSR = "ENABLED";
    FD1P3AX result_r_31___i216 (.D(result_r_ns_0__15__N_3[215]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i216.GSR = "ENABLED";
    FD1P3AX result_r_31___i217 (.D(result_r_ns_0__15__N_3[216]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i217.GSR = "ENABLED";
    FD1P3AX result_r_31___i218 (.D(result_r_ns_0__15__N_3[217]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i218.GSR = "ENABLED";
    FD1P3AX result_r_31___i219 (.D(result_r_ns_0__15__N_3[218]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i219.GSR = "ENABLED";
    FD1P3AX result_r_31___i220 (.D(result_r_ns_0__15__N_3[219]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i220.GSR = "ENABLED";
    FD1P3AX result_r_31___i221 (.D(result_r_ns_0__15__N_3[220]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i221.GSR = "ENABLED";
    FD1P3AX result_r_31___i222 (.D(result_r_ns_0__15__N_3[221]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i222.GSR = "ENABLED";
    FD1P3AX result_r_31___i223 (.D(result_r_ns_0__15__N_3[222]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i223.GSR = "ENABLED";
    FD1P3AX result_r_31___i224 (.D(result_r_ns_0__15__N_3[223]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[18] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i224.GSR = "ENABLED";
    FD1P3AX result_r_31___i225 (.D(result_r_ns_0__15__N_3[224]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i225.GSR = "ENABLED";
    FD1P3AX result_r_31___i226 (.D(result_r_ns_0__15__N_3[225]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i226.GSR = "ENABLED";
    FD1P3AX result_r_31___i227 (.D(result_r_ns_0__15__N_3[226]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i227.GSR = "ENABLED";
    FD1P3AX result_r_31___i228 (.D(result_r_ns_0__15__N_3[227]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i228.GSR = "ENABLED";
    FD1P3AX result_r_31___i229 (.D(result_r_ns_0__15__N_3[228]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i229.GSR = "ENABLED";
    FD1P3AX result_r_31___i230 (.D(result_r_ns_0__15__N_3[229]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i230.GSR = "ENABLED";
    FD1P3AX result_r_31___i231 (.D(result_r_ns_0__15__N_3[230]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i231.GSR = "ENABLED";
    FD1P3AX result_r_31___i232 (.D(result_r_ns_0__15__N_3[231]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i232.GSR = "ENABLED";
    FD1P3AX result_r_31___i233 (.D(result_r_ns_0__15__N_3[232]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i233.GSR = "ENABLED";
    FD1P3AX result_r_31___i234 (.D(result_r_ns_0__15__N_3[233]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i234.GSR = "ENABLED";
    FD1P3AX result_r_31___i235 (.D(result_r_ns_0__15__N_3[234]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i235.GSR = "ENABLED";
    FD1P3AX result_r_31___i236 (.D(result_r_ns_0__15__N_3[235]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i236.GSR = "ENABLED";
    FD1P3AX result_r_31___i237 (.D(result_r_ns_0__15__N_3[236]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i237.GSR = "ENABLED";
    FD1P3AX result_r_31___i238 (.D(result_r_ns_0__15__N_3[237]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i238.GSR = "ENABLED";
    FD1P3AX result_r_31___i239 (.D(result_r_ns_0__15__N_3[238]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i239.GSR = "ENABLED";
    FD1P3AX result_r_31___i240 (.D(result_r_ns_0__15__N_3[239]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[17] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i240.GSR = "ENABLED";
    FD1P3AX result_r_31___i241 (.D(result_r_ns_0__15__N_3[240]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i241.GSR = "ENABLED";
    FD1P3AX result_r_31___i242 (.D(result_r_ns_0__15__N_3[241]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i242.GSR = "ENABLED";
    FD1P3AX result_r_31___i243 (.D(result_r_ns_0__15__N_3[242]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i243.GSR = "ENABLED";
    FD1P3AX result_r_31___i244 (.D(result_r_ns_0__15__N_3[243]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i244.GSR = "ENABLED";
    FD1P3AX result_r_31___i245 (.D(result_r_ns_0__15__N_3[244]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i245.GSR = "ENABLED";
    FD1P3AX result_r_31___i246 (.D(result_r_ns_0__15__N_3[245]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i246.GSR = "ENABLED";
    FD1P3AX result_r_31___i247 (.D(result_r_ns_0__15__N_3[246]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i247.GSR = "ENABLED";
    FD1P3AX result_r_31___i248 (.D(result_r_ns_0__15__N_3[247]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i248.GSR = "ENABLED";
    FD1P3AX result_r_31___i249 (.D(result_r_ns_0__15__N_3[248]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i249.GSR = "ENABLED";
    FD1P3AX result_r_31___i250 (.D(result_r_ns_0__15__N_3[249]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i250.GSR = "ENABLED";
    FD1P3AX result_r_31___i251 (.D(result_r_ns_0__15__N_3[250]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i251.GSR = "ENABLED";
    FD1P3AX result_r_31___i252 (.D(result_r_ns_0__15__N_3[251]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i252.GSR = "ENABLED";
    FD1P3AX result_r_31___i253 (.D(result_r_ns_0__15__N_3[252]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i253.GSR = "ENABLED";
    FD1P3AX result_r_31___i254 (.D(result_r_ns_0__15__N_3[253]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i254.GSR = "ENABLED";
    FD1P3AX result_r_31___i255 (.D(result_r_ns_0__15__N_3[254]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i255.GSR = "ENABLED";
    FD1P3AX result_r_31___i256 (.D(result_r_ns_0__15__N_3[255]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[16] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i256.GSR = "ENABLED";
    FD1P3AX result_r_31___i257 (.D(result_r_ns_0__15__N_3[256]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i257.GSR = "ENABLED";
    FD1P3AX result_r_31___i258 (.D(result_r_ns_0__15__N_3[257]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i258.GSR = "ENABLED";
    FD1P3AX result_r_31___i259 (.D(result_r_ns_0__15__N_3[258]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i259.GSR = "ENABLED";
    FD1P3AX result_r_31___i260 (.D(result_r_ns_0__15__N_3[259]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i260.GSR = "ENABLED";
    FD1P3AX result_r_31___i261 (.D(result_r_ns_0__15__N_3[260]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i261.GSR = "ENABLED";
    FD1P3AX result_r_31___i262 (.D(result_r_ns_0__15__N_3[261]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i262.GSR = "ENABLED";
    FD1P3AX result_r_31___i263 (.D(result_r_ns_0__15__N_3[262]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i263.GSR = "ENABLED";
    FD1P3AX result_r_31___i264 (.D(result_r_ns_0__15__N_3[263]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i264.GSR = "ENABLED";
    FD1P3AX result_r_31___i265 (.D(result_r_ns_0__15__N_3[264]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i265.GSR = "ENABLED";
    FD1P3AX result_r_31___i266 (.D(result_r_ns_0__15__N_3[265]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i266.GSR = "ENABLED";
    FD1P3AX result_r_31___i267 (.D(result_r_ns_0__15__N_3[266]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i267.GSR = "ENABLED";
    FD1P3AX result_r_31___i268 (.D(result_r_ns_0__15__N_3[267]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i268.GSR = "ENABLED";
    FD1P3AX result_r_31___i269 (.D(result_r_ns_0__15__N_3[268]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i269.GSR = "ENABLED";
    FD1P3AX result_r_31___i270 (.D(result_r_ns_0__15__N_3[269]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i270.GSR = "ENABLED";
    FD1P3AX result_r_31___i271 (.D(result_r_ns_0__15__N_3[270]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i271.GSR = "ENABLED";
    FD1P3AX result_r_31___i272 (.D(result_r_ns_0__15__N_3[271]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[15] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i272.GSR = "ENABLED";
    FD1P3AX result_r_31___i273 (.D(result_r_ns_0__15__N_3[272]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i273.GSR = "ENABLED";
    FD1P3AX result_r_31___i274 (.D(result_r_ns_0__15__N_3[273]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i274.GSR = "ENABLED";
    FD1P3AX result_r_31___i275 (.D(result_r_ns_0__15__N_3[274]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i275.GSR = "ENABLED";
    FD1P3AX result_r_31___i276 (.D(result_r_ns_0__15__N_3[275]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i276.GSR = "ENABLED";
    FD1P3AX result_r_31___i277 (.D(result_r_ns_0__15__N_3[276]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i277.GSR = "ENABLED";
    FD1P3AX result_r_31___i278 (.D(result_r_ns_0__15__N_3[277]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i278.GSR = "ENABLED";
    FD1P3AX result_r_31___i279 (.D(result_r_ns_0__15__N_3[278]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i279.GSR = "ENABLED";
    FD1P3AX result_r_31___i280 (.D(result_r_ns_0__15__N_3[279]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i280.GSR = "ENABLED";
    FD1P3AX result_r_31___i281 (.D(result_r_ns_0__15__N_3[280]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i281.GSR = "ENABLED";
    FD1P3AX result_r_31___i282 (.D(result_r_ns_0__15__N_3[281]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i282.GSR = "ENABLED";
    FD1P3AX result_r_31___i283 (.D(result_r_ns_0__15__N_3[282]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i283.GSR = "ENABLED";
    FD1P3AX result_r_31___i284 (.D(result_r_ns_0__15__N_3[283]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i284.GSR = "ENABLED";
    FD1P3AX result_r_31___i285 (.D(result_r_ns_0__15__N_3[284]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i285.GSR = "ENABLED";
    FD1P3AX result_r_31___i286 (.D(result_r_ns_0__15__N_3[285]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i286.GSR = "ENABLED";
    FD1P3AX result_r_31___i287 (.D(result_r_ns_0__15__N_3[286]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i287.GSR = "ENABLED";
    FD1P3AX result_r_31___i288 (.D(result_r_ns_0__15__N_3[287]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[14] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i288.GSR = "ENABLED";
    FD1P3AX result_r_31___i289 (.D(result_r_ns_0__15__N_3[288]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i289.GSR = "ENABLED";
    FD1P3AX result_r_31___i290 (.D(result_r_ns_0__15__N_3[289]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i290.GSR = "ENABLED";
    FD1P3AX result_r_31___i291 (.D(result_r_ns_0__15__N_3[290]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i291.GSR = "ENABLED";
    FD1P3AX result_r_31___i292 (.D(result_r_ns_0__15__N_3[291]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i292.GSR = "ENABLED";
    FD1P3AX result_r_31___i293 (.D(result_r_ns_0__15__N_3[292]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i293.GSR = "ENABLED";
    FD1P3AX result_r_31___i294 (.D(result_r_ns_0__15__N_3[293]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i294.GSR = "ENABLED";
    FD1P3AX result_r_31___i295 (.D(result_r_ns_0__15__N_3[294]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i295.GSR = "ENABLED";
    FD1P3AX result_r_31___i296 (.D(result_r_ns_0__15__N_3[295]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i296.GSR = "ENABLED";
    FD1P3AX result_r_31___i297 (.D(result_r_ns_0__15__N_3[296]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i297.GSR = "ENABLED";
    FD1P3AX result_r_31___i298 (.D(result_r_ns_0__15__N_3[297]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i298.GSR = "ENABLED";
    FD1P3AX result_r_31___i299 (.D(result_r_ns_0__15__N_3[298]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i299.GSR = "ENABLED";
    FD1P3AX result_r_31___i300 (.D(result_r_ns_0__15__N_3[299]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i300.GSR = "ENABLED";
    FD1P3AX result_r_31___i301 (.D(result_r_ns_0__15__N_3[300]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i301.GSR = "ENABLED";
    FD1P3AX result_r_31___i302 (.D(result_r_ns_0__15__N_3[301]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i302.GSR = "ENABLED";
    FD1P3AX result_r_31___i303 (.D(result_r_ns_0__15__N_3[302]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i303.GSR = "ENABLED";
    FD1P3AX result_r_31___i304 (.D(result_r_ns_0__15__N_3[303]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[13] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i304.GSR = "ENABLED";
    FD1P3AX result_r_31___i305 (.D(result_r_ns_0__15__N_3[304]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i305.GSR = "ENABLED";
    FD1P3AX result_r_31___i306 (.D(result_r_ns_0__15__N_3[305]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i306.GSR = "ENABLED";
    FD1P3AX result_r_31___i307 (.D(result_r_ns_0__15__N_3[306]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i307.GSR = "ENABLED";
    FD1P3AX result_r_31___i308 (.D(result_r_ns_0__15__N_3[307]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i308.GSR = "ENABLED";
    FD1P3AX result_r_31___i309 (.D(result_r_ns_0__15__N_3[308]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i309.GSR = "ENABLED";
    FD1P3AX result_r_31___i310 (.D(result_r_ns_0__15__N_3[309]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i310.GSR = "ENABLED";
    FD1P3AX result_r_31___i311 (.D(result_r_ns_0__15__N_3[310]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i311.GSR = "ENABLED";
    FD1P3AX result_r_31___i312 (.D(result_r_ns_0__15__N_3[311]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i312.GSR = "ENABLED";
    FD1P3AX result_r_31___i313 (.D(result_r_ns_0__15__N_3[312]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i313.GSR = "ENABLED";
    FD1P3AX result_r_31___i314 (.D(result_r_ns_0__15__N_3[313]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i314.GSR = "ENABLED";
    FD1P3AX result_r_31___i315 (.D(result_r_ns_0__15__N_3[314]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i315.GSR = "ENABLED";
    FD1P3AX result_r_31___i316 (.D(result_r_ns_0__15__N_3[315]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i316.GSR = "ENABLED";
    FD1P3AX result_r_31___i317 (.D(result_r_ns_0__15__N_3[316]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i317.GSR = "ENABLED";
    FD1P3AX result_r_31___i318 (.D(result_r_ns_0__15__N_3[317]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i318.GSR = "ENABLED";
    FD1P3AX result_r_31___i319 (.D(result_r_ns_0__15__N_3[318]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i319.GSR = "ENABLED";
    FD1P3AX result_r_31___i320 (.D(result_r_ns_0__15__N_3[319]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[12] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i320.GSR = "ENABLED";
    FD1P3AX result_r_31___i321 (.D(result_r_ns_0__15__N_3[320]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i321.GSR = "ENABLED";
    FD1P3AX result_r_31___i322 (.D(result_r_ns_0__15__N_3[321]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i322.GSR = "ENABLED";
    FD1P3AX result_r_31___i323 (.D(result_r_ns_0__15__N_3[322]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i323.GSR = "ENABLED";
    FD1P3AX result_r_31___i324 (.D(result_r_ns_0__15__N_3[323]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i324.GSR = "ENABLED";
    FD1P3AX result_r_31___i325 (.D(result_r_ns_0__15__N_3[324]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i325.GSR = "ENABLED";
    FD1P3AX result_r_31___i326 (.D(result_r_ns_0__15__N_3[325]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i326.GSR = "ENABLED";
    FD1P3AX result_r_31___i327 (.D(result_r_ns_0__15__N_3[326]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i327.GSR = "ENABLED";
    FD1P3AX result_r_31___i328 (.D(result_r_ns_0__15__N_3[327]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i328.GSR = "ENABLED";
    FD1P3AX result_r_31___i329 (.D(result_r_ns_0__15__N_3[328]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i329.GSR = "ENABLED";
    FD1P3AX result_r_31___i330 (.D(result_r_ns_0__15__N_3[329]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i330.GSR = "ENABLED";
    FD1P3AX result_r_31___i331 (.D(result_r_ns_0__15__N_3[330]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i331.GSR = "ENABLED";
    FD1P3AX result_r_31___i332 (.D(result_r_ns_0__15__N_3[331]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i332.GSR = "ENABLED";
    FD1P3AX result_r_31___i333 (.D(result_r_ns_0__15__N_3[332]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i333.GSR = "ENABLED";
    FD1P3AX result_r_31___i334 (.D(result_r_ns_0__15__N_3[333]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i334.GSR = "ENABLED";
    FD1P3AX result_r_31___i335 (.D(result_r_ns_0__15__N_3[334]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i335.GSR = "ENABLED";
    FD1P3AX result_r_31___i336 (.D(result_r_ns_0__15__N_3[335]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[11] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i336.GSR = "ENABLED";
    FD1P3AX result_r_31___i337 (.D(result_r_ns_0__15__N_3[336]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i337.GSR = "ENABLED";
    FD1P3AX result_r_31___i338 (.D(result_r_ns_0__15__N_3[337]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i338.GSR = "ENABLED";
    FD1P3AX result_r_31___i339 (.D(result_r_ns_0__15__N_3[338]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i339.GSR = "ENABLED";
    FD1P3AX result_r_31___i340 (.D(result_r_ns_0__15__N_3[339]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i340.GSR = "ENABLED";
    FD1P3AX result_r_31___i341 (.D(result_r_ns_0__15__N_3[340]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i341.GSR = "ENABLED";
    FD1P3AX result_r_31___i342 (.D(result_r_ns_0__15__N_3[341]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i342.GSR = "ENABLED";
    FD1P3AX result_r_31___i343 (.D(result_r_ns_0__15__N_3[342]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i343.GSR = "ENABLED";
    FD1P3AX result_r_31___i344 (.D(result_r_ns_0__15__N_3[343]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i344.GSR = "ENABLED";
    FD1P3AX result_r_31___i345 (.D(result_r_ns_0__15__N_3[344]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i345.GSR = "ENABLED";
    FD1P3AX result_r_31___i346 (.D(result_r_ns_0__15__N_3[345]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i346.GSR = "ENABLED";
    FD1P3AX result_r_31___i347 (.D(result_r_ns_0__15__N_3[346]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i347.GSR = "ENABLED";
    FD1P3AX result_r_31___i348 (.D(result_r_ns_0__15__N_3[347]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i348.GSR = "ENABLED";
    FD1P3AX result_r_31___i349 (.D(result_r_ns_0__15__N_3[348]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i349.GSR = "ENABLED";
    FD1P3AX result_r_31___i350 (.D(result_r_ns_0__15__N_3[349]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i350.GSR = "ENABLED";
    FD1P3AX result_r_31___i351 (.D(result_r_ns_0__15__N_3[350]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i351.GSR = "ENABLED";
    FD1P3AX result_r_31___i352 (.D(result_r_ns_0__15__N_3[351]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[10] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i352.GSR = "ENABLED";
    FD1P3AX result_r_31___i353 (.D(result_r_ns_0__15__N_3[352]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i353.GSR = "ENABLED";
    FD1P3AX result_r_31___i354 (.D(result_r_ns_0__15__N_3[353]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i354.GSR = "ENABLED";
    FD1P3AX result_r_31___i355 (.D(result_r_ns_0__15__N_3[354]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i355.GSR = "ENABLED";
    FD1P3AX result_r_31___i356 (.D(result_r_ns_0__15__N_3[355]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i356.GSR = "ENABLED";
    FD1P3AX result_r_31___i357 (.D(result_r_ns_0__15__N_3[356]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i357.GSR = "ENABLED";
    FD1P3AX result_r_31___i358 (.D(result_r_ns_0__15__N_3[357]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i358.GSR = "ENABLED";
    FD1P3AX result_r_31___i359 (.D(result_r_ns_0__15__N_3[358]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i359.GSR = "ENABLED";
    FD1P3AX result_r_31___i360 (.D(result_r_ns_0__15__N_3[359]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i360.GSR = "ENABLED";
    FD1P3AX result_r_31___i361 (.D(result_r_ns_0__15__N_3[360]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i361.GSR = "ENABLED";
    FD1P3AX result_r_31___i362 (.D(result_r_ns_0__15__N_3[361]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i362.GSR = "ENABLED";
    FD1P3AX result_r_31___i363 (.D(result_r_ns_0__15__N_3[362]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i363.GSR = "ENABLED";
    FD1P3AX result_r_31___i364 (.D(result_r_ns_0__15__N_3[363]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i364.GSR = "ENABLED";
    FD1P3AX result_r_31___i365 (.D(result_r_ns_0__15__N_3[364]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i365.GSR = "ENABLED";
    FD1P3AX result_r_31___i366 (.D(result_r_ns_0__15__N_3[365]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i366.GSR = "ENABLED";
    FD1P3AX result_r_31___i367 (.D(result_r_ns_0__15__N_3[366]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i367.GSR = "ENABLED";
    FD1P3AX result_r_31___i368 (.D(result_r_ns_0__15__N_3[367]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[9] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i368.GSR = "ENABLED";
    FD1P3AX result_r_31___i369 (.D(result_r_ns_0__15__N_3[368]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i369.GSR = "ENABLED";
    FD1P3AX result_r_31___i370 (.D(result_r_ns_0__15__N_3[369]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i370.GSR = "ENABLED";
    FD1P3AX result_r_31___i371 (.D(result_r_ns_0__15__N_3[370]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i371.GSR = "ENABLED";
    FD1P3AX result_r_31___i372 (.D(result_r_ns_0__15__N_3[371]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i372.GSR = "ENABLED";
    FD1P3AX result_r_31___i373 (.D(result_r_ns_0__15__N_3[372]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i373.GSR = "ENABLED";
    FD1P3AX result_r_31___i374 (.D(result_r_ns_0__15__N_3[373]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i374.GSR = "ENABLED";
    FD1P3AX result_r_31___i375 (.D(result_r_ns_0__15__N_3[374]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i375.GSR = "ENABLED";
    FD1P3AX result_r_31___i376 (.D(result_r_ns_0__15__N_3[375]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i376.GSR = "ENABLED";
    FD1P3AX result_r_31___i377 (.D(result_r_ns_0__15__N_3[376]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i377.GSR = "ENABLED";
    FD1P3AX result_r_31___i378 (.D(result_r_ns_0__15__N_3[377]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i378.GSR = "ENABLED";
    FD1P3AX result_r_31___i379 (.D(result_r_ns_0__15__N_3[378]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i379.GSR = "ENABLED";
    FD1P3AX result_r_31___i380 (.D(result_r_ns_0__15__N_3[379]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i380.GSR = "ENABLED";
    FD1P3AX result_r_31___i381 (.D(result_r_ns_0__15__N_3[380]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i381.GSR = "ENABLED";
    FD1P3AX result_r_31___i382 (.D(result_r_ns_0__15__N_3[381]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i382.GSR = "ENABLED";
    FD1P3AX result_r_31___i383 (.D(result_r_ns_0__15__N_3[382]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i383.GSR = "ENABLED";
    FD1P3AX result_r_31___i384 (.D(result_r_ns_0__15__N_3[383]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[8] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i384.GSR = "ENABLED";
    FD1P3AX result_r_31___i385 (.D(result_r_ns_0__15__N_3[384]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i385.GSR = "ENABLED";
    FD1P3AX result_r_31___i386 (.D(result_r_ns_0__15__N_3[385]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i386.GSR = "ENABLED";
    FD1P3AX result_r_31___i387 (.D(result_r_ns_0__15__N_3[386]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i387.GSR = "ENABLED";
    FD1P3AX result_r_31___i388 (.D(result_r_ns_0__15__N_3[387]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i388.GSR = "ENABLED";
    FD1P3AX result_r_31___i389 (.D(result_r_ns_0__15__N_3[388]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i389.GSR = "ENABLED";
    FD1P3AX result_r_31___i390 (.D(result_r_ns_0__15__N_3[389]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i390.GSR = "ENABLED";
    FD1P3AX result_r_31___i391 (.D(result_r_ns_0__15__N_3[390]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i391.GSR = "ENABLED";
    FD1P3AX result_r_31___i392 (.D(result_r_ns_0__15__N_3[391]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i392.GSR = "ENABLED";
    FD1P3AX result_r_31___i393 (.D(result_r_ns_0__15__N_3[392]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i393.GSR = "ENABLED";
    FD1P3AX result_r_31___i394 (.D(result_r_ns_0__15__N_3[393]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i394.GSR = "ENABLED";
    FD1P3AX result_r_31___i395 (.D(result_r_ns_0__15__N_3[394]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i395.GSR = "ENABLED";
    FD1P3AX result_r_31___i396 (.D(result_r_ns_0__15__N_3[395]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i396.GSR = "ENABLED";
    FD1P3AX result_r_31___i397 (.D(result_r_ns_0__15__N_3[396]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i397.GSR = "ENABLED";
    FD1P3AX result_r_31___i398 (.D(result_r_ns_0__15__N_3[397]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i398.GSR = "ENABLED";
    FD1P3AX result_r_31___i399 (.D(result_r_ns_0__15__N_3[398]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i399.GSR = "ENABLED";
    FD1P3AX result_r_31___i400 (.D(result_r_ns_0__15__N_3[399]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[7] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i400.GSR = "ENABLED";
    FD1P3AX result_r_31___i401 (.D(result_r_ns_0__15__N_3[400]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i401.GSR = "ENABLED";
    FD1P3AX result_r_31___i402 (.D(result_r_ns_0__15__N_3[401]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i402.GSR = "ENABLED";
    FD1P3AX result_r_31___i403 (.D(result_r_ns_0__15__N_3[402]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i403.GSR = "ENABLED";
    FD1P3AX result_r_31___i404 (.D(result_r_ns_0__15__N_3[403]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i404.GSR = "ENABLED";
    FD1P3AX result_r_31___i405 (.D(result_r_ns_0__15__N_3[404]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i405.GSR = "ENABLED";
    FD1P3AX result_r_31___i406 (.D(result_r_ns_0__15__N_3[405]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i406.GSR = "ENABLED";
    FD1P3AX result_r_31___i407 (.D(result_r_ns_0__15__N_3[406]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i407.GSR = "ENABLED";
    FD1P3AX result_r_31___i408 (.D(result_r_ns_0__15__N_3[407]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i408.GSR = "ENABLED";
    FD1P3AX result_r_31___i409 (.D(result_r_ns_0__15__N_3[408]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i409.GSR = "ENABLED";
    FD1P3AX result_r_31___i410 (.D(result_r_ns_0__15__N_3[409]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i410.GSR = "ENABLED";
    FD1P3AX result_r_31___i411 (.D(result_r_ns_0__15__N_3[410]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i411.GSR = "ENABLED";
    FD1P3AX result_r_31___i412 (.D(result_r_ns_0__15__N_3[411]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i412.GSR = "ENABLED";
    FD1P3AX result_r_31___i413 (.D(result_r_ns_0__15__N_3[412]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i413.GSR = "ENABLED";
    FD1P3AX result_r_31___i414 (.D(result_r_ns_0__15__N_3[413]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i414.GSR = "ENABLED";
    FD1P3AX result_r_31___i415 (.D(result_r_ns_0__15__N_3[414]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i415.GSR = "ENABLED";
    FD1P3AX result_r_31___i416 (.D(result_r_ns_0__15__N_3[415]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[6] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i416.GSR = "ENABLED";
    FD1P3AX result_r_31___i417 (.D(result_r_ns_0__15__N_3[416]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i417.GSR = "ENABLED";
    FD1P3AX result_r_31___i418 (.D(result_r_ns_0__15__N_3[417]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i418.GSR = "ENABLED";
    FD1P3AX result_r_31___i419 (.D(result_r_ns_0__15__N_3[418]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i419.GSR = "ENABLED";
    FD1P3AX result_r_31___i420 (.D(result_r_ns_0__15__N_3[419]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i420.GSR = "ENABLED";
    FD1P3AX result_r_31___i421 (.D(result_r_ns_0__15__N_3[420]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i421.GSR = "ENABLED";
    FD1P3AX result_r_31___i422 (.D(result_r_ns_0__15__N_3[421]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i422.GSR = "ENABLED";
    FD1P3AX result_r_31___i423 (.D(result_r_ns_0__15__N_3[422]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i423.GSR = "ENABLED";
    FD1P3AX result_r_31___i424 (.D(result_r_ns_0__15__N_3[423]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i424.GSR = "ENABLED";
    FD1P3AX result_r_31___i425 (.D(result_r_ns_0__15__N_3[424]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i425.GSR = "ENABLED";
    FD1P3AX result_r_31___i426 (.D(result_r_ns_0__15__N_3[425]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i426.GSR = "ENABLED";
    FD1P3AX result_r_31___i427 (.D(result_r_ns_0__15__N_3[426]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i427.GSR = "ENABLED";
    FD1P3AX result_r_31___i428 (.D(result_r_ns_0__15__N_3[427]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i428.GSR = "ENABLED";
    FD1P3AX result_r_31___i429 (.D(result_r_ns_0__15__N_3[428]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i429.GSR = "ENABLED";
    FD1P3AX result_r_31___i430 (.D(result_r_ns_0__15__N_3[429]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i430.GSR = "ENABLED";
    FD1P3AX result_r_31___i431 (.D(result_r_ns_0__15__N_3[430]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i431.GSR = "ENABLED";
    FD1P3AX result_r_31___i432 (.D(result_r_ns_0__15__N_3[431]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[5] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i432.GSR = "ENABLED";
    FD1P3AX result_r_31___i433 (.D(result_r_ns_0__15__N_3[432]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i433.GSR = "ENABLED";
    FD1P3AX result_r_31___i434 (.D(result_r_ns_0__15__N_3[433]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i434.GSR = "ENABLED";
    FD1P3AX result_r_31___i435 (.D(result_r_ns_0__15__N_3[434]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i435.GSR = "ENABLED";
    FD1P3AX result_r_31___i436 (.D(result_r_ns_0__15__N_3[435]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i436.GSR = "ENABLED";
    FD1P3AX result_r_31___i437 (.D(result_r_ns_0__15__N_3[436]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i437.GSR = "ENABLED";
    FD1P3AX result_r_31___i438 (.D(result_r_ns_0__15__N_3[437]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i438.GSR = "ENABLED";
    FD1P3AX result_r_31___i439 (.D(result_r_ns_0__15__N_3[438]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i439.GSR = "ENABLED";
    FD1P3AX result_r_31___i440 (.D(result_r_ns_0__15__N_3[439]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i440.GSR = "ENABLED";
    FD1P3AX result_r_31___i441 (.D(result_r_ns_0__15__N_3[440]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i441.GSR = "ENABLED";
    FD1P3AX result_r_31___i442 (.D(result_r_ns_0__15__N_3[441]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i442.GSR = "ENABLED";
    FD1P3AX result_r_31___i443 (.D(result_r_ns_0__15__N_3[442]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i443.GSR = "ENABLED";
    FD1P3AX result_r_31___i444 (.D(result_r_ns_0__15__N_3[443]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i444.GSR = "ENABLED";
    FD1P3AX result_r_31___i445 (.D(result_r_ns_0__15__N_3[444]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i445.GSR = "ENABLED";
    FD1P3AX result_r_31___i446 (.D(result_r_ns_0__15__N_3[445]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i446.GSR = "ENABLED";
    FD1P3AX result_r_31___i447 (.D(result_r_ns_0__15__N_3[446]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i447.GSR = "ENABLED";
    FD1P3AX result_r_31___i448 (.D(result_r_ns_0__15__N_3[447]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[4] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i448.GSR = "ENABLED";
    FD1P3AX result_r_31___i449 (.D(result_r_ns_0__15__N_3[448]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i449.GSR = "ENABLED";
    FD1P3AX result_r_31___i450 (.D(result_r_ns_0__15__N_3[449]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i450.GSR = "ENABLED";
    FD1P3AX result_r_31___i451 (.D(result_r_ns_0__15__N_3[450]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i451.GSR = "ENABLED";
    FD1P3AX result_r_31___i452 (.D(result_r_ns_0__15__N_3[451]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i452.GSR = "ENABLED";
    FD1P3AX result_r_31___i453 (.D(result_r_ns_0__15__N_3[452]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i453.GSR = "ENABLED";
    FD1P3AX result_r_31___i454 (.D(result_r_ns_0__15__N_3[453]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i454.GSR = "ENABLED";
    FD1P3AX result_r_31___i455 (.D(result_r_ns_0__15__N_3[454]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i455.GSR = "ENABLED";
    FD1P3AX result_r_31___i456 (.D(result_r_ns_0__15__N_3[455]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i456.GSR = "ENABLED";
    FD1P3AX result_r_31___i457 (.D(result_r_ns_0__15__N_3[456]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i457.GSR = "ENABLED";
    FD1P3AX result_r_31___i458 (.D(result_r_ns_0__15__N_3[457]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i458.GSR = "ENABLED";
    FD1P3AX result_r_31___i459 (.D(result_r_ns_0__15__N_3[458]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i459.GSR = "ENABLED";
    FD1P3AX result_r_31___i460 (.D(result_r_ns_0__15__N_3[459]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i460.GSR = "ENABLED";
    FD1P3AX result_r_31___i461 (.D(result_r_ns_0__15__N_3[460]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i461.GSR = "ENABLED";
    FD1P3AX result_r_31___i462 (.D(result_r_ns_0__15__N_3[461]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i462.GSR = "ENABLED";
    FD1P3AX result_r_31___i463 (.D(result_r_ns_0__15__N_3[462]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i463.GSR = "ENABLED";
    FD1P3AX result_r_31___i464 (.D(result_r_ns_0__15__N_3[463]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[3] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i464.GSR = "ENABLED";
    FD1P3AX result_r_31___i465 (.D(result_r_ns_0__15__N_3[464]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i465.GSR = "ENABLED";
    FD1P3AX result_r_31___i466 (.D(result_r_ns_0__15__N_3[465]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i466.GSR = "ENABLED";
    FD1P3AX result_r_31___i467 (.D(result_r_ns_0__15__N_3[466]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i467.GSR = "ENABLED";
    FD1P3AX result_r_31___i468 (.D(result_r_ns_0__15__N_3[467]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i468.GSR = "ENABLED";
    FD1P3AX result_r_31___i469 (.D(result_r_ns_0__15__N_3[468]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i469.GSR = "ENABLED";
    FD1P3AX result_r_31___i470 (.D(result_r_ns_0__15__N_3[469]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i470.GSR = "ENABLED";
    FD1P3AX result_r_31___i471 (.D(result_r_ns_0__15__N_3[470]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i471.GSR = "ENABLED";
    FD1P3AX result_r_31___i472 (.D(result_r_ns_0__15__N_3[471]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i472.GSR = "ENABLED";
    FD1P3AX result_r_31___i473 (.D(result_r_ns_0__15__N_3[472]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i473.GSR = "ENABLED";
    FD1P3AX result_r_31___i474 (.D(result_r_ns_0__15__N_3[473]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i474.GSR = "ENABLED";
    FD1P3AX result_r_31___i475 (.D(result_r_ns_0__15__N_3[474]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i475.GSR = "ENABLED";
    FD1P3AX result_r_31___i476 (.D(result_r_ns_0__15__N_3[475]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i476.GSR = "ENABLED";
    FD1P3AX result_r_31___i477 (.D(result_r_ns_0__15__N_3[476]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i477.GSR = "ENABLED";
    FD1P3AX result_r_31___i478 (.D(result_r_ns_0__15__N_3[477]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i478.GSR = "ENABLED";
    FD1P3AX result_r_31___i479 (.D(result_r_ns_0__15__N_3[478]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i479.GSR = "ENABLED";
    FD1P3AX result_r_31___i480 (.D(result_r_ns_0__15__N_3[479]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[2] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i480.GSR = "ENABLED";
    FD1P3AX result_r_31___i481 (.D(result_r_ns_0__15__N_3[480]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i481.GSR = "ENABLED";
    FD1P3AX result_r_31___i482 (.D(result_r_ns_0__15__N_3[481]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i482.GSR = "ENABLED";
    FD1P3AX result_r_31___i483 (.D(result_r_ns_0__15__N_3[482]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i483.GSR = "ENABLED";
    FD1P3AX result_r_31___i484 (.D(result_r_ns_0__15__N_3[483]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i484.GSR = "ENABLED";
    FD1P3AX result_r_31___i485 (.D(result_r_ns_0__15__N_3[484]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i485.GSR = "ENABLED";
    FD1P3AX result_r_31___i486 (.D(result_r_ns_0__15__N_3[485]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i486.GSR = "ENABLED";
    FD1P3AX result_r_31___i487 (.D(result_r_ns_0__15__N_3[486]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i487.GSR = "ENABLED";
    FD1P3AX result_r_31___i488 (.D(result_r_ns_0__15__N_3[487]), .SP(clk_c_enable_2259), 
            .CK(clk_c), .Q(\result_r[1] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i488.GSR = "ENABLED";
    FD1P3AX result_r_31___i489 (.D(result_r_ns_0__15__N_3[488]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i489.GSR = "ENABLED";
    FD1P3AX result_r_31___i490 (.D(result_r_ns_0__15__N_3[489]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i490.GSR = "ENABLED";
    FD1P3AX result_r_31___i491 (.D(result_r_ns_0__15__N_3[490]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i491.GSR = "ENABLED";
    FD1P3AX result_r_31___i492 (.D(result_r_ns_0__15__N_3[491]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i492.GSR = "ENABLED";
    FD1P3AX result_r_31___i493 (.D(result_r_ns_0__15__N_3[492]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i493.GSR = "ENABLED";
    FD1P3AX result_r_31___i494 (.D(result_r_ns_0__15__N_3[493]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i494.GSR = "ENABLED";
    FD1P3AX result_r_31___i495 (.D(result_r_ns_0__15__N_3[494]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i495.GSR = "ENABLED";
    FD1P3AX result_r_31___i496 (.D(result_r_ns_0__15__N_3[495]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[1] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i496.GSR = "ENABLED";
    FD1P3AX result_r_31___i497 (.D(result_r_ns_0__15__N_3[496]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i497.GSR = "ENABLED";
    FD1P3AX result_r_31___i498 (.D(result_r_ns_0__15__N_3[497]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i498.GSR = "ENABLED";
    FD1P3AX result_r_31___i499 (.D(result_r_ns_0__15__N_3[498]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i499.GSR = "ENABLED";
    FD1P3AX result_r_31___i500 (.D(result_r_ns_0__15__N_3[499]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i500.GSR = "ENABLED";
    FD1P3AX result_r_31___i501 (.D(result_r_ns_0__15__N_3[500]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i501.GSR = "ENABLED";
    FD1P3AX result_r_31___i502 (.D(result_r_ns_0__15__N_3[501]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i502.GSR = "ENABLED";
    FD1P3AX result_r_31___i503 (.D(result_r_ns_0__15__N_3[502]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [6]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i503.GSR = "ENABLED";
    FD1P3AX result_r_31___i504 (.D(result_r_ns_0__15__N_3[503]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [7]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i504.GSR = "ENABLED";
    FD1P3AX result_r_31___i505 (.D(result_r_ns_0__15__N_3[504]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [8]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i505.GSR = "ENABLED";
    FD1P3AX result_r_31___i506 (.D(result_r_ns_0__15__N_3[505]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [9]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i506.GSR = "ENABLED";
    FD1P3AX result_r_31___i507 (.D(result_r_ns_0__15__N_3[506]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [10]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i507.GSR = "ENABLED";
    FD1P3AX result_r_31___i508 (.D(result_r_ns_0__15__N_3[507]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [11]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i508.GSR = "ENABLED";
    FD1P3AX result_r_31___i509 (.D(result_r_ns_0__15__N_3[508]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [12]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i509.GSR = "ENABLED";
    FD1P3AX result_r_31___i510 (.D(result_r_ns_0__15__N_3[509]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [13]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i510.GSR = "ENABLED";
    FD1P3AX result_r_31___i511 (.D(result_r_ns_0__15__N_3[510]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [14]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i511.GSR = "ENABLED";
    FD1P3AX result_r_31___i512 (.D(result_r_ns_0__15__N_3[511]), .SP(clk_c_enable_2283), 
            .CK(clk_c), .Q(\result_r[0] [15]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam result_r_31___i512.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i2 (.D(next_dout_r_15__N_1029[1]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_1));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i2.GSR = "ENABLED";
    PFUMX i15546 (.BLUT(n33920), .ALUT(n33921), .C0(y_1_delay[1]), .Z(n33930));
    LUT4 i2534_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[505])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2534_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15599_3_lut (.A(\result_r[26] [9]), .B(\result_r[27] [9]), .C(y_1_delay[0]), 
         .Z(n33983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15599_3_lut.init = 16'hcaca;
    LUT4 i2526_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[506])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2526_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2518_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[507])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2518_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15432_3_lut (.A(\result_r[2] [14]), .B(\result_r[3] [14]), .C(y_1_delay[0]), 
         .Z(n33816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15432_3_lut.init = 16'hcaca;
    LUT4 i2510_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[508])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2510_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15297 (.BLUT(n33670), .ALUT(n33671), .C0(y_1_delay[1]), .Z(n33681));
    PFUMX i15204 (.BLUT(n33577), .ALUT(n33578), .C0(y_1_delay[1]), .Z(n33588));
    LUT4 i15598_3_lut (.A(\result_r[24] [9]), .B(\result_r[25] [9]), .C(y_1_delay[0]), 
         .Z(n33982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15598_3_lut.init = 16'hcaca;
    LUT4 i15091_3_lut (.A(\result_i[2] [10]), .B(\result_i[3] [10]), .C(y_1_delay[0]), 
         .Z(n33475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15091_3_lut.init = 16'hcaca;
    LUT4 i15090_3_lut (.A(\result_i[0] [10]), .B(\result_i[1] [10]), .C(y_1_delay[0]), 
         .Z(n33474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15090_3_lut.init = 16'hcaca;
    LUT4 i15010_3_lut (.A(\result_i[26] [13]), .B(\result_i[27] [13]), .C(y_1_delay[0]), 
         .Z(n33394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15010_3_lut.init = 16'hcaca;
    LUT4 i15009_3_lut (.A(\result_i[24] [13]), .B(\result_i[25] [13]), .C(y_1_delay[0]), 
         .Z(n33393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15009_3_lut.init = 16'hcaca;
    LUT4 i15413_3_lut (.A(\result_r[26] [15]), .B(\result_r[27] [15]), .C(y_1_delay[0]), 
         .Z(n33797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15413_3_lut.init = 16'hcaca;
    LUT4 i15412_3_lut (.A(\result_r[24] [15]), .B(\result_r[25] [15]), .C(y_1_delay[0]), 
         .Z(n33796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15412_3_lut.init = 16'hcaca;
    LUT4 i15723_3_lut (.A(\result_r[26] [5]), .B(\result_r[27] [5]), .C(y_1_delay[0]), 
         .Z(n34107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15723_3_lut.init = 16'hcaca;
    LUT4 i15722_3_lut (.A(\result_r[24] [5]), .B(\result_r[25] [5]), .C(y_1_delay[0]), 
         .Z(n34106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15722_3_lut.init = 16'hcaca;
    LUT4 i15411_3_lut (.A(\result_r[22] [15]), .B(\result_r[23] [15]), .C(y_1_delay[0]), 
         .Z(n33795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15411_3_lut.init = 16'hcaca;
    LUT4 i15410_3_lut (.A(\result_r[20] [15]), .B(\result_r[21] [15]), .C(y_1_delay[0]), 
         .Z(n33794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15410_3_lut.init = 16'hcaca;
    LUT4 i15008_3_lut (.A(\result_i[22] [13]), .B(\result_i[23] [13]), .C(y_1_delay[0]), 
         .Z(n33392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15008_3_lut.init = 16'hcaca;
    LUT4 i15007_3_lut (.A(\result_i[20] [13]), .B(\result_i[21] [13]), .C(y_1_delay[0]), 
         .Z(n33391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15007_3_lut.init = 16'hcaca;
    LUT4 i15721_3_lut (.A(\result_r[22] [5]), .B(\result_r[23] [5]), .C(y_1_delay[0]), 
         .Z(n34105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15721_3_lut.init = 16'hcaca;
    LUT4 i15720_3_lut (.A(\result_r[20] [5]), .B(\result_r[21] [5]), .C(y_1_delay[0]), 
         .Z(n34104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15720_3_lut.init = 16'hcaca;
    LUT4 i15409_3_lut (.A(\result_r[18] [15]), .B(\result_r[19] [15]), .C(y_1_delay[0]), 
         .Z(n33793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15409_3_lut.init = 16'hcaca;
    LUT4 i2502_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [13]), 
         .D(out_i[21]), .Z(result_i_ns_0__15__N_517[509])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2502_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15431_3_lut (.A(\result_r[0] [14]), .B(\result_r[1] [14]), .C(y_1_delay[0]), 
         .Z(n33815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15431_3_lut.init = 16'hcaca;
    LUT4 i2494_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [14]), 
         .D(out_i[22]), .Z(result_i_ns_0__15__N_517[510])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2494_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15408_3_lut (.A(\result_r[16] [15]), .B(\result_r[17] [15]), .C(y_1_delay[0]), 
         .Z(n33792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15408_3_lut.init = 16'hcaca;
    LUT4 i15407_3_lut (.A(\result_r[14] [15]), .B(\result_r[15] [15]), .C(y_1_delay[0]), 
         .Z(n33791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15407_3_lut.init = 16'hcaca;
    PFUMX i15205 (.BLUT(n33579), .ALUT(n33580), .C0(y_1_delay[1]), .Z(n33589));
    LUT4 i15406_3_lut (.A(\result_r[12] [15]), .B(\result_r[13] [15]), .C(y_1_delay[0]), 
         .Z(n33790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15406_3_lut.init = 16'hcaca;
    LUT4 i15006_3_lut (.A(\result_i[18] [13]), .B(\result_i[19] [13]), .C(y_1_delay[0]), 
         .Z(n33390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15006_3_lut.init = 16'hcaca;
    LUT4 i15005_3_lut (.A(\result_i[16] [13]), .B(\result_i[17] [13]), .C(y_1_delay[0]), 
         .Z(n33389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15005_3_lut.init = 16'hcaca;
    LUT4 i15103_3_lut (.A(\result_i[26] [10]), .B(\result_i[27] [10]), .C(y_1_delay[0]), 
         .Z(n33487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15103_3_lut.init = 16'hcaca;
    LUT4 i2486_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_i[0] [15]), 
         .D(out_i[23]), .Z(result_i_ns_0__15__N_517[511])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2486_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15547 (.BLUT(n33922), .ALUT(n33923), .C0(y_1_delay[1]), .Z(n33931));
    LUT4 i15229_3_lut (.A(\result_i[30] [6]), .B(\result_i[31] [6]), .C(y_1_delay[0]), 
         .Z(n33613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15229_3_lut.init = 16'hcaca;
    LUT4 i15405_3_lut (.A(\result_r[10] [15]), .B(\result_r[11] [15]), .C(y_1_delay[0]), 
         .Z(n33789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15405_3_lut.init = 16'hcaca;
    PFUMX i15206 (.BLUT(n33581), .ALUT(n33582), .C0(y_1_delay[1]), .Z(n33590));
    PFUMX i15298 (.BLUT(n33672), .ALUT(n33673), .C0(y_1_delay[1]), .Z(n33682));
    LUT4 i15012_3_lut (.A(\result_i[30] [13]), .B(\result_i[31] [13]), .C(y_1_delay[0]), 
         .Z(n33396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15012_3_lut.init = 16'hcaca;
    LUT4 i6697_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [0]), 
         .D(out_r[8]), .Z(result_r_ns_0__15__N_3[496])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6697_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15404_3_lut (.A(\result_r[8] [15]), .B(\result_r[9] [15]), .C(y_1_delay[0]), 
         .Z(n33788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15404_3_lut.init = 16'hcaca;
    LUT4 i6769_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[487])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6769_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15004_3_lut (.A(\result_i[14] [13]), .B(\result_i[15] [13]), .C(y_1_delay[0]), 
         .Z(n33388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15004_3_lut.init = 16'hcaca;
    LUT4 i15003_3_lut (.A(\result_i[12] [13]), .B(\result_i[13] [13]), .C(y_1_delay[0]), 
         .Z(n33387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15003_3_lut.init = 16'hcaca;
    LUT4 i15002_3_lut (.A(\result_i[10] [13]), .B(\result_i[11] [13]), .C(y_1_delay[0]), 
         .Z(n33386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15002_3_lut.init = 16'hcaca;
    LUT4 i15001_3_lut (.A(\result_i[8] [13]), .B(\result_i[9] [13]), .C(y_1_delay[0]), 
         .Z(n33385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15001_3_lut.init = 16'hcaca;
    LUT4 i15000_3_lut (.A(\result_i[6] [13]), .B(\result_i[7] [13]), .C(y_1_delay[0]), 
         .Z(n33384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15000_3_lut.init = 16'hcaca;
    LUT4 i14999_3_lut (.A(\result_i[4] [13]), .B(\result_i[5] [13]), .C(y_1_delay[0]), 
         .Z(n33383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14999_3_lut.init = 16'hcaca;
    LUT4 i6689_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [1]), 
         .D(out_r[9]), .Z(result_r_ns_0__15__N_3[497])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6689_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15719_3_lut (.A(\result_r[18] [5]), .B(\result_r[19] [5]), .C(y_1_delay[0]), 
         .Z(n34103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15719_3_lut.init = 16'hcaca;
    LUT4 i15718_3_lut (.A(\result_r[16] [5]), .B(\result_r[17] [5]), .C(y_1_delay[0]), 
         .Z(n34102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15718_3_lut.init = 16'hcaca;
    LUT4 i15102_3_lut (.A(\result_i[24] [10]), .B(\result_i[25] [10]), .C(y_1_delay[0]), 
         .Z(n33486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15102_3_lut.init = 16'hcaca;
    LUT4 i14998_3_lut (.A(\result_i[2] [13]), .B(\result_i[3] [13]), .C(y_1_delay[0]), 
         .Z(n33382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14998_3_lut.init = 16'hcaca;
    LUT4 i14997_3_lut (.A(\result_i[0] [13]), .B(\result_i[1] [13]), .C(y_1_delay[0]), 
         .Z(n33381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14997_3_lut.init = 16'hcaca;
    LUT4 i15011_3_lut (.A(\result_i[28] [13]), .B(\result_i[29] [13]), .C(y_1_delay[0]), 
         .Z(n33395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15011_3_lut.init = 16'hcaca;
    LUT4 i15403_3_lut (.A(\result_r[6] [15]), .B(\result_r[7] [15]), .C(y_1_delay[0]), 
         .Z(n33787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15403_3_lut.init = 16'hcaca;
    LUT4 i15402_3_lut (.A(\result_r[4] [15]), .B(\result_r[5] [15]), .C(y_1_delay[0]), 
         .Z(n33786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15402_3_lut.init = 16'hcaca;
    LUT4 i15401_3_lut (.A(\result_r[2] [15]), .B(\result_r[3] [15]), .C(y_1_delay[0]), 
         .Z(n33785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15401_3_lut.init = 16'hcaca;
    LUT4 i15400_3_lut (.A(\result_r[0] [15]), .B(\result_r[1] [15]), .C(y_1_delay[0]), 
         .Z(n33784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15400_3_lut.init = 16'hcaca;
    PFUMX i15850 (.BLUT(n34218), .ALUT(n34219), .C0(y_1_delay[1]), .Z(n34234));
    LUT4 i14950_3_lut (.A(\result_i[30] [15]), .B(\result_i[31] [15]), .C(y_1_delay[0]), 
         .Z(n33334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14950_3_lut.init = 16'hcaca;
    LUT4 i6681_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [2]), 
         .D(out_r[10]), .Z(result_r_ns_0__15__N_3[498])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6681_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14949_3_lut (.A(\result_i[28] [15]), .B(\result_i[29] [15]), .C(y_1_delay[0]), 
         .Z(n33333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14949_3_lut.init = 16'hcaca;
    LUT4 i6673_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [3]), 
         .D(out_r[11]), .Z(result_r_ns_0__15__N_3[499])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6673_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15136_3_lut (.A(\result_i[30] [9]), .B(\result_i[31] [9]), .C(y_1_delay[0]), 
         .Z(n33520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15136_3_lut.init = 16'hcaca;
    PFUMX i15851 (.BLUT(n34220), .ALUT(n34221), .C0(y_1_delay[1]), .Z(n34235));
    LUT4 i15101_3_lut (.A(\result_i[22] [10]), .B(\result_i[23] [10]), .C(y_1_delay[0]), 
         .Z(n33485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15101_3_lut.init = 16'hcaca;
    LUT4 i15414_3_lut (.A(\result_r[28] [15]), .B(\result_r[29] [15]), .C(y_1_delay[0]), 
         .Z(n33798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15414_3_lut.init = 16'hcaca;
    LUT4 i6665_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [4]), 
         .D(out_r[12]), .Z(result_r_ns_0__15__N_3[500])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6665_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i15852 (.BLUT(n34222), .ALUT(n34223), .C0(y_1_delay[1]), .Z(n34236));
    PFUMX i15853 (.BLUT(n34224), .ALUT(n34225), .C0(y_1_delay[1]), .Z(n34237));
    LUT4 i15100_3_lut (.A(\result_i[20] [10]), .B(\result_i[21] [10]), .C(y_1_delay[0]), 
         .Z(n33484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15100_3_lut.init = 16'hcaca;
    LUT4 i15228_3_lut (.A(\result_i[28] [6]), .B(\result_i[29] [6]), .C(y_1_delay[0]), 
         .Z(n33612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15228_3_lut.init = 16'hcaca;
    LUT4 i6657_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [5]), 
         .D(out_r[13]), .Z(result_r_ns_0__15__N_3[501])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6657_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15099_3_lut (.A(\result_i[18] [10]), .B(\result_i[19] [10]), .C(y_1_delay[0]), 
         .Z(n33483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15099_3_lut.init = 16'hcaca;
    VLO i1 (.Z(GND_net));
    PFUMX i15854 (.BLUT(n34226), .ALUT(n34227), .C0(y_1_delay[1]), .Z(n34238));
    PFUMX i15855 (.BLUT(n34228), .ALUT(n34229), .C0(y_1_delay[1]), .Z(n34239));
    LUT4 i6649_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [6]), 
         .D(out_r[14]), .Z(result_r_ns_0__15__N_3[502])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6649_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15098_3_lut (.A(\result_i[16] [10]), .B(\result_i[17] [10]), .C(y_1_delay[0]), 
         .Z(n33482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15098_3_lut.init = 16'hcaca;
    LUT4 i6641_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [7]), 
         .D(out_r[15]), .Z(result_r_ns_0__15__N_3[503])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6641_3_lut_4_lut.init = 16'hf1e0;
    shift_2 shift_2 (.shift_2_dout_r({shift_2_dout_r}), .clk_c(clk_c), .clk_c_enable_1396(clk_c_enable_1396), 
            .\dout_i_23__N_5777[0] (dout_i_23__N_5777[0]), .\dout_r_23__N_5681[0] (dout_r_23__N_5681[0]), 
            .valid(valid_adj_7001), .clk_c_enable_2299(clk_c_enable_2299), 
            .VCC_net(VCC_net), .\dout_i_23__N_5777[1] (dout_i_23__N_5777[1]), 
            .\dout_i_23__N_5777[2] (dout_i_23__N_5777[2]), .\dout_i_23__N_5777[3] (dout_i_23__N_5777[3]), 
            .\dout_i_23__N_5777[4] (dout_i_23__N_5777[4]), .\dout_i_23__N_5777[5] (dout_i_23__N_5777[5]), 
            .\dout_i_23__N_5777[6] (dout_i_23__N_5777[6]), .\dout_i_23__N_5777[7] (dout_i_23__N_5777[7]), 
            .\dout_i_23__N_5777[8] (dout_i_23__N_5777[8]), .\dout_i_23__N_5777[9] (dout_i_23__N_5777[9]), 
            .\dout_i_23__N_5777[10] (dout_i_23__N_5777[10]), .\dout_i_23__N_5777[11] (dout_i_23__N_5777[11]), 
            .\dout_i_23__N_5777[12] (dout_i_23__N_5777[12]), .\dout_i_23__N_5777[13] (dout_i_23__N_5777[13]), 
            .\dout_i_23__N_5777[14] (dout_i_23__N_5777[14]), .\dout_i_23__N_5777[15] (dout_i_23__N_5777[15]), 
            .\dout_i_23__N_5777[16] (dout_i_23__N_5777[16]), .\dout_i_23__N_5777[17] (dout_i_23__N_5777[17]), 
            .\dout_i_23__N_5777[18] (dout_i_23__N_5777[18]), .\dout_i_23__N_5777[19] (dout_i_23__N_5777[19]), 
            .\dout_i_23__N_5777[20] (dout_i_23__N_5777[20]), .\dout_i_23__N_5777[21] (dout_i_23__N_5777[21]), 
            .\dout_i_23__N_5777[22] (dout_i_23__N_5777[22]), .\dout_i_23__N_5777[23] (dout_i_23__N_5777[23]), 
            .\dout_r_23__N_5681[1] (dout_r_23__N_5681[1]), .\dout_r_23__N_5681[2] (dout_r_23__N_5681[2]), 
            .\dout_r_23__N_5681[3] (dout_r_23__N_5681[3]), .\dout_r_23__N_5681[4] (dout_r_23__N_5681[4]), 
            .\dout_r_23__N_5681[5] (dout_r_23__N_5681[5]), .\dout_r_23__N_5681[6] (dout_r_23__N_5681[6]), 
            .\dout_r_23__N_5681[7] (dout_r_23__N_5681[7]), .\dout_r_23__N_5681[8] (dout_r_23__N_5681[8]), 
            .\dout_r_23__N_5681[9] (dout_r_23__N_5681[9]), .\dout_r_23__N_5681[10] (dout_r_23__N_5681[10]), 
            .\dout_r_23__N_5681[11] (dout_r_23__N_5681[11]), .\dout_r_23__N_5681[12] (dout_r_23__N_5681[12]), 
            .\dout_r_23__N_5681[13] (dout_r_23__N_5681[13]), .\dout_r_23__N_5681[14] (dout_r_23__N_5681[14]), 
            .\dout_r_23__N_5681[15] (dout_r_23__N_5681[15]), .\dout_r_23__N_5681[16] (dout_r_23__N_5681[16]), 
            .\dout_r_23__N_5681[17] (dout_r_23__N_5681[17]), .\dout_r_23__N_5681[18] (dout_r_23__N_5681[18]), 
            .\dout_r_23__N_5681[19] (dout_r_23__N_5681[19]), .\dout_r_23__N_5681[20] (dout_r_23__N_5681[20]), 
            .\dout_r_23__N_5681[21] (dout_r_23__N_5681[21]), .\dout_r_23__N_5681[22] (dout_r_23__N_5681[22]), 
            .\dout_r_23__N_5681[23] (dout_r_23__N_5681[23]), .n34841(n34841), 
            .shift_2_dout_i({shift_2_dout_i})) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(198[9] 205[2])
    shift_4 shift_4 (.clk_c(clk_c), .clk_c_enable_1373(clk_c_enable_1373), 
            .\dout_r_23__N_5203[0] (dout_r_23__N_5203[0]), .\dout_i_23__N_5395[0] (dout_i_23__N_5395[0]), 
            .valid(valid_adj_6771), .clk_c_enable_2305(clk_c_enable_2305), 
            .VCC_net(VCC_net), .\dout_r_23__N_5203[1] (dout_r_23__N_5203[1]), 
            .\dout_r_23__N_5203[2] (dout_r_23__N_5203[2]), .\dout_r_23__N_5203[3] (dout_r_23__N_5203[3]), 
            .\dout_r_23__N_5203[4] (dout_r_23__N_5203[4]), .\dout_r_23__N_5203[5] (dout_r_23__N_5203[5]), 
            .\dout_r_23__N_5203[6] (dout_r_23__N_5203[6]), .\dout_r_23__N_5203[7] (dout_r_23__N_5203[7]), 
            .\dout_r_23__N_5203[8] (dout_r_23__N_5203[8]), .\dout_r_23__N_5203[9] (dout_r_23__N_5203[9]), 
            .\dout_r_23__N_5203[10] (dout_r_23__N_5203[10]), .\dout_r_23__N_5203[11] (dout_r_23__N_5203[11]), 
            .\dout_r_23__N_5203[12] (dout_r_23__N_5203[12]), .\dout_r_23__N_5203[13] (dout_r_23__N_5203[13]), 
            .\dout_r_23__N_5203[14] (dout_r_23__N_5203[14]), .\dout_r_23__N_5203[15] (dout_r_23__N_5203[15]), 
            .\dout_r_23__N_5203[16] (dout_r_23__N_5203[16]), .\dout_r_23__N_5203[17] (dout_r_23__N_5203[17]), 
            .\dout_r_23__N_5203[18] (dout_r_23__N_5203[18]), .\dout_r_23__N_5203[19] (dout_r_23__N_5203[19]), 
            .\dout_r_23__N_5203[20] (dout_r_23__N_5203[20]), .\dout_r_23__N_5203[21] (dout_r_23__N_5203[21]), 
            .\dout_r_23__N_5203[22] (dout_r_23__N_5203[22]), .\dout_r_23__N_5203[23] (dout_r_23__N_5203[23]), 
            .\dout_i_23__N_5395[1] (dout_i_23__N_5395[1]), .\dout_i_23__N_5395[2] (dout_i_23__N_5395[2]), 
            .\dout_i_23__N_5395[3] (dout_i_23__N_5395[3]), .\dout_i_23__N_5395[4] (dout_i_23__N_5395[4]), 
            .\dout_i_23__N_5395[5] (dout_i_23__N_5395[5]), .\dout_i_23__N_5395[6] (dout_i_23__N_5395[6]), 
            .\dout_i_23__N_5395[7] (dout_i_23__N_5395[7]), .\dout_i_23__N_5395[8] (dout_i_23__N_5395[8]), 
            .\dout_i_23__N_5395[9] (dout_i_23__N_5395[9]), .\dout_i_23__N_5395[10] (dout_i_23__N_5395[10]), 
            .\dout_i_23__N_5395[11] (dout_i_23__N_5395[11]), .\dout_i_23__N_5395[12] (dout_i_23__N_5395[12]), 
            .\dout_i_23__N_5395[13] (dout_i_23__N_5395[13]), .\dout_i_23__N_5395[14] (dout_i_23__N_5395[14]), 
            .\dout_i_23__N_5395[15] (dout_i_23__N_5395[15]), .\dout_i_23__N_5395[16] (dout_i_23__N_5395[16]), 
            .\dout_i_23__N_5395[17] (dout_i_23__N_5395[17]), .\dout_i_23__N_5395[18] (dout_i_23__N_5395[18]), 
            .\dout_i_23__N_5395[19] (dout_i_23__N_5395[19]), .\dout_i_23__N_5395[20] (dout_i_23__N_5395[20]), 
            .\dout_i_23__N_5395[21] (dout_i_23__N_5395[21]), .\dout_i_23__N_5395[22] (dout_i_23__N_5395[22]), 
            .\dout_i_23__N_5395[23] (dout_i_23__N_5395[23]), .n34842(n34842), 
            .shift_4_dout_r({shift_4_dout_r}), .shift_4_dout_i({shift_4_dout_i})) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(164[9] 171[2])
    ROM_8 rom8 (.n29816(n29816), .n29815(n29815), .n34532(n34532), .\rom8_state[0] (rom8_state[0]), 
          .s_count({s_count}), .clk_c(clk_c), .clk_c_enable_2285(clk_c_enable_2285), 
          .clk_c_enable_2310(clk_c_enable_2310), .n34726(n34726), .n34788(n34788), 
          .\rom8_w_i[12] (rom8_w_i[12]), .n29782(n29782), .n5(n5), .n29824(n29824), 
          .n29823(n29823), .n29822(n29822), .n34842(n34842), .n30191(n30191), 
          .GND_net(GND_net), .VCC_net(VCC_net), .n34762(n34762), .n34761(n34761), 
          .n34760(n34760), .\rom8_w_i[1] (rom8_w_i[1]), .n34785(n34785), 
          .n34734(n34734), .\rom8_w_i[4] (rom8_w_i[4]), .\rom8_w_i[3] (rom8_w_i[3]), 
          .n34787(n34787), .\rom8_w_i[0] (rom8_w_i[0]), .\rom8_w_i[6] (rom8_w_i[6]), 
          .n34742(n34742), .\rom8_w_i[2] (rom8_w_i[2]), .n6(n6_adj_7292), 
          .n34778(n34778), .\rom8_w_r[0] (rom8_w_r[0]), .\rom8_w_r[7] (rom8_w_r[7]), 
          .n34752(n34752), .n34753(n34753), .\rom8_w_r[4] (rom8_w_r[4]), 
          .\rom8_w_r[3] (rom8_w_r[3]), .\rom8_w_r[6] (rom8_w_r[6]), .n34779(n34779), 
          .\rom8_w_r[1] (rom8_w_r[1]), .n34754(n34754), .\rom8_w_r[8] (rom8_w_r[8]), 
          .\rom8_w_r[5] (rom8_w_r[5]), .\rom8_w_r[10] (rom8_w_r[10]), .n34794(n34794), 
          .n34755(n34755), .n34756(n34756), .clk_c_enable_2305(clk_c_enable_2305), 
          .n30040(n30040)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(139[7] 146[2])
    LUT4 i6633_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[504])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6633_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6625_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[505])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6625_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14948_3_lut (.A(\result_i[26] [15]), .B(\result_i[27] [15]), .C(y_1_delay[0]), 
         .Z(n33332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14948_3_lut.init = 16'hcaca;
    LUT4 i6617_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [10]), 
         .D(out_r[18]), .Z(result_r_ns_0__15__N_3[506])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6617_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6609_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [11]), 
         .D(out_r[19]), .Z(result_r_ns_0__15__N_3[507])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6609_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15717_3_lut (.A(\result_r[14] [5]), .B(\result_r[15] [5]), .C(y_1_delay[0]), 
         .Z(n34101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15717_3_lut.init = 16'hcaca;
    LUT4 i6601_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [12]), 
         .D(out_r[20]), .Z(result_r_ns_0__15__N_3[508])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6601_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6593_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [13]), 
         .D(out_r[21]), .Z(result_r_ns_0__15__N_3[509])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6593_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6585_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [14]), 
         .D(out_r[22]), .Z(result_r_ns_0__15__N_3[510])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6585_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6577_3_lut_4_lut (.A(n34741), .B(n34703), .C(\result_r[0] [15]), 
         .D(out_r[23]), .Z(result_r_ns_0__15__N_3[511])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6577_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15597_3_lut (.A(\result_r[22] [9]), .B(\result_r[23] [9]), .C(y_1_delay[0]), 
         .Z(n33981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15597_3_lut.init = 16'hcaca;
    LUT4 i2735_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [0]), 
         .D(out_i[8]), .Z(result_i_ns_0__15__N_517[480])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2735_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15596_3_lut (.A(\result_r[20] [9]), .B(\result_r[21] [9]), .C(y_1_delay[0]), 
         .Z(n33980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15596_3_lut.init = 16'hcaca;
    PFUMX i15144 (.BLUT(n33519), .ALUT(n33520), .C0(y_1_delay[1]), .Z(n33528));
    PFUMX i15856 (.BLUT(n34230), .ALUT(n34231), .C0(y_1_delay[1]), .Z(n34240));
    PFUMX i15571 (.BLUT(n33939), .ALUT(n33940), .C0(y_1_delay[1]), .Z(n33955));
    LUT4 i2727_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [1]), 
         .D(out_i[9]), .Z(result_i_ns_0__15__N_517[481])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2727_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15097_3_lut (.A(\result_i[14] [10]), .B(\result_i[15] [10]), .C(y_1_delay[0]), 
         .Z(n33481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15097_3_lut.init = 16'hcaca;
    LUT4 i2719_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [2]), 
         .D(out_i[10]), .Z(result_i_ns_0__15__N_517[482])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2719_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15591_3_lut (.A(\result_r[10] [9]), .B(\result_r[11] [9]), .C(y_1_delay[0]), 
         .Z(n33975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15591_3_lut.init = 16'hcaca;
    LUT4 i15096_3_lut (.A(\result_i[12] [10]), .B(\result_i[13] [10]), .C(y_1_delay[0]), 
         .Z(n33480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15096_3_lut.init = 16'hcaca;
    PFUMX i15299 (.BLUT(n33674), .ALUT(n33675), .C0(y_1_delay[1]), .Z(n33683));
    PFUMX i15572 (.BLUT(n33941), .ALUT(n33942), .C0(y_1_delay[1]), .Z(n33956));
    LUT4 i2711_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [3]), 
         .D(out_i[11]), .Z(result_i_ns_0__15__N_517[483])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2711_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2703_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [4]), 
         .D(out_i[12]), .Z(result_i_ns_0__15__N_517[484])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2703_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2695_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [5]), 
         .D(out_i[13]), .Z(result_i_ns_0__15__N_517[485])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2695_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2687_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [6]), 
         .D(out_i[14]), .Z(result_i_ns_0__15__N_517[486])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2687_3_lut_4_lut.init = 16'hf2d0;
    FD1P3AX dout_r_i0_i3 (.D(next_dout_r_15__N_1029[2]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_2));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i3.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i4 (.D(next_dout_r_15__N_1029[3]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_3));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i4.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i5 (.D(next_dout_r_15__N_1029[4]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_4));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i5.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i6 (.D(next_dout_r_15__N_1029[5]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_5));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i6.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i7 (.D(next_dout_r_15__N_1029[6]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_6));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i7.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i8 (.D(next_dout_r_15__N_1029[7]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_7));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i8.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i9 (.D(next_dout_r_15__N_1029[8]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_8));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i9.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i10 (.D(next_dout_r_15__N_1029[9]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_9));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i10.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i11 (.D(next_dout_r_15__N_1029[10]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_10));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i11.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i12 (.D(next_dout_r_15__N_1029[11]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_11));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i12.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i13 (.D(next_dout_r_15__N_1029[12]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_12));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i13.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i14 (.D(next_dout_r_15__N_1029[13]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_13));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i14.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i15 (.D(next_dout_r_15__N_1029[14]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_14));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i15.GSR = "ENABLED";
    FD1P3AX dout_r_i0_i16 (.D(next_dout_r_15__N_1029[15]), .SP(next_out_valid), 
            .CK(clk_c), .Q(dout_r_c_15));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(282[10] 298[8])
    defparam dout_r_i0_i16.GSR = "ENABLED";
    LUT4 i2679_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [7]), 
         .D(out_i[15]), .Z(result_i_ns_0__15__N_517[487])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2679_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15857 (.BLUT(n34232), .ALUT(n34233), .C0(y_1_delay[1]), .Z(n34241));
    LUT4 i2671_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [8]), 
         .D(out_i[16]), .Z(result_i_ns_0__15__N_517[488])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2671_3_lut_4_lut.init = 16'hf2d0;
    radix2_U3 radix_no1 (.op_r_23__N_1106({op_r_23__N_1106}), .\count[5] (count[5]), 
            .\count[4] (count[4]), .\op_r_23__N_1082[8] (op_r_23__N_1082[8]), 
            .\radix_no1_op_r[0] (radix_no1_op_r[0]), .\op_r_23__N_1082[9] (op_r_23__N_1082[9]), 
            .\radix_no1_op_r[1] (radix_no1_op_r[1]), .GND_net(GND_net), 
            .\op_r_23__N_1268[0] (op_r_23__N_1268[0]), .\op_r_23__N_1268[1] (op_r_23__N_1268[1]), 
            .\op_r_23__N_1268[2] (op_r_23__N_1268[2]), .\op_r_23__N_1268[3] (op_r_23__N_1268[3]), 
            .\op_r_23__N_1268[4] (op_r_23__N_1268[4]), .\op_r_23__N_1268[5] (op_r_23__N_1268[5]), 
            .\op_r_23__N_1268[6] (op_r_23__N_1268[6]), .\op_r_23__N_1268[7] (op_r_23__N_1268[7]), 
            .\op_r_23__N_1268[8] (op_r_23__N_1268[8]), .\op_r_23__N_1268[9] (op_r_23__N_1268[9]), 
            .\op_r_23__N_1268[10] (op_r_23__N_1268[10]), .\op_r_23__N_1268[11] (op_r_23__N_1268[11]), 
            .\op_r_23__N_1268[12] (op_r_23__N_1268[12]), .\op_r_23__N_1268[13] (op_r_23__N_1268[13]), 
            .\op_r_23__N_1268[14] (op_r_23__N_1268[14]), .\op_r_23__N_1268[15] (op_r_23__N_1268[15]), 
            .\op_r_23__N_1268[16] (op_r_23__N_1268[16]), .\op_r_23__N_1268[17] (op_r_23__N_1268[17]), 
            .VCC_net(VCC_net), .\op_r_23__N_1082[10] (op_r_23__N_1082[10]), 
            .\radix_no1_op_r[2] (radix_no1_op_r[2]), .\op_r_23__N_1082[11] (op_r_23__N_1082[11]), 
            .\radix_no1_op_r[3] (radix_no1_op_r[3]), .\op_r_23__N_1082[12] (op_r_23__N_1082[12]), 
            .\radix_no1_op_r[4] (radix_no1_op_r[4]), .\op_i_23__N_1310[0] (op_i_23__N_1310[0]), 
            .\op_i_23__N_1310[1] (op_i_23__N_1310[1]), .\op_i_23__N_1310[2] (op_i_23__N_1310[2]), 
            .\op_i_23__N_1310[3] (op_i_23__N_1310[3]), .\op_i_23__N_1310[4] (op_i_23__N_1310[4]), 
            .\op_i_23__N_1310[5] (op_i_23__N_1310[5]), .n89(n89_adj_7164), 
            .n88(n88_adj_7165), .n87(n87_adj_7166), .n86(n86_adj_7216), 
            .n85(n85_adj_7217), .n84(n84_adj_7218), .n83(n83_adj_7219), 
            .n82(n82_adj_7220), .n81(n81_adj_7221), .n80(n80_adj_7222), 
            .n79(n79_adj_7223), .n78(n78_adj_7224), .n77(n77_adj_7225), 
            .n76(n76_adj_7226), .n75(n75_adj_7227), .n74(n74_adj_7228), 
            .n73(n73_adj_7229), .n72(n72_adj_7230), .n71(n71_adj_7231), 
            .n70(n70_adj_7232), .n69(n69_adj_7233), .n68(n68_adj_7234), 
            .n67(n67_adj_7235), .n66(n66_adj_7236), .n65(n65_adj_7237), 
            .\rom16_w_i[8] (rom16_w_i[8]), .n9983(n9983), .n9984(n9984), 
            .n9985(n9985), .n9986(n9986), .n9987(n9987), .n9988(n9988), 
            .\rom16_w_i[0] (rom16_w_i[0]), .\rom16_w_i[1] (rom16_w_i[1]), 
            .\rom16_w_i[2] (rom16_w_i[2]), .\rom16_w_i[3] (rom16_w_i[3]), 
            .\rom16_w_i[4] (rom16_w_i[4]), .\rom16_w_i[5] (rom16_w_i[5]), 
            .\rom16_w_i[6] (rom16_w_i[6]), .\rom16_w_i[7] (rom16_w_i[7]), 
            .\op_r_23__N_1082[13] (op_r_23__N_1082[13]), .\radix_no1_op_r[5] (radix_no1_op_r[5]), 
            .\op_r_23__N_1226[0] (op_r_23__N_1226[0]), .\op_r_23__N_1226[1] (op_r_23__N_1226[1]), 
            .\op_r_23__N_1226[2] (op_r_23__N_1226[2]), .\op_r_23__N_1226[3] (op_r_23__N_1226[3]), 
            .\op_r_23__N_1226[4] (op_r_23__N_1226[4]), .\op_r_23__N_1226[5] (op_r_23__N_1226[5]), 
            .\op_r_23__N_1226[6] (op_r_23__N_1226[6]), .\op_r_23__N_1226[7] (op_r_23__N_1226[7]), 
            .\op_r_23__N_1226[8] (op_r_23__N_1226[8]), .\op_r_23__N_1226[9] (op_r_23__N_1226[9]), 
            .\op_r_23__N_1226[10] (op_r_23__N_1226[10]), .\op_r_23__N_1226[11] (op_r_23__N_1226[11]), 
            .\op_r_23__N_1226[12] (op_r_23__N_1226[12]), .\op_r_23__N_1226[13] (op_r_23__N_1226[13]), 
            .\op_r_23__N_1226[14] (op_r_23__N_1226[14]), .\op_r_23__N_1226[15] (op_r_23__N_1226[15]), 
            .\op_r_23__N_1226[16] (op_r_23__N_1226[16]), .\op_r_23__N_1226[17] (op_r_23__N_1226[17]), 
            .\op_r_23__N_1226[18] (op_r_23__N_1226[18]), .\op_r_23__N_1226[19] (op_r_23__N_1226[19]), 
            .\op_r_23__N_1226[20] (op_r_23__N_1226[20]), .\op_r_23__N_1226[21] (op_r_23__N_1226[21]), 
            .\op_r_23__N_1226[22] (op_r_23__N_1226[22]), .\op_r_23__N_1226[23] (op_r_23__N_1226[23]), 
            .\op_r_23__N_1226[24] (op_r_23__N_1226[24]), .\op_r_23__N_1226[25] (op_r_23__N_1226[25]), 
            .\op_r_23__N_1226[26] (op_r_23__N_1226[26]), .\op_r_23__N_1226[27] (op_r_23__N_1226[27]), 
            .\op_r_23__N_1226[28] (op_r_23__N_1226[28]), .\op_r_23__N_1226[29] (op_r_23__N_1226[29]), 
            .\op_r_23__N_1226[30] (op_r_23__N_1226[30]), .\op_r_23__N_1226[31] (op_r_23__N_1226[31]), 
            .\op_r_23__N_1082[14] (op_r_23__N_1082[14]), .\radix_no1_op_r[6] (radix_no1_op_r[6]), 
            .\op_r_23__N_1268[18] (op_r_23__N_1268[18]), .\op_r_23__N_1268[19] (op_r_23__N_1268[19]), 
            .\op_r_23__N_1268[20] (op_r_23__N_1268[20]), .\op_r_23__N_1268[21] (op_r_23__N_1268[21]), 
            .\op_r_23__N_1268[22] (op_r_23__N_1268[22]), .\op_r_23__N_1268[23] (op_r_23__N_1268[23]), 
            .\op_r_23__N_1268[24] (op_r_23__N_1268[24]), .\op_r_23__N_1268[25] (op_r_23__N_1268[25]), 
            .\op_r_23__N_1268[26] (op_r_23__N_1268[26]), .\op_r_23__N_1268[27] (op_r_23__N_1268[27]), 
            .\op_r_23__N_1268[28] (op_r_23__N_1268[28]), .\op_r_23__N_1268[29] (op_r_23__N_1268[29]), 
            .\op_r_23__N_1268[30] (op_r_23__N_1268[30]), .\op_r_23__N_1268[31] (op_r_23__N_1268[31]), 
            .\rom16_w_r[9] (rom16_w_r[9]), .n12332(n12332), .n12333(n12333), 
            .n12334(n12334), .n12335(n12335), .n12336(n12336), .n12337(n12337), 
            .n12338(n12338), .\rom16_w_r[0] (rom16_w_r[0]), .\rom16_w_r[1] (rom16_w_r[1]), 
            .\rom16_w_r[2] (rom16_w_r[2]), .\rom16_w_r[3] (rom16_w_r[3]), 
            .\rom16_w_r[4] (rom16_w_r[4]), .\rom16_w_r[5] (rom16_w_r[5]), 
            .\rom16_w_r[6] (rom16_w_r[6]), .\rom16_w_r[7] (rom16_w_r[7]), 
            .\rom16_w_r[8] (rom16_w_r[8]), .n12314(n12314), .n12315(n12315), 
            .n12316(n12316), .n12317(n12317), .n12318(n12318), .n12319(n12319), 
            .n12320(n12320), .n12321(n12321), .n12322(n12322), .n12323(n12323), 
            .n12324(n12324), .n12325(n12325), .n12326(n12326), .n12327(n12327), 
            .n12328(n12328), .n12329(n12329), .n12330(n12330), .n12331(n12331), 
            .\op_r_23__N_1082[15] (op_r_23__N_1082[15]), .\radix_no1_op_r[7] (radix_no1_op_r[7]), 
            .op_i_23__N_1154({op_i_23__N_1154}), .\op_i_23__N_1130[8] (op_i_23__N_1130[8]), 
            .\radix_no1_op_i[0] (radix_no1_op_i[0]), .\op_i_23__N_1130[9] (op_i_23__N_1130[9]), 
            .\radix_no1_op_i[1] (radix_no1_op_i[1]), .\op_i_23__N_1130[10] (op_i_23__N_1130[10]), 
            .\radix_no1_op_i[2] (radix_no1_op_i[2]), .\op_i_23__N_1130[11] (op_i_23__N_1130[11]), 
            .\radix_no1_op_i[3] (radix_no1_op_i[3]), .\op_i_23__N_1130[12] (op_i_23__N_1130[12]), 
            .\radix_no1_op_i[4] (radix_no1_op_i[4]), .\op_i_23__N_1130[13] (op_i_23__N_1130[13]), 
            .\radix_no1_op_i[5] (radix_no1_op_i[5]), .\op_i_23__N_1130[14] (op_i_23__N_1130[14]), 
            .\radix_no1_op_i[6] (radix_no1_op_i[6]), .\op_i_23__N_1130[15] (op_i_23__N_1130[15]), 
            .\radix_no1_op_i[7] (radix_no1_op_i[7]), .n8593(n8593), .n8592(n8592), 
            .n8591(n8591), .n8590(n8590), .n8589(n8589), .n8588(n8588), 
            .n8587(n8587), .n8586(n8586), .n8585(n8585), .n8584(n8584), 
            .n8583(n8583), .n8582(n8582), .n8581(n8581), .n8580(n8580), 
            .n8579(n8579), .n8578(n8578), .n8577(n8577), .n8576(n8576), 
            .n8575(n8575), .n8574(n8574), .n8573(n8573), .n8572(n8572), 
            .n8571(n8571), .n8570(n8570), .n8569(n8569), .n8568(n8568), 
            .n319(n319), .n9989(n9989), .n9990(n9990), .n9991(n9991), 
            .n9992(n9992), .n9993(n9993), .n9994(n9994), .n9995(n9995), 
            .n9996(n9996), .n9997(n9997), .n9998(n9998), .n9999(n9999), 
            .n10000(n10000), .n10001(n10001), .n10002(n10002), .n10003(n10003), 
            .n10004(n10004), .n10005(n10005), .n10006(n10006), .\shift_16_dout_i[8] (shift_16_dout_i[8]), 
            .\shift_16_dout_i[9] (shift_16_dout_i[9]), .\shift_16_dout_i[10] (shift_16_dout_i[10]), 
            .\shift_16_dout_i[11] (shift_16_dout_i[11]), .\shift_16_dout_i[12] (shift_16_dout_i[12]), 
            .\shift_16_dout_i[13] (shift_16_dout_i[13]), .\shift_16_dout_i[14] (shift_16_dout_i[14]), 
            .\shift_16_dout_i[15] (shift_16_dout_i[15]), .\shift_16_dout_i[16] (shift_16_dout_i[16]), 
            .\shift_16_dout_i[17] (shift_16_dout_i[17]), .n12344(n12344), 
            .n12345(n12345), .n12346(n12346), .n12347(n12347), .n12348(n12348), 
            .n12349(n12349), .n12350(n12350), .n12351(n12351), .n12352(n12352), 
            .n12353(n12353), .n12368(n12368), .\shift_16_dout_i[18] (shift_16_dout_i[18]), 
            .\shift_16_dout_i[19] (shift_16_dout_i[19]), .\shift_16_dout_i[20] (shift_16_dout_i[20]), 
            .\shift_16_dout_i[21] (shift_16_dout_i[21]), .\shift_16_dout_i[22] (shift_16_dout_i[22]), 
            .\shift_16_dout_i[23] (shift_16_dout_i[23]), .clk_c_enable_2310(clk_c_enable_2310), 
            .n34755(n34755), .\shift_8_dout_r[22] (shift_8_dout_r[22]), 
            .n7539(n7539), .n34756(n34756), .\op_r_23__N_1082[30] (op_r_23__N_1082_adj_7327[30]), 
            .n31574(n31574), .\shift_8_dout_r[23] (shift_8_dout_r[23]), 
            .n7538(n7538), .\op_r_23__N_1082[31] (op_r_23__N_1082_adj_7327[31]), 
            .n31572(n31572), .\shift_8_dout_i[22] (shift_8_dout_i[22]), 
            .n7486(n7486), .\op_i_23__N_1130[30] (op_i_23__N_1130_adj_7330[30]), 
            .n31378(n31378), .\shift_8_dout_i[23] (shift_8_dout_i[23]), 
            .n7485(n7485), .\op_i_23__N_1130[31] (op_i_23__N_1130_adj_7330[31]), 
            .n31376(n31376), .\shift_8_dout_r[20] (shift_8_dout_r[20]), 
            .n7541(n7541), .\op_r_23__N_1082[28] (op_r_23__N_1082_adj_7327[28]), 
            .n31578(n31578), .\shift_8_dout_r[21] (shift_8_dout_r[21]), 
            .n7540(n7540), .\op_r_23__N_1082[29] (op_r_23__N_1082_adj_7327[29]), 
            .n31576(n31576), .\shift_8_dout_i[20] (shift_8_dout_i[20]), 
            .n7488(n7488), .\op_i_23__N_1130[28] (op_i_23__N_1130_adj_7330[28]), 
            .n31382(n31382), .\shift_8_dout_i[21] (shift_8_dout_i[21]), 
            .n7487(n7487), .\op_i_23__N_1130[29] (op_i_23__N_1130_adj_7330[29]), 
            .n31380(n31380), .\shift_8_dout_r[18] (shift_8_dout_r[18]), 
            .n7543(n7543), .\op_r_23__N_1082[26] (op_r_23__N_1082_adj_7327[26]), 
            .n31582(n31582), .\shift_8_dout_r[19] (shift_8_dout_r[19]), 
            .n7542(n7542), .\op_r_23__N_1082[27] (op_r_23__N_1082_adj_7327[27]), 
            .n31580(n31580), .\shift_8_dout_i[18] (shift_8_dout_i[18]), 
            .n7490(n7490), .\op_i_23__N_1130[26] (op_i_23__N_1130_adj_7330[26]), 
            .n31386(n31386), .\shift_8_dout_i[19] (shift_8_dout_i[19]), 
            .n7489(n7489), .\op_i_23__N_1130[27] (op_i_23__N_1130_adj_7330[27]), 
            .n31384(n31384), .\shift_8_dout_r[16] (shift_8_dout_r[16]), 
            .n7545(n7545), .\op_r_23__N_1082[24] (op_r_23__N_1082_adj_7327[24]), 
            .n31586(n31586), .\shift_8_dout_r[17] (shift_8_dout_r[17]), 
            .n7544(n7544), .\op_r_23__N_1082[25] (op_r_23__N_1082_adj_7327[25]), 
            .n31584(n31584), .\shift_8_dout_i[16] (shift_8_dout_i[16]), 
            .n7492(n7492), .\op_i_23__N_1130[24] (op_i_23__N_1130_adj_7330[24]), 
            .n31390(n31390), .\shift_8_dout_i[17] (shift_8_dout_i[17]), 
            .n7491(n7491), .\op_i_23__N_1130[25] (op_i_23__N_1130_adj_7330[25]), 
            .n31388(n31388), .\shift_8_dout_r[14] (shift_8_dout_r[14]), 
            .n7547(n7547), .\op_r_23__N_1082[22] (op_r_23__N_1082_adj_7327[22]), 
            .n31590(n31590), .\shift_8_dout_r[15] (shift_8_dout_r[15]), 
            .n7546(n7546), .\op_r_23__N_1082[23] (op_r_23__N_1082_adj_7327[23]), 
            .n31588(n31588), .\shift_8_dout_i[14] (shift_8_dout_i[14]), 
            .n7494(n7494), .\op_i_23__N_1130[22] (op_i_23__N_1130_adj_7330[22]), 
            .n31394(n31394), .\shift_8_dout_i[15] (shift_8_dout_i[15]), 
            .n7493(n7493), .\op_i_23__N_1130[23] (op_i_23__N_1130_adj_7330[23]), 
            .n31392(n31392), .\shift_8_dout_r[12] (shift_8_dout_r[12]), 
            .n7549(n7549), .\op_r_23__N_1082[20] (op_r_23__N_1082_adj_7327[20]), 
            .n31594(n31594), .\shift_8_dout_r[13] (shift_8_dout_r[13]), 
            .n7548(n7548), .\op_r_23__N_1082[21] (op_r_23__N_1082_adj_7327[21]), 
            .n31592(n31592), .\shift_8_dout_i[12] (shift_8_dout_i[12]), 
            .n7496(n7496), .\op_i_23__N_1130[20] (op_i_23__N_1130_adj_7330[20]), 
            .n31398(n31398), .\shift_8_dout_i[13] (shift_8_dout_i[13]), 
            .n7495(n7495), .\op_i_23__N_1130[21] (op_i_23__N_1130_adj_7330[21]), 
            .n31396(n31396), .\shift_8_dout_r[10] (shift_8_dout_r[10]), 
            .n7551(n7551), .\op_r_23__N_1082[18] (op_r_23__N_1082_adj_7327[18]), 
            .n31598(n31598), .\shift_8_dout_r[11] (shift_8_dout_r[11]), 
            .n7550(n7550), .\op_r_23__N_1082[19] (op_r_23__N_1082_adj_7327[19]), 
            .n31596(n31596), .\shift_8_dout_i[10] (shift_8_dout_i[10]), 
            .n7498(n7498), .\op_i_23__N_1130[18] (op_i_23__N_1130_adj_7330[18]), 
            .n31402(n31402), .\shift_8_dout_i[11] (shift_8_dout_i[11]), 
            .n7497(n7497), .\op_i_23__N_1130[19] (op_i_23__N_1130_adj_7330[19]), 
            .n31400(n31400), .\shift_8_dout_r[8] (shift_8_dout_r[8]), .n7553(n7553), 
            .\op_r_23__N_1082[16] (op_r_23__N_1082_adj_7327[16]), .n31602(n31602), 
            .\shift_8_dout_r[9] (shift_8_dout_r[9]), .n7552(n7552), .\op_r_23__N_1082[17] (op_r_23__N_1082_adj_7327[17]), 
            .n31600(n31600), .\shift_8_dout_i[8] (shift_8_dout_i[8]), .n7500(n7500), 
            .\op_i_23__N_1130[16] (op_i_23__N_1130_adj_7330[16]), .n31406(n31406), 
            .\shift_8_dout_i[9] (shift_8_dout_i[9]), .n7499(n7499), .\op_i_23__N_1130[17] (op_i_23__N_1130_adj_7330[17]), 
            .n31404(n31404), .\din_r_reg[8] (din_r_reg[8]), .\delay_r_23__N_1178[8] (delay_r_23__N_1178[8]), 
            .\dout_r_23__N_2506[8] (dout_r_23__N_2506[8]), .\din_r_reg[9] (din_r_reg[9]), 
            .\delay_r_23__N_1178[9] (delay_r_23__N_1178[9]), .\dout_r_23__N_2506[9] (dout_r_23__N_2506[9]), 
            .\din_r_reg[10] (din_r_reg[10]), .\delay_r_23__N_1178[10] (delay_r_23__N_1178[10]), 
            .\dout_r_23__N_2506[10] (dout_r_23__N_2506[10]), .\din_r_reg[11] (din_r_reg[11]), 
            .\delay_r_23__N_1178[11] (delay_r_23__N_1178[11]), .\dout_r_23__N_2506[11] (dout_r_23__N_2506[11]), 
            .\din_r_reg[12] (din_r_reg[12]), .\delay_r_23__N_1178[12] (delay_r_23__N_1178[12]), 
            .\dout_r_23__N_2506[12] (dout_r_23__N_2506[12]), .\din_r_reg[13] (din_r_reg[13]), 
            .\delay_r_23__N_1178[13] (delay_r_23__N_1178[13]), .\dout_r_23__N_2506[13] (dout_r_23__N_2506[13]), 
            .\din_r_reg[14] (din_r_reg[14]), .\delay_r_23__N_1178[14] (delay_r_23__N_1178[14]), 
            .\dout_r_23__N_2506[14] (dout_r_23__N_2506[14]), .\din_r_reg[15] (din_r_reg[15]), 
            .\delay_r_23__N_1178[15] (delay_r_23__N_1178[15]), .\dout_r_23__N_2506[15] (dout_r_23__N_2506[15]), 
            .\din_r_reg[16] (din_r_reg[16]), .\delay_r_23__N_1178[16] (delay_r_23__N_1178[16]), 
            .\dout_r_23__N_2506[16] (dout_r_23__N_2506[16]), .\din_r_reg[17] (din_r_reg[17]), 
            .\delay_r_23__N_1178[17] (delay_r_23__N_1178[17]), .\dout_r_23__N_2506[17] (dout_r_23__N_2506[17]), 
            .\din_r_reg[18] (din_r_reg[18]), .\delay_r_23__N_1178[18] (delay_r_23__N_1178[18]), 
            .\dout_r_23__N_2506[18] (dout_r_23__N_2506[18]), .\din_r_reg[23] (din_r_reg[23]), 
            .\delay_r_23__N_1178[19] (delay_r_23__N_1178[19]), .\dout_r_23__N_2506[19] (dout_r_23__N_2506[19]), 
            .\delay_r_23__N_1178[20] (delay_r_23__N_1178[20]), .\dout_r_23__N_2506[20] (dout_r_23__N_2506[20]), 
            .\delay_r_23__N_1178[21] (delay_r_23__N_1178[21]), .\dout_r_23__N_2506[21] (dout_r_23__N_2506[21]), 
            .\delay_r_23__N_1178[22] (delay_r_23__N_1178[22]), .\dout_r_23__N_2506[22] (dout_r_23__N_2506[22]), 
            .\delay_r_23__N_1178[23] (delay_r_23__N_1178[23]), .\dout_r_23__N_2506[23] (dout_r_23__N_2506[23]), 
            .\din_i_reg[8] (din_i_reg[8]), .\delay_i_23__N_1202[8] (delay_i_23__N_1202[8]), 
            .\dout_i_23__N_3274[8] (dout_i_23__N_3274[8]), .\din_i_reg[9] (din_i_reg[9]), 
            .\delay_i_23__N_1202[9] (delay_i_23__N_1202[9]), .\dout_i_23__N_3274[9] (dout_i_23__N_3274[9]), 
            .\din_i_reg[10] (din_i_reg[10]), .\delay_i_23__N_1202[10] (delay_i_23__N_1202[10]), 
            .\dout_i_23__N_3274[10] (dout_i_23__N_3274[10]), .\din_i_reg[11] (din_i_reg[11]), 
            .\delay_i_23__N_1202[11] (delay_i_23__N_1202[11]), .\dout_i_23__N_3274[11] (dout_i_23__N_3274[11]), 
            .\din_i_reg[12] (din_i_reg[12]), .\delay_i_23__N_1202[12] (delay_i_23__N_1202[12]), 
            .\dout_i_23__N_3274[12] (dout_i_23__N_3274[12]), .\din_i_reg[13] (din_i_reg[13]), 
            .\delay_i_23__N_1202[13] (delay_i_23__N_1202[13]), .\dout_i_23__N_3274[13] (dout_i_23__N_3274[13]), 
            .\din_i_reg[14] (din_i_reg[14]), .\delay_i_23__N_1202[14] (delay_i_23__N_1202[14]), 
            .\dout_i_23__N_3274[14] (dout_i_23__N_3274[14]), .\din_i_reg[15] (din_i_reg[15]), 
            .\delay_i_23__N_1202[15] (delay_i_23__N_1202[15]), .\dout_i_23__N_3274[15] (dout_i_23__N_3274[15]), 
            .\din_i_reg[16] (din_i_reg[16]), .\delay_i_23__N_1202[16] (delay_i_23__N_1202[16]), 
            .\dout_i_23__N_3274[16] (dout_i_23__N_3274[16]), .\din_i_reg[17] (din_i_reg[17]), 
            .\delay_i_23__N_1202[17] (delay_i_23__N_1202[17]), .\dout_i_23__N_3274[17] (dout_i_23__N_3274[17]), 
            .\din_i_reg[18] (din_i_reg[18]), .\delay_i_23__N_1202[18] (delay_i_23__N_1202[18]), 
            .\dout_i_23__N_3274[18] (dout_i_23__N_3274[18]), .\din_i_reg[23] (din_i_reg[23]), 
            .\delay_i_23__N_1202[19] (delay_i_23__N_1202[19]), .\dout_i_23__N_3274[19] (dout_i_23__N_3274[19]), 
            .\delay_i_23__N_1202[20] (delay_i_23__N_1202[20]), .\dout_i_23__N_3274[20] (dout_i_23__N_3274[20]), 
            .\delay_i_23__N_1202[21] (delay_i_23__N_1202[21]), .\dout_i_23__N_3274[21] (dout_i_23__N_3274[21]), 
            .\delay_i_23__N_1202[22] (delay_i_23__N_1202[22]), .\dout_i_23__N_3274[22] (dout_i_23__N_3274[22]), 
            .\delay_i_23__N_1202[23] (delay_i_23__N_1202[23]), .\dout_i_23__N_3274[23] (dout_i_23__N_3274[23]), 
            .n34659(n34659), .n34652(n34652), .n34651(n34651), .n34650(n34650), 
            .n34649(n34649), .n34642(n34642), .n34641(n34641), .n34640(n34640), 
            .n34639(n34639), .n34630(n34630), .n34629(n34629), .n34628(n34628), 
            .n34627(n34627), .n34618(n34618), .n34617(n34617), .n34616(n34616), 
            .n34615(n34615), .n34660(n34660), .n34661(n34661), .n34662(n34662), 
            .n34669(n34669), .n34670(n34670), .n34671(n34671), .n34672(n34672), 
            .n34675(n34675), .n34676(n34676), .n34677(n34677), .n34678(n34678), 
            .n34683(n34683), .n34684(n34684), .n34685(n34685), .n34686(n34686), 
            .valid(valid), .clk_c_enable_1419(clk_c_enable_1419)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(82[8] 95[2])
    PFUMX i15573 (.BLUT(n33943), .ALUT(n33944), .C0(y_1_delay[1]), .Z(n33957));
    LUT4 i15095_3_lut (.A(\result_i[10] [10]), .B(\result_i[11] [10]), .C(y_1_delay[0]), 
         .Z(n33479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15095_3_lut.init = 16'hcaca;
    LUT4 i2663_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [9]), 
         .D(out_i[17]), .Z(result_i_ns_0__15__N_517[489])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2663_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15574 (.BLUT(n33945), .ALUT(n33946), .C0(y_1_delay[1]), .Z(n33958));
    radix2_U0 radix_no4 (.\op_r_23__N_1106[14] (op_r_23__N_1106_adj_7370[14]), 
            .n34841(n34841), .n30179(n30179), .\delay_r_23__N_1178[14] (delay_r_23__N_1178_adj_7427[14]), 
            .\dout_r_23__N_5681[14] (dout_r_23__N_5681[14]), .\op_i_23__N_1154[13] (op_i_23__N_1154_adj_7371[13]), 
            .\delay_i_23__N_1202[13] (delay_i_23__N_1202_adj_7428[13]), .\dout_i_23__N_5777[13] (dout_i_23__N_5777[13]), 
            .\op_r_23__N_1106[21] (op_r_23__N_1106_adj_7370[21]), .\delay_r_23__N_1178[21] (delay_r_23__N_1178_adj_7427[21]), 
            .\dout_r_23__N_5681[21] (dout_r_23__N_5681[21]), .\op_i_23__N_1154[12] (op_i_23__N_1154_adj_7371[12]), 
            .\delay_i_23__N_1202[12] (delay_i_23__N_1202_adj_7428[12]), .\dout_i_23__N_5777[12] (dout_i_23__N_5777[12]), 
            .\op_r_23__N_1226[0] (op_r_23__N_1226_adj_7432[0]), .\op_r_23__N_1226[1] (op_r_23__N_1226_adj_7432[1]), 
            .\op_r_23__N_1226[2] (op_r_23__N_1226_adj_7432[2]), .\op_r_23__N_1226[3] (op_r_23__N_1226_adj_7432[3]), 
            .\op_r_23__N_1226[4] (op_r_23__N_1226_adj_7432[4]), .\op_r_23__N_1226[5] (op_r_23__N_1226_adj_7432[5]), 
            .\op_r_23__N_1226[6] (op_r_23__N_1226_adj_7432[6]), .\op_r_23__N_1226[7] (op_r_23__N_1226_adj_7432[7]), 
            .\op_r_23__N_1226[8] (op_r_23__N_1226_adj_7432[8]), .\op_r_23__N_1226[9] (op_r_23__N_1226_adj_7432[9]), 
            .\op_r_23__N_1226[10] (op_r_23__N_1226_adj_7432[10]), .\op_r_23__N_1226[11] (op_r_23__N_1226_adj_7432[11]), 
            .\op_r_23__N_1226[12] (op_r_23__N_1226_adj_7432[12]), .\op_r_23__N_1226[13] (op_r_23__N_1226_adj_7432[13]), 
            .\op_r_23__N_1226[14] (op_r_23__N_1226_adj_7432[14]), .\op_r_23__N_1226[15] (op_r_23__N_1226_adj_7432[15]), 
            .\op_r_23__N_1226[16] (op_r_23__N_1226_adj_7432[16]), .\op_r_23__N_1226[17] (op_r_23__N_1226_adj_7432[17]), 
            .\op_r_23__N_1226[18] (op_r_23__N_1226_adj_7432[18]), .\op_r_23__N_1226[19] (op_r_23__N_1226_adj_7432[19]), 
            .\op_r_23__N_1226[20] (op_r_23__N_1226_adj_7432[20]), .\op_r_23__N_1226[21] (op_r_23__N_1226_adj_7432[21]), 
            .\op_r_23__N_1226[22] (op_r_23__N_1226_adj_7432[22]), .\op_r_23__N_1226[23] (op_r_23__N_1226_adj_7432[23]), 
            .\op_r_23__N_1226[24] (op_r_23__N_1226_adj_7432[24]), .\op_r_23__N_1226[25] (op_r_23__N_1226_adj_7432[25]), 
            .\op_r_23__N_1226[26] (op_r_23__N_1226_adj_7432[26]), .\op_r_23__N_1226[27] (op_r_23__N_1226_adj_7432[27]), 
            .\op_r_23__N_1226[28] (op_r_23__N_1226_adj_7432[28]), .\op_r_23__N_1226[29] (op_r_23__N_1226_adj_7432[29]), 
            .\op_r_23__N_1226[30] (op_r_23__N_1226_adj_7432[30]), .\op_r_23__N_1226[31] (op_r_23__N_1226_adj_7432[31]), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n12170(n12170), .n12171(n12171), 
            .n12172(n12172), .n12173(n12173), .n12174(n12174), .n12175(n12175), 
            .n12176(n12176), .\rom2_w_r[8] (rom2_w_r[8]), .n12152(n12152), 
            .n12153(n12153), .n12154(n12154), .n12155(n12155), .n12156(n12156), 
            .n12157(n12157), .n12158(n12158), .n12159(n12159), .n12160(n12160), 
            .n12161(n12161), .n12162(n12162), .n12163(n12163), .n12164(n12164), 
            .n12165(n12165), .n12166(n12166), .n12167(n12167), .n12168(n12168), 
            .n12169(n12169), .\op_r_23__N_1106[15] (op_r_23__N_1106_adj_7370[15]), 
            .\delay_r_23__N_1178[15] (delay_r_23__N_1178_adj_7427[15]), .\dout_r_23__N_5681[15] (dout_r_23__N_5681[15]), 
            .\op_r_23__N_1106[13] (op_r_23__N_1106_adj_7370[13]), .\delay_r_23__N_1178[13] (delay_r_23__N_1178_adj_7427[13]), 
            .\dout_r_23__N_5681[13] (dout_r_23__N_5681[13]), .\op_r_23__N_1106[12] (op_r_23__N_1106_adj_7370[12]), 
            .\delay_r_23__N_1178[12] (delay_r_23__N_1178_adj_7427[12]), .\dout_r_23__N_5681[12] (dout_r_23__N_5681[12]), 
            .\op_i_23__N_1154[11] (op_i_23__N_1154_adj_7371[11]), .\delay_i_23__N_1202[11] (delay_i_23__N_1202_adj_7428[11]), 
            .\dout_i_23__N_5777[11] (dout_i_23__N_5777[11]), .\op_r_23__N_1106[20] (op_r_23__N_1106_adj_7370[20]), 
            .\delay_r_23__N_1178[20] (delay_r_23__N_1178_adj_7427[20]), .\dout_r_23__N_5681[20] (dout_r_23__N_5681[20]), 
            .\op_i_23__N_1154[10] (op_i_23__N_1154_adj_7371[10]), .\delay_i_23__N_1202[10] (delay_i_23__N_1202_adj_7428[10]), 
            .\dout_i_23__N_5777[10] (dout_i_23__N_5777[10]), .n34795(n34795), 
            .n114(n114), .shift_2_dout_i({shift_2_dout_i}), .\op_r_23__N_1268[0] (op_r_23__N_1268_adj_7430[0]), 
            .\op_r_23__N_1268[1] (op_r_23__N_1268_adj_7430[1]), .\op_r_23__N_1268[2] (op_r_23__N_1268_adj_7430[2]), 
            .\op_r_23__N_1268[3] (op_r_23__N_1268_adj_7430[3]), .\op_r_23__N_1268[4] (op_r_23__N_1268_adj_7430[4]), 
            .\op_r_23__N_1268[5] (op_r_23__N_1268_adj_7430[5]), .\op_r_23__N_1268[6] (op_r_23__N_1268_adj_7430[6]), 
            .\op_r_23__N_1268[7] (op_r_23__N_1268_adj_7430[7]), .\op_r_23__N_1268[8] (op_r_23__N_1268_adj_7430[8]), 
            .\op_r_23__N_1268[9] (op_r_23__N_1268_adj_7430[9]), .\op_r_23__N_1268[10] (op_r_23__N_1268_adj_7430[10]), 
            .\op_r_23__N_1268[11] (op_r_23__N_1268_adj_7430[11]), .\op_r_23__N_1268[12] (op_r_23__N_1268_adj_7430[12]), 
            .\op_r_23__N_1268[13] (op_r_23__N_1268_adj_7430[13]), .\op_r_23__N_1268[14] (op_r_23__N_1268_adj_7430[14]), 
            .\op_r_23__N_1268[15] (op_r_23__N_1268_adj_7430[15]), .\op_r_23__N_1268[16] (op_r_23__N_1268_adj_7430[16]), 
            .\op_r_23__N_1268[17] (op_r_23__N_1268_adj_7430[17]), .\op_r_23__N_1268[18] (op_r_23__N_1268_adj_7430[18]), 
            .\op_r_23__N_1268[19] (op_r_23__N_1268_adj_7430[19]), .\op_r_23__N_1268[20] (op_r_23__N_1268_adj_7430[20]), 
            .\op_r_23__N_1268[21] (op_r_23__N_1268_adj_7430[21]), .\op_r_23__N_1268[22] (op_r_23__N_1268_adj_7430[22]), 
            .\op_r_23__N_1268[23] (op_r_23__N_1268_adj_7430[23]), .\op_r_23__N_1268[24] (op_r_23__N_1268_adj_7430[24]), 
            .\op_r_23__N_1268[25] (op_r_23__N_1268_adj_7430[25]), .\op_r_23__N_1268[26] (op_r_23__N_1268_adj_7430[26]), 
            .\op_r_23__N_1268[27] (op_r_23__N_1268_adj_7430[27]), .\op_r_23__N_1268[28] (op_r_23__N_1268_adj_7430[28]), 
            .\op_r_23__N_1268[29] (op_r_23__N_1268_adj_7430[29]), .\op_r_23__N_1268[30] (op_r_23__N_1268_adj_7430[30]), 
            .\op_r_23__N_1268[31] (op_r_23__N_1268_adj_7430[31]), .n8977(n8977), 
            .n8976(n8976), .n8975(n8975), .n8974(n8974), .n8973(n8973), 
            .n8972(n8972), .n8971(n8971), .n8970(n8970), .n8969(n8969), 
            .n8968(n8968), .n8967(n8967), .n8966(n8966), .n8965(n8965), 
            .n8964(n8964), .n8963(n8963), .n8962(n8962), .n8961(n8961), 
            .n8960(n8960), .n8959(n8959), .n8958(n8958), .n8957(n8957), 
            .n8956(n8956), .n8955(n8955), .n8954(n8954), .n8953(n8953), 
            .n8952(n8952), .\op_i_23__N_1154[19] (op_i_23__N_1154_adj_7371[19]), 
            .\delay_i_23__N_1202[19] (delay_i_23__N_1202_adj_7428[19]), .\dout_i_23__N_5777[19] (dout_i_23__N_5777[19]), 
            .n319(n319_adj_6944), .\rom4_w_i[12] (rom4_w_i[12]), .n114_adj_33(n114_adj_7263), 
            .n11126(n11126), .n11127(n11127), .n11128(n11128), .n11129(n11129), 
            .n11130(n11130), .n11131(n11131), .n11132(n11132), .n11133(n11133), 
            .n11134(n11134), .n11135(n11135), .n11136(n11136), .n11137(n11137), 
            .n11138(n11138), .n11139(n11139), .n11140(n11140), .n11141(n11141), 
            .n11142(n11142), .n11143(n11143), .n120(n120), .n126(n126), 
            .\op_i_23__N_1310[0] (op_i_23__N_1310_adj_7435[0]), .n123(n123), 
            .n117(n117), .n111(n111), .\op_i_23__N_1310[2] (op_i_23__N_1310_adj_7435[2]), 
            .\op_i_23__N_1310[3] (op_i_23__N_1310_adj_7435[3]), .\op_i_23__N_1310[4] (op_i_23__N_1310_adj_7435[4]), 
            .\op_i_23__N_1310[5] (op_i_23__N_1310_adj_7435[5]), .n89(n89_adj_7261), 
            .n87(n87_adj_7259), .n88(n88_adj_7260), .n85(n85_adj_7257), 
            .n86(n86_adj_7258), .n83(n83_adj_7255), .n84(n84_adj_7256), 
            .n81(n81_adj_7253), .n82(n82_adj_7254), .n79(n79_adj_7251), 
            .n80(n80_adj_7252), .n77(n77_adj_7249), .n78(n78_adj_7250), 
            .n75(n75_adj_7247), .n76(n76_adj_7248), .n73(n73_adj_7245), 
            .n74(n74_adj_7246), .n71(n71_adj_7243), .n72(n72_adj_7244), 
            .n69(n69_adj_7241), .n70(n70_adj_7242), .n67(n67_adj_7239), 
            .n68(n68_adj_7240), .n65(n65), .n66(n66_adj_7238), .\op_i_23__N_1310[1] (op_i_23__N_1310_adj_7435[1]), 
            .n120_adj_34(n120_adj_7265), .n126_adj_35(n126_adj_7267), .n34777(n34777), 
            .\op_i_23__N_1310[0]_adj_36 (op_i_23__N_1310_adj_7380[0]), .n123_adj_37(n123_adj_7266), 
            .n117_adj_38(n117_adj_7264), .n111_adj_39(n111_adj_7262), .\op_i_23__N_1310[2]_adj_40 (op_i_23__N_1310_adj_7380[2]), 
            .\op_i_23__N_1310[3]_adj_41 (op_i_23__N_1310_adj_7380[3]), .\op_i_23__N_1310[4]_adj_42 (op_i_23__N_1310_adj_7380[4]), 
            .\op_i_23__N_1310[5]_adj_43 (op_i_23__N_1310_adj_7380[5]), .n89_adj_44(n89_adj_7291), 
            .n87_adj_45(n87_adj_7289), .n88_adj_46(n88_adj_7290), .n85_adj_47(n85_adj_7287), 
            .n86_adj_48(n86_adj_7288), .n83_adj_49(n83_adj_7285), .n84_adj_50(n84_adj_7286), 
            .n81_adj_51(n81_adj_7283), .n82_adj_52(n82_adj_7284), .n79_adj_53(n79_adj_7281), 
            .n80_adj_54(n80_adj_7282), .n77_adj_55(n77_adj_7279), .n78_adj_56(n78_adj_7280), 
            .n75_adj_57(n75_adj_7277), .n76_adj_58(n76_adj_7278), .n73_adj_59(n73_adj_7275), 
            .n74_adj_60(n74_adj_7276), .n71_adj_61(n71_adj_7273), .n72_adj_62(n72_adj_7274), 
            .n69_adj_63(n69_adj_7271), .n70_adj_64(n70_adj_7272), .n67_adj_65(n67_adj_7269), 
            .n68_adj_66(n68_adj_7270), .n65_adj_67(n65_adj_6772), .n66_adj_68(n66_adj_7268), 
            .\op_i_23__N_1310[1]_adj_69 (op_i_23__N_1310_adj_7380[1]), .\op_r_23__N_1106[19] (op_r_23__N_1106_adj_7370[19]), 
            .\delay_r_23__N_1178[19] (delay_r_23__N_1178_adj_7427[19]), .\dout_r_23__N_5681[19] (dout_r_23__N_5681[19]), 
            .\op_r_23__N_1106[11] (op_r_23__N_1106_adj_7370[11]), .\delay_r_23__N_1178[11] (delay_r_23__N_1178_adj_7427[11]), 
            .\dout_r_23__N_5681[11] (dout_r_23__N_5681[11]), .\op_r_23__N_1106[10] (op_r_23__N_1106_adj_7370[10]), 
            .\delay_r_23__N_1178[10] (delay_r_23__N_1178_adj_7427[10]), .\dout_r_23__N_5681[10] (dout_r_23__N_5681[10]), 
            .\op_i_23__N_1154[9] (op_i_23__N_1154_adj_7371[9]), .\delay_i_23__N_1202[9] (delay_i_23__N_1202_adj_7428[9]), 
            .\dout_i_23__N_5777[9] (dout_i_23__N_5777[9]), .\op_r_23__N_1106[18] (op_r_23__N_1106_adj_7370[18]), 
            .\delay_r_23__N_1178[18] (delay_r_23__N_1178_adj_7427[18]), .\dout_r_23__N_5681[18] (dout_r_23__N_5681[18]), 
            .\op_i_23__N_1154[8] (op_i_23__N_1154_adj_7371[8]), .\delay_i_23__N_1202[8] (delay_i_23__N_1202_adj_7428[8]), 
            .\dout_i_23__N_5777[8] (dout_i_23__N_5777[8]), .\op_r_23__N_1106[9] (op_r_23__N_1106_adj_7370[9]), 
            .\delay_r_23__N_1178[9] (delay_r_23__N_1178_adj_7427[9]), .\dout_r_23__N_5681[9] (dout_r_23__N_5681[9]), 
            .\op_r_23__N_1106[8] (op_r_23__N_1106_adj_7370[8]), .\delay_r_23__N_1178[8] (delay_r_23__N_1178_adj_7427[8]), 
            .\dout_r_23__N_5681[8] (dout_r_23__N_5681[8]), .\op_i_23__N_1154[7] (op_i_23__N_1154_adj_7371[7]), 
            .\delay_i_23__N_1202[7] (delay_i_23__N_1202_adj_7428[7]), .\dout_i_23__N_5777[7] (dout_i_23__N_5777[7]), 
            .\op_i_23__N_1154[6] (op_i_23__N_1154_adj_7371[6]), .\delay_i_23__N_1202[6] (delay_i_23__N_1202_adj_7428[6]), 
            .\dout_i_23__N_5777[6] (dout_i_23__N_5777[6]), .\op_i_23__N_1154[17] (op_i_23__N_1154_adj_7371[17]), 
            .\delay_i_23__N_1202[17] (delay_i_23__N_1202_adj_7428[17]), .\dout_i_23__N_5777[17] (dout_i_23__N_5777[17]), 
            .\op_i_23__N_1154[23] (op_i_23__N_1154_adj_7371[23]), .\delay_i_23__N_1202[23] (delay_i_23__N_1202_adj_7428[23]), 
            .\dout_i_23__N_5777[23] (dout_i_23__N_5777[23]), .\op_r_23__N_1106[23] (op_r_23__N_1106_adj_7370[23]), 
            .\delay_r_23__N_1178[23] (delay_r_23__N_1178_adj_7427[23]), .\dout_r_23__N_5681[23] (dout_r_23__N_5681[23]), 
            .\op_r_23__N_1106[22] (op_r_23__N_1106_adj_7370[22]), .\delay_r_23__N_1178[22] (delay_r_23__N_1178_adj_7427[22]), 
            .\dout_r_23__N_5681[22] (dout_r_23__N_5681[22]), .\op_i_23__N_1154[21] (op_i_23__N_1154_adj_7371[21]), 
            .\delay_i_23__N_1202[21] (delay_i_23__N_1202_adj_7428[21]), .\dout_i_23__N_5777[21] (dout_i_23__N_5777[21]), 
            .\op_i_23__N_1154[16] (op_i_23__N_1154_adj_7371[16]), .\delay_i_23__N_1202[16] (delay_i_23__N_1202_adj_7428[16]), 
            .\dout_i_23__N_5777[16] (dout_i_23__N_5777[16]), .\op_i_23__N_1154[20] (op_i_23__N_1154_adj_7371[20]), 
            .\delay_i_23__N_1202[20] (delay_i_23__N_1202_adj_7428[20]), .\dout_i_23__N_5777[20] (dout_i_23__N_5777[20]), 
            .\op_i_23__N_1154[5] (op_i_23__N_1154_adj_7371[5]), .\delay_i_23__N_1202[5] (delay_i_23__N_1202_adj_7428[5]), 
            .\dout_i_23__N_5777[5] (dout_i_23__N_5777[5]), .\op_i_23__N_1154[4] (op_i_23__N_1154_adj_7371[4]), 
            .\delay_i_23__N_1202[4] (delay_i_23__N_1202_adj_7428[4]), .\dout_i_23__N_5777[4] (dout_i_23__N_5777[4]), 
            .\op_i_23__N_1154[3] (op_i_23__N_1154_adj_7371[3]), .\delay_i_23__N_1202[3] (delay_i_23__N_1202_adj_7428[3]), 
            .\dout_i_23__N_5777[3] (dout_i_23__N_5777[3]), .\op_i_23__N_1154[22] (op_i_23__N_1154_adj_7371[22]), 
            .\delay_i_23__N_1202[22] (delay_i_23__N_1202_adj_7428[22]), .\dout_i_23__N_5777[22] (dout_i_23__N_5777[22]), 
            .\op_r_23__N_1106[7] (op_r_23__N_1106_adj_7370[7]), .\delay_r_23__N_1178[7] (delay_r_23__N_1178_adj_7427[7]), 
            .\dout_r_23__N_5681[7] (dout_r_23__N_5681[7]), .\op_r_23__N_1106[6] (op_r_23__N_1106_adj_7370[6]), 
            .\delay_r_23__N_1178[6] (delay_r_23__N_1178_adj_7427[6]), .\dout_r_23__N_5681[6] (dout_r_23__N_5681[6]), 
            .\op_r_23__N_1106[5] (op_r_23__N_1106_adj_7370[5]), .\delay_r_23__N_1178[5] (delay_r_23__N_1178_adj_7427[5]), 
            .\dout_r_23__N_5681[5] (dout_r_23__N_5681[5]), .\op_r_23__N_1106[4] (op_r_23__N_1106_adj_7370[4]), 
            .\delay_r_23__N_1178[4] (delay_r_23__N_1178_adj_7427[4]), .\dout_r_23__N_5681[4] (dout_r_23__N_5681[4]), 
            .\op_r_23__N_1106[17] (op_r_23__N_1106_adj_7370[17]), .\delay_r_23__N_1178[17] (delay_r_23__N_1178_adj_7427[17]), 
            .\dout_r_23__N_5681[17] (dout_r_23__N_5681[17]), .\op_r_23__N_1106[3] (op_r_23__N_1106_adj_7370[3]), 
            .\delay_r_23__N_1178[3] (delay_r_23__N_1178_adj_7427[3]), .\dout_r_23__N_5681[3] (dout_r_23__N_5681[3]), 
            .\op_r_23__N_1106[2] (op_r_23__N_1106_adj_7370[2]), .\delay_r_23__N_1178[2] (delay_r_23__N_1178_adj_7427[2]), 
            .\dout_r_23__N_5681[2] (dout_r_23__N_5681[2]), .\op_r_23__N_1106[16] (op_r_23__N_1106_adj_7370[16]), 
            .\delay_r_23__N_1178[16] (delay_r_23__N_1178_adj_7427[16]), .\dout_r_23__N_5681[16] (dout_r_23__N_5681[16]), 
            .\op_r_23__N_1106[1] (op_r_23__N_1106_adj_7370[1]), .\delay_r_23__N_1178[1] (delay_r_23__N_1178_adj_7427[1]), 
            .\dout_r_23__N_5681[1] (dout_r_23__N_5681[1]), .\op_i_23__N_1154[15] (op_i_23__N_1154_adj_7371[15]), 
            .\delay_i_23__N_1202[15] (delay_i_23__N_1202_adj_7428[15]), .\dout_i_23__N_5777[15] (dout_i_23__N_5777[15]), 
            .\op_i_23__N_1154[14] (op_i_23__N_1154_adj_7371[14]), .\delay_i_23__N_1202[14] (delay_i_23__N_1202_adj_7428[14]), 
            .\dout_i_23__N_5777[14] (dout_i_23__N_5777[14])) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(183[8] 196[2])
    LUT4 i15595_3_lut (.A(\result_r[18] [9]), .B(\result_r[19] [9]), .C(y_1_delay[0]), 
         .Z(n33979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15595_3_lut.init = 16'hcaca;
    LUT4 i2655_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [10]), 
         .D(out_i[18]), .Z(result_i_ns_0__15__N_517[490])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2655_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15575 (.BLUT(n33947), .ALUT(n33948), .C0(y_1_delay[1]), .Z(n33959));
    LUT4 i15094_3_lut (.A(\result_i[8] [10]), .B(\result_i[9] [10]), .C(y_1_delay[0]), 
         .Z(n33478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15094_3_lut.init = 16'hcaca;
    LUT4 i854_2_lut_rep_440 (.A(count_y[1]), .B(count_y[0]), .Z(n34802)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i854_2_lut_rep_440.init = 16'heeee;
    LUT4 i861_2_lut_rep_408_3_lut (.A(count_y[1]), .B(count_y[0]), .C(count_y[2]), 
         .Z(n34770)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(47[14:56])
    defparam i861_2_lut_rep_408_3_lut.init = 16'hfefe;
    PFUMX i15576 (.BLUT(n33949), .ALUT(n33950), .C0(y_1_delay[1]), .Z(n33960));
    LUT4 i2647_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [11]), 
         .D(out_i[19]), .Z(result_i_ns_0__15__N_517[491])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2647_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i2639_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_i[1] [12]), 
         .D(out_i[20]), .Z(result_i_ns_0__15__N_517[492])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i2639_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15577 (.BLUT(n33951), .ALUT(n33952), .C0(y_1_delay[1]), .Z(n33961));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i15594_3_lut (.A(\result_r[16] [9]), .B(\result_r[17] [9]), .C(y_1_delay[0]), 
         .Z(n33978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15594_3_lut.init = 16'hcaca;
    PFUMX i15578 (.BLUT(n33953), .ALUT(n33954), .C0(y_1_delay[1]), .Z(n33962));
    LUT4 i6761_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [8]), 
         .D(out_r[16]), .Z(result_r_ns_0__15__N_3[488])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6761_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i15230 (.BLUT(n33598), .ALUT(n33599), .C0(y_1_delay[1]), .Z(n33614));
    PFUMX i15231 (.BLUT(n33600), .ALUT(n33601), .C0(y_1_delay[1]), .Z(n33615));
    PFUMX i15232 (.BLUT(n33602), .ALUT(n33603), .C0(y_1_delay[1]), .Z(n33616));
    PFUMX i15044 (.BLUT(n33412), .ALUT(n33413), .C0(y_1_delay[1]), .Z(n33428));
    PFUMX i15233 (.BLUT(n33604), .ALUT(n33605), .C0(y_1_delay[1]), .Z(n33617));
    PFUMX i15602 (.BLUT(n33970), .ALUT(n33971), .C0(y_1_delay[1]), .Z(n33986));
    PFUMX i15603 (.BLUT(n33972), .ALUT(n33973), .C0(y_1_delay[1]), .Z(n33987));
    PFUMX i15234 (.BLUT(n33606), .ALUT(n33607), .C0(y_1_delay[1]), .Z(n33618));
    PFUMX i15235 (.BLUT(n33608), .ALUT(n33609), .C0(y_1_delay[1]), .Z(n33619));
    PFUMX i15045 (.BLUT(n33414), .ALUT(n33415), .C0(y_1_delay[1]), .Z(n33429));
    LUT4 i6753_3_lut_4_lut (.A(n34741), .B(n34715), .C(\result_r[1] [9]), 
         .D(out_r[17]), .Z(result_r_ns_0__15__N_3[489])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(312[9] 444[16])
    defparam i6753_3_lut_4_lut.init = 16'hf2d0;
    shift_8 shift_8 (.clk_c(clk_c), .clk_c_enable_1419(clk_c_enable_1419), 
            .\dout_i_23__N_4670[0] (dout_i_23__N_4670[0]), .\dout_r_23__N_4286[0] (dout_r_23__N_4286[0]), 
            .valid(valid), .clk_c_enable_2310(clk_c_enable_2310), .VCC_net(VCC_net), 
            .\dout_i_23__N_4670[1] (dout_i_23__N_4670[1]), .\dout_i_23__N_4670[2] (dout_i_23__N_4670[2]), 
            .\dout_i_23__N_4670[3] (dout_i_23__N_4670[3]), .\dout_i_23__N_4670[4] (dout_i_23__N_4670[4]), 
            .\dout_i_23__N_4670[5] (dout_i_23__N_4670[5]), .\dout_i_23__N_4670[6] (dout_i_23__N_4670[6]), 
            .\dout_i_23__N_4670[7] (dout_i_23__N_4670[7]), .\dout_i_23__N_4670[8] (dout_i_23__N_4670[8]), 
            .\dout_i_23__N_4670[9] (dout_i_23__N_4670[9]), .\dout_i_23__N_4670[10] (dout_i_23__N_4670[10]), 
            .\dout_i_23__N_4670[11] (dout_i_23__N_4670[11]), .\dout_i_23__N_4670[12] (dout_i_23__N_4670[12]), 
            .\dout_i_23__N_4670[13] (dout_i_23__N_4670[13]), .\dout_i_23__N_4670[14] (dout_i_23__N_4670[14]), 
            .\dout_i_23__N_4670[15] (dout_i_23__N_4670[15]), .\dout_i_23__N_4670[16] (dout_i_23__N_4670[16]), 
            .\dout_i_23__N_4670[17] (dout_i_23__N_4670[17]), .\dout_i_23__N_4670[18] (dout_i_23__N_4670[18]), 
            .\dout_i_23__N_4670[19] (dout_i_23__N_4670[19]), .\dout_i_23__N_4670[20] (dout_i_23__N_4670[20]), 
            .\dout_i_23__N_4670[21] (dout_i_23__N_4670[21]), .\dout_i_23__N_4670[22] (dout_i_23__N_4670[22]), 
            .\dout_i_23__N_4670[23] (dout_i_23__N_4670[23]), .\dout_r_23__N_4286[1] (dout_r_23__N_4286[1]), 
            .\dout_r_23__N_4286[2] (dout_r_23__N_4286[2]), .\dout_r_23__N_4286[3] (dout_r_23__N_4286[3]), 
            .\dout_r_23__N_4286[4] (dout_r_23__N_4286[4]), .\dout_r_23__N_4286[5] (dout_r_23__N_4286[5]), 
            .\dout_r_23__N_4286[6] (dout_r_23__N_4286[6]), .\dout_r_23__N_4286[7] (dout_r_23__N_4286[7]), 
            .\dout_r_23__N_4286[8] (dout_r_23__N_4286[8]), .\dout_r_23__N_4286[9] (dout_r_23__N_4286[9]), 
            .\dout_r_23__N_4286[10] (dout_r_23__N_4286[10]), .\dout_r_23__N_4286[11] (dout_r_23__N_4286[11]), 
            .\dout_r_23__N_4286[12] (dout_r_23__N_4286[12]), .\dout_r_23__N_4286[13] (dout_r_23__N_4286[13]), 
            .\dout_r_23__N_4286[14] (dout_r_23__N_4286[14]), .\dout_r_23__N_4286[15] (dout_r_23__N_4286[15]), 
            .\dout_r_23__N_4286[16] (dout_r_23__N_4286[16]), .\dout_r_23__N_4286[17] (dout_r_23__N_4286[17]), 
            .\dout_r_23__N_4286[18] (dout_r_23__N_4286[18]), .\dout_r_23__N_4286[19] (dout_r_23__N_4286[19]), 
            .\dout_r_23__N_4286[20] (dout_r_23__N_4286[20]), .\dout_r_23__N_4286[21] (dout_r_23__N_4286[21]), 
            .\dout_r_23__N_4286[22] (dout_r_23__N_4286[22]), .\dout_r_23__N_4286[23] (dout_r_23__N_4286[23]), 
            .shift_8_dout_i({shift_8_dout_i}), .shift_8_dout_r({shift_8_dout_r})) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(130[9] 137[2])
    LUT4 i15590_3_lut (.A(\result_r[8] [9]), .B(\result_r[9] [9]), .C(y_1_delay[0]), 
         .Z(n33974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15590_3_lut.init = 16'hcaca;
    PFUMX i15046 (.BLUT(n33416), .ALUT(n33417), .C0(y_1_delay[1]), .Z(n33430));
    PFUMX i15236 (.BLUT(n33610), .ALUT(n33611), .C0(y_1_delay[1]), .Z(n33620));
    radix2 radix_no5 (.dout_i_23__N_5974({dout_i_23__N_5974}), .GND_net(GND_net), 
           .VCC_net(VCC_net), .clk_c(clk_c), .n34738(n34738), .rst_n_N_2(rst_n_N_2), 
           .\op_r_23__N_1226[0] (op_r_23__N_1226_adj_7488[0]), .\op_r_23__N_1226[1] (op_r_23__N_1226_adj_7488[1]), 
           .\op_r_23__N_1226[2] (op_r_23__N_1226_adj_7488[2]), .\op_r_23__N_1226[3] (op_r_23__N_1226_adj_7488[3]), 
           .\op_r_23__N_1226[4] (op_r_23__N_1226_adj_7488[4]), .\op_r_23__N_1226[5] (op_r_23__N_1226_adj_7488[5]), 
           .\op_r_23__N_1226[6] (op_r_23__N_1226_adj_7488[6]), .\op_r_23__N_1226[7] (op_r_23__N_1226_adj_7488[7]), 
           .\op_r_23__N_1226[8] (op_r_23__N_1226_adj_7488[8]), .\op_r_23__N_1226[9] (op_r_23__N_1226_adj_7488[9]), 
           .\op_r_23__N_1226[10] (op_r_23__N_1226_adj_7488[10]), .\op_r_23__N_1226[11] (op_r_23__N_1226_adj_7488[11]), 
           .\op_r_23__N_1226[12] (op_r_23__N_1226_adj_7488[12]), .\op_r_23__N_1226[13] (op_r_23__N_1226_adj_7488[13]), 
           .\op_r_23__N_1226[14] (op_r_23__N_1226_adj_7488[14]), .\op_r_23__N_1226[15] (op_r_23__N_1226_adj_7488[15]), 
           .\op_r_23__N_1226[16] (op_r_23__N_1226_adj_7488[16]), .\op_r_23__N_1226[17] (op_r_23__N_1226_adj_7488[17]), 
           .\op_r_23__N_1226[18] (op_r_23__N_1226_adj_7488[18]), .\op_r_23__N_1226[19] (op_r_23__N_1226_adj_7488[19]), 
           .\op_r_23__N_1226[20] (op_r_23__N_1226_adj_7488[20]), .\op_r_23__N_1226[21] (op_r_23__N_1226_adj_7488[21]), 
           .\op_r_23__N_1226[22] (op_r_23__N_1226_adj_7488[22]), .\op_r_23__N_1226[23] (op_r_23__N_1226_adj_7488[23]), 
           .\op_r_23__N_1226[24] (op_r_23__N_1226_adj_7488[24]), .\op_r_23__N_1226[25] (op_r_23__N_1226_adj_7488[25]), 
           .\op_r_23__N_1226[26] (op_r_23__N_1226_adj_7488[26]), .\op_r_23__N_1226[27] (op_r_23__N_1226_adj_7488[27]), 
           .\op_r_23__N_1226[28] (op_r_23__N_1226_adj_7488[28]), .\op_r_23__N_1226[29] (op_r_23__N_1226_adj_7488[29]), 
           .\op_r_23__N_1226[30] (op_r_23__N_1226_adj_7488[30]), .\op_r_23__N_1226[31] (op_r_23__N_1226_adj_7488[31]), 
           .\op_i_23__N_1310[0] (op_i_23__N_1310_adj_7491[0]), .\op_i_23__N_1310[1] (op_i_23__N_1310_adj_7491[1]), 
           .\op_i_23__N_1310[2] (op_i_23__N_1310_adj_7491[2]), .\op_i_23__N_1310[3] (op_i_23__N_1310_adj_7491[3]), 
           .\op_i_23__N_1310[4] (op_i_23__N_1310_adj_7491[4]), .\op_i_23__N_1310[5] (op_i_23__N_1310_adj_7491[5]), 
           .n89(n89_adj_6552), .n88(n88_adj_6553), .n87(n87_adj_6554), 
           .n86(n86_adj_6555), .n85(n85_adj_6556), .n84(n84_adj_6557), 
           .n83(n83_adj_6558), .n82(n82_adj_6559), .n81(n81_adj_6560), 
           .n80(n80_adj_6561), .n79(n79_adj_6562), .n78(n78_adj_6563), 
           .n77(n77_adj_6564), .n76(n76_adj_6565), .n75(n75_adj_6566), 
           .n74(n74_adj_6567), .n73(n73_adj_6568), .n72(n72_adj_6569), 
           .n71(n71_adj_6570), .n70(n70_adj_6571), .n69(n69_adj_6572), 
           .n68(n68_adj_6573), .n67(n67_adj_6574), .n66(n66_adj_6575), 
           .n65(n65_adj_6576), .n11556(n11556), .n11557(n11557), .n11558(n11558), 
           .n11559(n11559), .n11560(n11560), .n11561(n11561), .n12083(n12083), 
           .n12084(n12084), .n12085(n12085), .n12086(n12086), .n12087(n12087), 
           .n12088(n12088), .n12089(n12089), .n12065(n12065), .n12066(n12066), 
           .n12067(n12067), .n12068(n12068), .n12069(n12069), .n12070(n12070), 
           .n12071(n12071), .n12072(n12072), .n12073(n12073), .n12074(n12074), 
           .n12075(n12075), .n12076(n12076), .n12077(n12077), .n12078(n12078), 
           .n12079(n12079), .n12080(n12080), .n12081(n12081), .n12082(n12082), 
           .\op_r_23__N_1268[0] (op_r_23__N_1268_adj_7486[0]), .\op_r_23__N_1268[1] (op_r_23__N_1268_adj_7486[1]), 
           .\op_r_23__N_1268[2] (op_r_23__N_1268_adj_7486[2]), .\op_r_23__N_1268[3] (op_r_23__N_1268_adj_7486[3]), 
           .\op_r_23__N_1268[4] (op_r_23__N_1268_adj_7486[4]), .\op_r_23__N_1268[5] (op_r_23__N_1268_adj_7486[5]), 
           .\op_r_23__N_1268[6] (op_r_23__N_1268_adj_7486[6]), .\op_r_23__N_1268[7] (op_r_23__N_1268_adj_7486[7]), 
           .\op_r_23__N_1268[8] (op_r_23__N_1268_adj_7486[8]), .\op_r_23__N_1268[9] (op_r_23__N_1268_adj_7486[9]), 
           .\op_r_23__N_1268[10] (op_r_23__N_1268_adj_7486[10]), .\op_r_23__N_1268[11] (op_r_23__N_1268_adj_7486[11]), 
           .\op_r_23__N_1268[12] (op_r_23__N_1268_adj_7486[12]), .\op_r_23__N_1268[13] (op_r_23__N_1268_adj_7486[13]), 
           .\op_r_23__N_1268[14] (op_r_23__N_1268_adj_7486[14]), .\op_r_23__N_1268[15] (op_r_23__N_1268_adj_7486[15]), 
           .\op_r_23__N_1268[16] (op_r_23__N_1268_adj_7486[16]), .\op_r_23__N_1268[17] (op_r_23__N_1268_adj_7486[17]), 
           .\op_r_23__N_1268[18] (op_r_23__N_1268_adj_7486[18]), .\op_r_23__N_1268[19] (op_r_23__N_1268_adj_7486[19]), 
           .\op_r_23__N_1268[20] (op_r_23__N_1268_adj_7486[20]), .\op_r_23__N_1268[21] (op_r_23__N_1268_adj_7486[21]), 
           .\op_r_23__N_1268[22] (op_r_23__N_1268_adj_7486[22]), .\op_r_23__N_1268[23] (op_r_23__N_1268_adj_7486[23]), 
           .\op_r_23__N_1268[24] (op_r_23__N_1268_adj_7486[24]), .\op_r_23__N_1268[25] (op_r_23__N_1268_adj_7486[25]), 
           .\op_r_23__N_1268[26] (op_r_23__N_1268_adj_7486[26]), .\op_r_23__N_1268[27] (op_r_23__N_1268_adj_7486[27]), 
           .\op_r_23__N_1268[28] (op_r_23__N_1268_adj_7486[28]), .\op_r_23__N_1268[29] (op_r_23__N_1268_adj_7486[29]), 
           .\op_r_23__N_1268[30] (op_r_23__N_1268_adj_7486[30]), .\op_r_23__N_1268[31] (op_r_23__N_1268_adj_7486[31]), 
           .n9105(n9105), .n9104(n9104), .n9103(n9103), .n9102(n9102), 
           .n9101(n9101), .n9100(n9100), .n9099(n9099), .n9098(n9098), 
           .n9097(n9097), .n9096(n9096), .n9095(n9095), .n9094(n9094), 
           .n9093(n9093), .n9092(n9092), .n9091(n9091), .n9090(n9090), 
           .n9089(n9089), .n9088(n9088), .n9087(n9087), .n9086(n9086), 
           .n9085(n9085), .n9084(n9084), .n9083(n9083), .n9082(n9082), 
           .n9081(n9081), .n9080(n9080), .n319(n319_adj_7163), .n11562(n11562), 
           .n11563(n11563), .n11564(n11564), .n11565(n11565), .n11566(n11566), 
           .n11567(n11567), .n11568(n11568), .n11569(n11569), .n11570(n11570), 
           .n11571(n11571), .n11572(n11572), .n11573(n11573), .n11574(n11574), 
           .n11575(n11575), .n11576(n11576), .n11577(n11577), .n11578(n11578), 
           .n11579(n11579), .n34843(n34843), .delay_i_23__N_1202({delay_i_23__N_1202_adj_7484}), 
           .\no5_state[0] (no5_state[0]), .op_i_23__N_1154({op_i_23__N_1154_adj_7426}), 
           .delay_r_23__N_1178({delay_r_23__N_1178_adj_7483}), .op_r_23__N_1106({op_r_23__N_1106_adj_7425}), 
           .dout_r_23__N_5926({dout_r_23__N_5926}), .s5_count(s5_count), 
           .r4_valid(r4_valid), .\op_i_23__N_1130[16] (op_i_23__N_1130_adj_7492[16]), 
           .\op_i_23__N_1154[8]_adj_1 (op_i_23__N_1154_adj_7482[8]), .\out_i[8] (out_i[8]), 
           .\op_i_23__N_1130[21] (op_i_23__N_1130_adj_7492[21]), .\op_i_23__N_1154[13]_adj_2 (op_i_23__N_1154_adj_7482[13]), 
           .\out_i[13] (out_i[13]), .\op_i_23__N_1130[20] (op_i_23__N_1130_adj_7492[20]), 
           .\op_i_23__N_1154[12]_adj_3 (op_i_23__N_1154_adj_7482[12]), .\out_i[12] (out_i[12]), 
           .\op_i_23__N_1130[19] (op_i_23__N_1130_adj_7492[19]), .\op_i_23__N_1154[11]_adj_4 (op_i_23__N_1154_adj_7482[11]), 
           .\out_i[11] (out_i[11]), .\op_i_23__N_1130[18] (op_i_23__N_1130_adj_7492[18]), 
           .\op_i_23__N_1154[10]_adj_5 (op_i_23__N_1154_adj_7482[10]), .\out_i[10] (out_i[10]), 
           .\op_i_23__N_1130[17] (op_i_23__N_1130_adj_7492[17]), .\op_i_23__N_1154[9]_adj_6 (op_i_23__N_1154_adj_7482[9]), 
           .\out_i[9] (out_i[9]), .\op_i_23__N_1130[31] (op_i_23__N_1130_adj_7492[31]), 
           .\op_i_23__N_1154[23]_adj_7 (op_i_23__N_1154_adj_7482[23]), .\out_i[23] (out_i[23]), 
           .\op_i_23__N_1130[30] (op_i_23__N_1130_adj_7492[30]), .\op_i_23__N_1154[22]_adj_8 (op_i_23__N_1154_adj_7482[22]), 
           .\out_i[22] (out_i[22]), .\op_i_23__N_1130[29] (op_i_23__N_1130_adj_7492[29]), 
           .\op_i_23__N_1154[21]_adj_9 (op_i_23__N_1154_adj_7482[21]), .\out_i[21] (out_i[21]), 
           .\op_i_23__N_1130[28] (op_i_23__N_1130_adj_7492[28]), .\op_i_23__N_1154[20]_adj_10 (op_i_23__N_1154_adj_7482[20]), 
           .\out_i[20] (out_i[20]), .\op_i_23__N_1130[27] (op_i_23__N_1130_adj_7492[27]), 
           .\op_i_23__N_1154[19]_adj_11 (op_i_23__N_1154_adj_7482[19]), .\out_i[19] (out_i[19]), 
           .\op_i_23__N_1130[26] (op_i_23__N_1130_adj_7492[26]), .\op_i_23__N_1154[18]_adj_12 (op_i_23__N_1154_adj_7482[18]), 
           .\out_i[18] (out_i[18]), .\op_i_23__N_1130[25] (op_i_23__N_1130_adj_7492[25]), 
           .\op_i_23__N_1154[17]_adj_13 (op_i_23__N_1154_adj_7482[17]), .\out_i[17] (out_i[17]), 
           .\op_i_23__N_1130[24] (op_i_23__N_1130_adj_7492[24]), .\op_i_23__N_1154[16]_adj_14 (op_i_23__N_1154_adj_7482[16]), 
           .\out_i[16] (out_i[16]), .\op_i_23__N_1130[23] (op_i_23__N_1130_adj_7492[23]), 
           .\op_i_23__N_1154[15]_adj_15 (op_i_23__N_1154_adj_7482[15]), .\out_i[15] (out_i[15]), 
           .\op_i_23__N_1130[22] (op_i_23__N_1130_adj_7492[22]), .\op_i_23__N_1154[14]_adj_16 (op_i_23__N_1154_adj_7482[14]), 
           .\out_i[14] (out_i[14]), .\op_r_23__N_1082[16] (op_r_23__N_1082_adj_7489[16]), 
           .\op_r_23__N_1106[8]_adj_17 (op_r_23__N_1106_adj_7481[8]), .\out_r[8] (out_r[8]), 
           .\op_r_23__N_1082[17] (op_r_23__N_1082_adj_7489[17]), .\op_r_23__N_1106[9]_adj_18 (op_r_23__N_1106_adj_7481[9]), 
           .\out_r[9] (out_r[9]), .\op_r_23__N_1082[18] (op_r_23__N_1082_adj_7489[18]), 
           .\op_r_23__N_1106[10]_adj_19 (op_r_23__N_1106_adj_7481[10]), .\out_r[10] (out_r[10]), 
           .\op_r_23__N_1082[19] (op_r_23__N_1082_adj_7489[19]), .\op_r_23__N_1106[11]_adj_20 (op_r_23__N_1106_adj_7481[11]), 
           .\out_r[11] (out_r[11]), .\op_r_23__N_1082[20] (op_r_23__N_1082_adj_7489[20]), 
           .\op_r_23__N_1106[12]_adj_21 (op_r_23__N_1106_adj_7481[12]), .\out_r[12] (out_r[12]), 
           .\op_r_23__N_1082[21] (op_r_23__N_1082_adj_7489[21]), .\op_r_23__N_1106[13]_adj_22 (op_r_23__N_1106_adj_7481[13]), 
           .\out_r[13] (out_r[13]), .\op_r_23__N_1082[22] (op_r_23__N_1082_adj_7489[22]), 
           .\op_r_23__N_1106[14]_adj_23 (op_r_23__N_1106_adj_7481[14]), .\out_r[14] (out_r[14]), 
           .\op_r_23__N_1082[23] (op_r_23__N_1082_adj_7489[23]), .\op_r_23__N_1106[15]_adj_24 (op_r_23__N_1106_adj_7481[15]), 
           .\out_r[15] (out_r[15]), .\op_r_23__N_1082[24] (op_r_23__N_1082_adj_7489[24]), 
           .\op_r_23__N_1106[16]_adj_25 (op_r_23__N_1106_adj_7481[16]), .\out_r[16] (out_r[16]), 
           .\op_r_23__N_1082[25] (op_r_23__N_1082_adj_7489[25]), .\op_r_23__N_1106[17]_adj_26 (op_r_23__N_1106_adj_7481[17]), 
           .\out_r[17] (out_r[17]), .\op_r_23__N_1082[26] (op_r_23__N_1082_adj_7489[26]), 
           .\op_r_23__N_1106[18]_adj_27 (op_r_23__N_1106_adj_7481[18]), .\out_r[18] (out_r[18]), 
           .\op_r_23__N_1082[27] (op_r_23__N_1082_adj_7489[27]), .\op_r_23__N_1106[19]_adj_28 (op_r_23__N_1106_adj_7481[19]), 
           .\out_r[19] (out_r[19]), .\op_r_23__N_1082[28] (op_r_23__N_1082_adj_7489[28]), 
           .\op_r_23__N_1106[20]_adj_29 (op_r_23__N_1106_adj_7481[20]), .\out_r[20] (out_r[20]), 
           .\op_r_23__N_1082[29] (op_r_23__N_1082_adj_7489[29]), .\op_r_23__N_1106[21]_adj_30 (op_r_23__N_1106_adj_7481[21]), 
           .\out_r[21] (out_r[21]), .\op_r_23__N_1082[30] (op_r_23__N_1082_adj_7489[30]), 
           .\op_r_23__N_1106[22]_adj_31 (op_r_23__N_1106_adj_7481[22]), .\out_r[22] (out_r[22]), 
           .\op_r_23__N_1082[31] (op_r_23__N_1082_adj_7489[31]), .\op_r_23__N_1106[23]_adj_32 (op_r_23__N_1106_adj_7481[23]), 
           .\out_r[23] (out_r[23])) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(217[8] 230[2])
    FD1P3AX count_y_689__i1 (.D(n34), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(count_y[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689__i1.GSR = "ENABLED";
    FD1P3AX count_y_689__i2 (.D(n33), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(count_y[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689__i2.GSR = "ENABLED";
    FD1P3AX count_y_689__i3 (.D(n32), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(count_y[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689__i3.GSR = "ENABLED";
    FD1P3AX count_y_689__i4 (.D(n31), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(count_y[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689__i4.GSR = "ENABLED";
    FD1P3AX count_y_689__i5 (.D(n30), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(count_y[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(251[43:57])
    defparam count_y_689__i5.GSR = "ENABLED";
    ROM_16 rom16 (.clk_c(clk_c), .n34737(n34737), .n30203(n30203), .\rom16_w_i[5] (rom16_w_i[5]), 
           .\count[4] (count[4]), .n30207(n30207), .n33013(n33013), .n30197(n30197), 
           .n34736(n34736), .n32928(n32928), .\count[5] (count[5]), .n34735(n34735), 
           .\rom16_w_i[1] (rom16_w_i[1]), .\rom16_w_i[6] (rom16_w_i[6]), 
           .n20089(n20089), .\rom16_w_r[1] (rom16_w_r[1]), .n28589(n28589), 
           .\rom16_w_r[2] (rom16_w_r[2]), .n20095(n20095), .\rom16_w_r[3] (rom16_w_r[3]), 
           .n20103(n20103), .\rom16_w_r[4] (rom16_w_r[4]), .n28591(n28591), 
           .\rom16_w_r[5] (rom16_w_r[5]), .\rom16_w_r[8] (rom16_w_r[8]), 
           .n17(n17), .GND_net(GND_net), .VCC_net(VCC_net), .in_valid_reg(in_valid_reg), 
           .n34713(n34713), .\rom16_w_i[8] (rom16_w_i[8]), .n34727(n34727), 
           .\rom16_w_i[0] (rom16_w_i[0]), .\rom16_w_r[6] (rom16_w_r[6]), 
           .n30499(n30499), .\rom16_w_i[2] (rom16_w_i[2]), .\rom16_w_i[3] (rom16_w_i[3]), 
           .n33030(n33030), .\rom16_w_i[4] (rom16_w_i[4]), .n34729(n34729), 
           .\rom16_w_i[7] (rom16_w_i[7]), .n34730(n34730), .n34789(n34789), 
           .\rom16_w_r[9] (rom16_w_r[9]), .n33051(n33051), .n28598(n28598), 
           .\rom16_w_r[0] (rom16_w_r[0]), .n34757(n34757), .n34733(n34733), 
           .\op_i_23__N_1130[17] (op_i_23__N_1130[17]), .\din_i_reg[9] (din_i_reg[9]), 
           .n31698(n31698), .\op_i_23__N_1130[16] (op_i_23__N_1130[16]), 
           .\din_i_reg[8] (din_i_reg[8]), .n31700(n31700), .\op_i_23__N_1130[19] (op_i_23__N_1130[19]), 
           .\din_i_reg[11] (din_i_reg[11]), .n31694(n31694), .\op_i_23__N_1130[18] (op_i_23__N_1130[18]), 
           .\din_i_reg[10] (din_i_reg[10]), .n31696(n31696), .\op_i_23__N_1130[21] (op_i_23__N_1130[21]), 
           .\din_i_reg[13] (din_i_reg[13]), .n31690(n31690), .\op_i_23__N_1130[20] (op_i_23__N_1130[20]), 
           .\din_i_reg[12] (din_i_reg[12]), .n31692(n31692), .\op_i_23__N_1130[23] (op_i_23__N_1130[23]), 
           .\din_i_reg[15] (din_i_reg[15]), .n31686(n31686), .\op_i_23__N_1130[22] (op_i_23__N_1130[22]), 
           .\din_i_reg[14] (din_i_reg[14]), .n31688(n31688), .\op_i_23__N_1130[25] (op_i_23__N_1130[25]), 
           .\din_i_reg[17] (din_i_reg[17]), .n31682(n31682), .\op_i_23__N_1130[24] (op_i_23__N_1130[24]), 
           .\din_i_reg[16] (din_i_reg[16]), .n31684(n31684), .\op_i_23__N_1130[27] (op_i_23__N_1130[27]), 
           .\din_i_reg[23] (din_i_reg[23]), .n31678(n31678), .\op_i_23__N_1130[26] (op_i_23__N_1130[26]), 
           .\din_i_reg[18] (din_i_reg[18]), .n31680(n31680), .\op_i_23__N_1130[29] (op_i_23__N_1130[29]), 
           .n31674(n31674), .\op_i_23__N_1130[28] (op_i_23__N_1130[28]), 
           .n31676(n31676), .\op_i_23__N_1130[31] (op_i_23__N_1130[31]), 
           .n31670(n31670), .\op_i_23__N_1130[30] (op_i_23__N_1130[30]), 
           .n31672(n31672), .\op_r_23__N_1082[17] (op_r_23__N_1082[17]), 
           .\din_r_reg[9] (din_r_reg[9]), .n31731(n31731), .\op_r_23__N_1082[16] (op_r_23__N_1082[16]), 
           .\din_r_reg[8] (din_r_reg[8]), .n31733(n31733), .\rom16_w_r[7] (rom16_w_r[7]), 
           .\op_r_23__N_1082[30] (op_r_23__N_1082[30]), .\din_r_reg[23] (din_r_reg[23]), 
           .n31705(n31705), .\op_r_23__N_1082[31] (op_r_23__N_1082[31]), 
           .n31703(n31703), .\op_r_23__N_1082[28] (op_r_23__N_1082[28]), 
           .n31709(n31709), .\op_r_23__N_1082[29] (op_r_23__N_1082[29]), 
           .n31707(n31707), .\op_r_23__N_1082[26] (op_r_23__N_1082[26]), 
           .\din_r_reg[18] (din_r_reg[18]), .n31713(n31713), .\op_r_23__N_1082[27] (op_r_23__N_1082[27]), 
           .n31711(n31711), .\op_r_23__N_1082[24] (op_r_23__N_1082[24]), 
           .\din_r_reg[16] (din_r_reg[16]), .n31717(n31717), .\op_r_23__N_1082[25] (op_r_23__N_1082[25]), 
           .\din_r_reg[17] (din_r_reg[17]), .n31715(n31715), .\op_r_23__N_1082[22] (op_r_23__N_1082[22]), 
           .\din_r_reg[14] (din_r_reg[14]), .n31721(n31721), .\op_r_23__N_1082[23] (op_r_23__N_1082[23]), 
           .\din_r_reg[15] (din_r_reg[15]), .n31719(n31719), .\op_r_23__N_1082[20] (op_r_23__N_1082[20]), 
           .\din_r_reg[12] (din_r_reg[12]), .n31725(n31725), .\op_r_23__N_1082[21] (op_r_23__N_1082[21]), 
           .\din_r_reg[13] (din_r_reg[13]), .n31723(n31723), .\op_r_23__N_1082[18] (op_r_23__N_1082[18]), 
           .\din_r_reg[10] (din_r_reg[10]), .n31729(n31729), .\op_r_23__N_1082[19] (op_r_23__N_1082[19]), 
           .\din_r_reg[11] (din_r_reg[11]), .n31727(n31727), .n34759(n34759)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(106[8] 113[2])
    shift_16 shift_16 (.clk_c(clk_c), .in_valid_reg(in_valid_reg), .VCC_net(VCC_net), 
            .\op_i_23__N_1154[7] (op_i_23__N_1154[7]), .\op_i_23__N_1154[6] (op_i_23__N_1154[6]), 
            .\op_i_23__N_1154[5] (op_i_23__N_1154[5]), .\op_i_23__N_1154[4] (op_i_23__N_1154[4]), 
            .\op_i_23__N_1154[3] (op_i_23__N_1154[3]), .\op_i_23__N_1154[2] (op_i_23__N_1154[2]), 
            .\op_i_23__N_1154[1] (op_i_23__N_1154[1]), .\op_r_23__N_1106[7] (op_r_23__N_1106[7]), 
            .\op_r_23__N_1106[6] (op_r_23__N_1106[6]), .\op_r_23__N_1106[5] (op_r_23__N_1106[5]), 
            .\op_r_23__N_1106[4] (op_r_23__N_1106[4]), .\op_r_23__N_1106[3] (op_r_23__N_1106[3]), 
            .\op_r_23__N_1106[2] (op_r_23__N_1106[2]), .\op_r_23__N_1106[1] (op_r_23__N_1106[1]), 
            .\op_i_23__N_1154[0] (op_i_23__N_1154[0]), .\op_r_23__N_1106[0] (op_r_23__N_1106[0]), 
            .\dout_r_23__N_2506[8] (dout_r_23__N_2506[8]), .\dout_r_23__N_2506[9] (dout_r_23__N_2506[9]), 
            .\dout_r_23__N_2506[10] (dout_r_23__N_2506[10]), .\dout_r_23__N_2506[11] (dout_r_23__N_2506[11]), 
            .\dout_r_23__N_2506[12] (dout_r_23__N_2506[12]), .\dout_r_23__N_2506[13] (dout_r_23__N_2506[13]), 
            .\dout_r_23__N_2506[14] (dout_r_23__N_2506[14]), .\dout_r_23__N_2506[15] (dout_r_23__N_2506[15]), 
            .\dout_r_23__N_2506[16] (dout_r_23__N_2506[16]), .\dout_r_23__N_2506[17] (dout_r_23__N_2506[17]), 
            .\dout_r_23__N_2506[18] (dout_r_23__N_2506[18]), .\dout_r_23__N_2506[19] (dout_r_23__N_2506[19]), 
            .\dout_r_23__N_2506[20] (dout_r_23__N_2506[20]), .\dout_r_23__N_2506[21] (dout_r_23__N_2506[21]), 
            .\dout_r_23__N_2506[22] (dout_r_23__N_2506[22]), .\dout_r_23__N_2506[23] (dout_r_23__N_2506[23]), 
            .\shift_16_dout_i[23] (shift_16_dout_i[23]), .\shift_16_dout_i[22] (shift_16_dout_i[22]), 
            .\shift_16_dout_i[21] (shift_16_dout_i[21]), .\shift_16_dout_i[20] (shift_16_dout_i[20]), 
            .\shift_16_dout_i[19] (shift_16_dout_i[19]), .\shift_16_dout_i[18] (shift_16_dout_i[18]), 
            .\shift_16_dout_i[17] (shift_16_dout_i[17]), .\shift_16_dout_i[16] (shift_16_dout_i[16]), 
            .\shift_16_dout_i[15] (shift_16_dout_i[15]), .\shift_16_dout_i[14] (shift_16_dout_i[14]), 
            .\shift_16_dout_i[13] (shift_16_dout_i[13]), .\shift_16_dout_i[12] (shift_16_dout_i[12]), 
            .\shift_16_dout_i[11] (shift_16_dout_i[11]), .\shift_16_dout_i[10] (shift_16_dout_i[10]), 
            .\shift_16_dout_i[9] (shift_16_dout_i[9]), .\shift_16_dout_i[8] (shift_16_dout_i[8]), 
            .\shift_16_dout_r[23] (shift_16_dout_r[23]), .\shift_16_dout_r[22] (shift_16_dout_r[22]), 
            .\shift_16_dout_r[21] (shift_16_dout_r[21]), .\shift_16_dout_r[20] (shift_16_dout_r[20]), 
            .\shift_16_dout_r[19] (shift_16_dout_r[19]), .\shift_16_dout_r[18] (shift_16_dout_r[18]), 
            .\shift_16_dout_r[17] (shift_16_dout_r[17]), .\shift_16_dout_r[16] (shift_16_dout_r[16]), 
            .\shift_16_dout_r[15] (shift_16_dout_r[15]), .\shift_16_dout_r[13] (shift_16_dout_r[13]), 
            .\shift_16_dout_r[12] (shift_16_dout_r[12]), .\shift_16_dout_r[11] (shift_16_dout_r[11]), 
            .\shift_16_dout_r[10] (shift_16_dout_r[10]), .\shift_16_dout_r[9] (shift_16_dout_r[9]), 
            .\shift_16_dout_r[8] (shift_16_dout_r[8]), .\shift_16_dout_r[14] (shift_16_dout_r[14]), 
            .\count[5] (count[5]), .\count[4] (count[4]), .\dout_i_23__N_3274[8] (dout_i_23__N_3274[8]), 
            .\dout_i_23__N_3274[9] (dout_i_23__N_3274[9]), .\dout_i_23__N_3274[10] (dout_i_23__N_3274[10]), 
            .\dout_i_23__N_3274[11] (dout_i_23__N_3274[11]), .\dout_i_23__N_3274[12] (dout_i_23__N_3274[12]), 
            .\dout_i_23__N_3274[13] (dout_i_23__N_3274[13]), .\dout_i_23__N_3274[14] (dout_i_23__N_3274[14]), 
            .\dout_i_23__N_3274[15] (dout_i_23__N_3274[15]), .\dout_i_23__N_3274[16] (dout_i_23__N_3274[16]), 
            .\dout_i_23__N_3274[17] (dout_i_23__N_3274[17]), .\dout_i_23__N_3274[18] (dout_i_23__N_3274[18]), 
            .\dout_i_23__N_3274[19] (dout_i_23__N_3274[19]), .\dout_i_23__N_3274[20] (dout_i_23__N_3274[20]), 
            .\dout_i_23__N_3274[21] (dout_i_23__N_3274[21]), .\dout_i_23__N_3274[22] (dout_i_23__N_3274[22]), 
            .\dout_i_23__N_3274[23] (dout_i_23__N_3274[23])) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(97[10] 104[2])
    ROM_2 rom2 (.clk_c(clk_c), .clk_c_enable_2299(clk_c_enable_2299), .clk_c_enable_2300(clk_c_enable_2300), 
          .n34839(n34839), .n34801(n34801), .n34843(n34843), .\s_count[1] (s_count_adj_7458[1]), 
          .GND_net(GND_net), .VCC_net(VCC_net), .\count[1] (count_adj_7456[1]), 
          .n34800(n34800), .\state_1__N_5843[1] (state_1__N_5843[1]), .n30179(n30179), 
          .valid(valid_adj_7215), .n34738(n34738), .n34795(n34795), .\rom2_w_r[8] (rom2_w_r[8]), 
          .n34769(n34769)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(207[7] 214[2])
    shift_1 shift_1 (.rst_n_c(rst_n_c), .rst_n_N_2(rst_n_N_2), .valid(valid_adj_7215), 
            .clk_c(clk_c), .n34738(n34738), .n34843(n34843), .dout_i_23__N_5974({dout_i_23__N_5974}), 
            .shift_1_dout_i({shift_1_dout_i}), .dout_r_23__N_5926({dout_r_23__N_5926}), 
            .shift_1_dout_r({shift_1_dout_r})) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(232[9] 239[2])
    ROM_4 rom4 (.n29820(n29820), .n29819(n29819), .n34520(n34520), .\rom4_state[0] (rom4_state[0]), 
          .state_1__N_5502(state_1__N_5502), .clk_c(clk_c), .clk_c_enable_2305(clk_c_enable_2305), 
          .s_count({s_count_adj_7402}), .\rom4_w_i[12] (rom4_w_i[12]), .GND_net(GND_net), 
          .VCC_net(VCC_net), .n29826(n29826), .n29828(n29828), .n29827(n29827), 
          .n34841(n34841), .\rom4_w_r[1] (rom4_w_r[1]), .n34776(n34776), 
          .\rom4_w_r[8] (rom4_w_r[8]), .n34777(n34777), .\rom4_w_r[5] (rom4_w_r[5]), 
          .n34799(n34799), .clk_c_enable_2299(clk_c_enable_2299), .n6514(n6514), 
          .n3(n3), .n30041(n30041)) /* synthesis syn_module_defined=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(173[7] 180[2])
    
endmodule
//
// Verilog Description of module radix2_U2
//

module radix2_U2 (op_r_23__N_1106, n34842, n3, shift_4_dout_r, n7431, 
            n6514, \op_r_23__N_1082[29] , n31429, op_i_23__N_1154, shift_4_dout_i, 
            n7590, \op_i_23__N_1130[26] , n31484, GND_net, \op_i_23__N_1310[0] , 
            \op_i_23__N_1310[1] , \op_i_23__N_1310[2] , \op_i_23__N_1310[3] , 
            \op_i_23__N_1310[4] , \op_i_23__N_1310[5] , n89, n88, n87, 
            n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, 
            n76, n75, n74, n73, n72, n71, n70, n69, n68, n67, 
            n66, n65, VCC_net, \rom8_w_i[12] , n11148, n11149, n11150, 
            n11151, n11152, n11153, \op_i_23__N_1130[27] , n31482, 
            \rom8_w_i[0] , \rom8_w_i[1] , \rom8_w_i[2] , \rom8_w_i[3] , 
            \rom8_w_i[4] , \rom8_w_i[6] , \op_r_23__N_1082[26] , n31435, 
            \op_r_23__N_1082[27] , n31433, shift_8_dout_i, n119, \op_r_23__N_1268[0] , 
            \op_r_23__N_1268[1] , \op_r_23__N_1268[2] , \op_r_23__N_1268[3] , 
            \op_r_23__N_1268[4] , \op_r_23__N_1268[5] , \op_r_23__N_1268[6] , 
            \op_r_23__N_1268[7] , \op_r_23__N_1268[8] , \op_r_23__N_1268[9] , 
            \op_r_23__N_1268[10] , \op_r_23__N_1268[11] , \op_r_23__N_1268[12] , 
            \op_r_23__N_1268[13] , \op_r_23__N_1268[14] , \op_r_23__N_1268[15] , 
            \op_r_23__N_1268[16] , \op_r_23__N_1268[17] , \op_r_23__N_1268[18] , 
            \op_r_23__N_1268[19] , \op_r_23__N_1268[20] , \op_r_23__N_1268[21] , 
            \op_r_23__N_1268[22] , \op_r_23__N_1268[23] , \op_r_23__N_1268[24] , 
            \op_r_23__N_1268[25] , \op_r_23__N_1268[26] , \op_r_23__N_1268[27] , 
            \op_r_23__N_1268[28] , \op_r_23__N_1268[29] , \op_r_23__N_1268[30] , 
            \op_r_23__N_1268[31] , \op_r_23__N_1226[0] , \op_r_23__N_1226[1] , 
            \op_r_23__N_1226[2] , \op_r_23__N_1226[3] , \op_r_23__N_1226[4] , 
            \op_r_23__N_1226[5] , \op_r_23__N_1226[6] , \op_r_23__N_1226[7] , 
            \op_r_23__N_1226[8] , \op_r_23__N_1226[9] , \op_r_23__N_1226[10] , 
            \op_r_23__N_1226[11] , \op_r_23__N_1226[12] , \op_r_23__N_1226[13] , 
            \op_r_23__N_1226[14] , \op_r_23__N_1226[15] , \op_r_23__N_1226[16] , 
            \op_r_23__N_1226[17] , \op_r_23__N_1226[18] , \op_r_23__N_1226[19] , 
            \op_r_23__N_1226[20] , \op_r_23__N_1226[21] , \op_r_23__N_1226[22] , 
            \op_r_23__N_1226[23] , \op_r_23__N_1226[24] , \op_r_23__N_1226[25] , 
            \op_r_23__N_1226[26] , \op_r_23__N_1226[27] , \op_r_23__N_1226[28] , 
            \op_r_23__N_1226[29] , \op_r_23__N_1226[30] , \op_r_23__N_1226[31] , 
            \op_i_23__N_1130[24] , n31488, \rom8_w_r[0] , \rom8_w_r[1] , 
            \rom8_w_r[7] , \rom8_w_r[3] , \rom8_w_r[4] , \rom8_w_r[5] , 
            \rom8_w_r[6] , \rom8_w_r[8] , \rom8_w_r[10] , n12270, n12271, 
            n12272, n12273, n12274, n12275, n12276, n12277, n12278, 
            n12279, n12280, n12281, n12282, n12283, n12284, n12285, 
            n12286, n12287, n8721, n8720, n8719, n8718, n8717, 
            n8716, n8715, n8714, n8713, n8712, n8711, n8710, n8709, 
            n8708, n8707, n8706, n8705, n8704, n8703, n8702, n8701, 
            n8700, n8699, n8698, n8697, n8696, n319, n11154, n11155, 
            n11156, n11157, n11158, n11159, n11160, n11161, n11162, 
            n11163, n11164, n11165, n11166, n11167, n11168, n11169, 
            n11170, n11171, n12444, n12445, n12446, n12447, n12448, 
            n12449, n12450, n12451, n12452, n12453, n12288, n12289, 
            n12290, n12291, n12292, n12293, n12294, \op_i_23__N_1130[25] , 
            n31486, \op_r_23__N_1082[24] , n31439, \op_r_23__N_1082[25] , 
            n31437, \op_i_23__N_1130[22] , n31492, \op_i_23__N_1130[23] , 
            n31490, \op_r_23__N_1082[22] , n31443, \op_r_23__N_1082[23] , 
            n31441, \op_i_23__N_1130[20] , n31496, \op_i_23__N_1130[21] , 
            n31494, \op_r_23__N_1082[20] , n31447, \op_r_23__N_1082[21] , 
            n31445, \op_i_23__N_1130[18] , n31500, \op_i_23__N_1130[19] , 
            n31498, \op_r_23__N_1082[18] , n31451, \op_r_23__N_1082[19] , 
            n31449, \op_i_23__N_1130[16] , n31504, \op_i_23__N_1130[17] , 
            n31502, \op_i_23__N_1130[31] , n31474, \op_r_23__N_1082[16] , 
            n31455, \op_r_23__N_1082[17] , n31453, \op_r_23__N_1082[30] , 
            n31427, \op_i_23__N_1130[30] , n31476, \op_r_23__N_1082[31] , 
            n31425, \rom8_state[0] , n34794, \radix_no1_op_i[1] , n7507, 
            \radix_no1_op_i[0] , n7508, \radix_no1_op_i[3] , n7505, 
            \radix_no1_op_i[2] , n7506, \radix_no1_op_i[5] , n7503, 
            \radix_no1_op_i[4] , n7504, \radix_no1_op_i[7] , n7501, 
            \radix_no1_op_i[6] , n7502, \radix_no1_op_r[1] , \shift_8_dout_r[1] , 
            n7560, \radix_no1_op_r[0] , \shift_8_dout_r[0] , n7561, 
            \radix_no1_op_r[3] , \shift_8_dout_r[3] , n7558, \radix_no1_op_r[2] , 
            \shift_8_dout_r[2] , n7559, \radix_no1_op_r[5] , \shift_8_dout_r[5] , 
            n7556, \radix_no1_op_r[4] , \shift_8_dout_r[4] , n7557, 
            \radix_no1_op_r[7] , \shift_8_dout_r[7] , n7554, \radix_no1_op_r[6] , 
            \shift_8_dout_r[6] , n7555, \op_i_23__N_1130[8] , n31422, 
            \op_i_23__N_1130[9] , n31420, \op_i_23__N_1130[13] , n31412, 
            \op_i_23__N_1130[10] , n31418, \op_i_23__N_1130[11] , n31416, 
            \op_i_23__N_1130[14] , n31410, \op_i_23__N_1130[15] , n31408, 
            \op_i_23__N_1130[12] , n31414, \op_r_23__N_1082[14] , n31606, 
            \op_r_23__N_1082[15] , n31604, \op_r_23__N_1082[12] , n31610, 
            \op_r_23__N_1082[13] , n31608, \op_r_23__N_1082[10] , n31614, 
            \op_r_23__N_1082[11] , n31612, \op_r_23__N_1082[8] , n31618, 
            \op_r_23__N_1082[9] , n31616, n34625, n34620, n34619, 
            n34614, n34613, n34608, n34607, n34606, n34605, n34600, 
            n34599, n34598, n34597, n34592, n34591, n34590, n34589, 
            n34626, n34631, n34632, n34637, n34638, n34643, n34644, 
            n34647, n34648, n34653, n34654, n34657, n34658, n34663, 
            n34664, n34681, n34682, n34687, n34688, n34691, n34692, 
            n34693, n34694, n34695, n34696, n34697, n34698, n34699, 
            n34700, n34701, n34702, valid, clk_c_enable_1373, \op_i_23__N_1130[14]_adj_70 , 
            n31508, \op_i_23__N_1130[15]_adj_71 , n31506, \op_r_23__N_1082[14]_adj_72 , 
            n31459, \op_r_23__N_1082[15]_adj_73 , n31457, \op_i_23__N_1130[13]_adj_74 , 
            n31510, \op_r_23__N_1082[12]_adj_75 , n31463, \op_r_23__N_1082[13]_adj_76 , 
            n31461, \op_i_23__N_1130[12]_adj_77 , n31512, \op_r_23__N_1082[28] , 
            n31431, \op_r_23__N_1082[10]_adj_78 , n31467, \op_r_23__N_1082[11]_adj_79 , 
            n31465, \op_i_23__N_1130[10]_adj_80 , n31516, \op_i_23__N_1130[11]_adj_81 , 
            n31514, \op_r_23__N_1082[8]_adj_82 , n31471, \op_r_23__N_1082[9]_adj_83 , 
            n31469, \op_i_23__N_1130[8]_adj_84 , n31520, \op_i_23__N_1130[9]_adj_85 , 
            n31518, \op_i_23__N_1130[29] , n31478, \op_i_23__N_1130[28] , 
            n31480) /* synthesis syn_module_defined=1 */ ;
    input [23:0]op_r_23__N_1106;
    input n34842;
    input n3;
    input [23:0]shift_4_dout_r;
    output [23:0]n7431;
    input n6514;
    input \op_r_23__N_1082[29] ;
    output n31429;
    input [23:0]op_i_23__N_1154;
    input [23:0]shift_4_dout_i;
    output [23:0]n7590;
    input \op_i_23__N_1130[26] ;
    output n31484;
    input GND_net;
    output \op_i_23__N_1310[0] ;
    output \op_i_23__N_1310[1] ;
    output \op_i_23__N_1310[2] ;
    output \op_i_23__N_1310[3] ;
    output \op_i_23__N_1310[4] ;
    output \op_i_23__N_1310[5] ;
    output n89;
    output n88;
    output n87;
    output n86;
    output n85;
    output n84;
    output n83;
    output n82;
    output n81;
    output n80;
    output n79;
    output n78;
    output n77;
    output n76;
    output n75;
    output n74;
    output n73;
    output n72;
    output n71;
    output n70;
    output n69;
    output n68;
    output n67;
    output n66;
    output n65;
    input VCC_net;
    input \rom8_w_i[12] ;
    input n11148;
    input n11149;
    input n11150;
    input n11151;
    input n11152;
    input n11153;
    input \op_i_23__N_1130[27] ;
    output n31482;
    input \rom8_w_i[0] ;
    input \rom8_w_i[1] ;
    input \rom8_w_i[2] ;
    input \rom8_w_i[3] ;
    input \rom8_w_i[4] ;
    input \rom8_w_i[6] ;
    input \op_r_23__N_1082[26] ;
    output n31435;
    input \op_r_23__N_1082[27] ;
    output n31433;
    input [23:0]shift_8_dout_i;
    input n119;
    output \op_r_23__N_1268[0] ;
    output \op_r_23__N_1268[1] ;
    output \op_r_23__N_1268[2] ;
    output \op_r_23__N_1268[3] ;
    output \op_r_23__N_1268[4] ;
    output \op_r_23__N_1268[5] ;
    output \op_r_23__N_1268[6] ;
    output \op_r_23__N_1268[7] ;
    output \op_r_23__N_1268[8] ;
    output \op_r_23__N_1268[9] ;
    output \op_r_23__N_1268[10] ;
    output \op_r_23__N_1268[11] ;
    output \op_r_23__N_1268[12] ;
    output \op_r_23__N_1268[13] ;
    output \op_r_23__N_1268[14] ;
    output \op_r_23__N_1268[15] ;
    output \op_r_23__N_1268[16] ;
    output \op_r_23__N_1268[17] ;
    output \op_r_23__N_1268[18] ;
    output \op_r_23__N_1268[19] ;
    output \op_r_23__N_1268[20] ;
    output \op_r_23__N_1268[21] ;
    output \op_r_23__N_1268[22] ;
    output \op_r_23__N_1268[23] ;
    output \op_r_23__N_1268[24] ;
    output \op_r_23__N_1268[25] ;
    output \op_r_23__N_1268[26] ;
    output \op_r_23__N_1268[27] ;
    output \op_r_23__N_1268[28] ;
    output \op_r_23__N_1268[29] ;
    output \op_r_23__N_1268[30] ;
    output \op_r_23__N_1268[31] ;
    output \op_r_23__N_1226[0] ;
    output \op_r_23__N_1226[1] ;
    output \op_r_23__N_1226[2] ;
    output \op_r_23__N_1226[3] ;
    output \op_r_23__N_1226[4] ;
    output \op_r_23__N_1226[5] ;
    output \op_r_23__N_1226[6] ;
    output \op_r_23__N_1226[7] ;
    output \op_r_23__N_1226[8] ;
    output \op_r_23__N_1226[9] ;
    output \op_r_23__N_1226[10] ;
    output \op_r_23__N_1226[11] ;
    output \op_r_23__N_1226[12] ;
    output \op_r_23__N_1226[13] ;
    output \op_r_23__N_1226[14] ;
    output \op_r_23__N_1226[15] ;
    output \op_r_23__N_1226[16] ;
    output \op_r_23__N_1226[17] ;
    output \op_r_23__N_1226[18] ;
    output \op_r_23__N_1226[19] ;
    output \op_r_23__N_1226[20] ;
    output \op_r_23__N_1226[21] ;
    output \op_r_23__N_1226[22] ;
    output \op_r_23__N_1226[23] ;
    output \op_r_23__N_1226[24] ;
    output \op_r_23__N_1226[25] ;
    output \op_r_23__N_1226[26] ;
    output \op_r_23__N_1226[27] ;
    output \op_r_23__N_1226[28] ;
    output \op_r_23__N_1226[29] ;
    output \op_r_23__N_1226[30] ;
    output \op_r_23__N_1226[31] ;
    input \op_i_23__N_1130[24] ;
    output n31488;
    input \rom8_w_r[0] ;
    input \rom8_w_r[1] ;
    input \rom8_w_r[7] ;
    input \rom8_w_r[3] ;
    input \rom8_w_r[4] ;
    input \rom8_w_r[5] ;
    input \rom8_w_r[6] ;
    input \rom8_w_r[8] ;
    input \rom8_w_r[10] ;
    input n12270;
    input n12271;
    input n12272;
    input n12273;
    input n12274;
    input n12275;
    input n12276;
    input n12277;
    input n12278;
    input n12279;
    input n12280;
    input n12281;
    input n12282;
    input n12283;
    input n12284;
    input n12285;
    input n12286;
    input n12287;
    output n8721;
    output n8720;
    output n8719;
    output n8718;
    output n8717;
    output n8716;
    output n8715;
    output n8714;
    output n8713;
    output n8712;
    output n8711;
    output n8710;
    output n8709;
    output n8708;
    output n8707;
    output n8706;
    output n8705;
    output n8704;
    output n8703;
    output n8702;
    output n8701;
    output n8700;
    output n8699;
    output n8698;
    output n8697;
    output n8696;
    input n319;
    input n11154;
    input n11155;
    input n11156;
    input n11157;
    input n11158;
    input n11159;
    input n11160;
    input n11161;
    input n11162;
    input n11163;
    input n11164;
    input n11165;
    input n11166;
    input n11167;
    input n11168;
    input n11169;
    input n11170;
    input n11171;
    input n12444;
    input n12445;
    input n12446;
    input n12447;
    input n12448;
    input n12449;
    input n12450;
    input n12451;
    input n12452;
    input n12453;
    input n12288;
    input n12289;
    input n12290;
    input n12291;
    input n12292;
    input n12293;
    input n12294;
    input \op_i_23__N_1130[25] ;
    output n31486;
    input \op_r_23__N_1082[24] ;
    output n31439;
    input \op_r_23__N_1082[25] ;
    output n31437;
    input \op_i_23__N_1130[22] ;
    output n31492;
    input \op_i_23__N_1130[23] ;
    output n31490;
    input \op_r_23__N_1082[22] ;
    output n31443;
    input \op_r_23__N_1082[23] ;
    output n31441;
    input \op_i_23__N_1130[20] ;
    output n31496;
    input \op_i_23__N_1130[21] ;
    output n31494;
    input \op_r_23__N_1082[20] ;
    output n31447;
    input \op_r_23__N_1082[21] ;
    output n31445;
    input \op_i_23__N_1130[18] ;
    output n31500;
    input \op_i_23__N_1130[19] ;
    output n31498;
    input \op_r_23__N_1082[18] ;
    output n31451;
    input \op_r_23__N_1082[19] ;
    output n31449;
    input \op_i_23__N_1130[16] ;
    output n31504;
    input \op_i_23__N_1130[17] ;
    output n31502;
    input \op_i_23__N_1130[31] ;
    output n31474;
    input \op_r_23__N_1082[16] ;
    output n31455;
    input \op_r_23__N_1082[17] ;
    output n31453;
    input \op_r_23__N_1082[30] ;
    output n31427;
    input \op_i_23__N_1130[30] ;
    output n31476;
    input \op_r_23__N_1082[31] ;
    output n31425;
    input \rom8_state[0] ;
    input n34794;
    input \radix_no1_op_i[1] ;
    output n7507;
    input \radix_no1_op_i[0] ;
    output n7508;
    input \radix_no1_op_i[3] ;
    output n7505;
    input \radix_no1_op_i[2] ;
    output n7506;
    input \radix_no1_op_i[5] ;
    output n7503;
    input \radix_no1_op_i[4] ;
    output n7504;
    input \radix_no1_op_i[7] ;
    output n7501;
    input \radix_no1_op_i[6] ;
    output n7502;
    input \radix_no1_op_r[1] ;
    input \shift_8_dout_r[1] ;
    output n7560;
    input \radix_no1_op_r[0] ;
    input \shift_8_dout_r[0] ;
    output n7561;
    input \radix_no1_op_r[3] ;
    input \shift_8_dout_r[3] ;
    output n7558;
    input \radix_no1_op_r[2] ;
    input \shift_8_dout_r[2] ;
    output n7559;
    input \radix_no1_op_r[5] ;
    input \shift_8_dout_r[5] ;
    output n7556;
    input \radix_no1_op_r[4] ;
    input \shift_8_dout_r[4] ;
    output n7557;
    input \radix_no1_op_r[7] ;
    input \shift_8_dout_r[7] ;
    output n7554;
    input \radix_no1_op_r[6] ;
    input \shift_8_dout_r[6] ;
    output n7555;
    input \op_i_23__N_1130[8] ;
    output n31422;
    input \op_i_23__N_1130[9] ;
    output n31420;
    input \op_i_23__N_1130[13] ;
    output n31412;
    input \op_i_23__N_1130[10] ;
    output n31418;
    input \op_i_23__N_1130[11] ;
    output n31416;
    input \op_i_23__N_1130[14] ;
    output n31410;
    input \op_i_23__N_1130[15] ;
    output n31408;
    input \op_i_23__N_1130[12] ;
    output n31414;
    input \op_r_23__N_1082[14] ;
    output n31606;
    input \op_r_23__N_1082[15] ;
    output n31604;
    input \op_r_23__N_1082[12] ;
    output n31610;
    input \op_r_23__N_1082[13] ;
    output n31608;
    input \op_r_23__N_1082[10] ;
    output n31614;
    input \op_r_23__N_1082[11] ;
    output n31612;
    input \op_r_23__N_1082[8] ;
    output n31618;
    input \op_r_23__N_1082[9] ;
    output n31616;
    output n34625;
    output n34620;
    output n34619;
    output n34614;
    output n34613;
    output n34608;
    output n34607;
    output n34606;
    output n34605;
    output n34600;
    output n34599;
    output n34598;
    output n34597;
    output n34592;
    output n34591;
    output n34590;
    output n34589;
    output n34626;
    output n34631;
    output n34632;
    output n34637;
    output n34638;
    output n34643;
    output n34644;
    output n34647;
    output n34648;
    output n34653;
    output n34654;
    output n34657;
    output n34658;
    output n34663;
    output n34664;
    output n34681;
    output n34682;
    output n34687;
    output n34688;
    output n34691;
    output n34692;
    output n34693;
    output n34694;
    output n34695;
    output n34696;
    output n34697;
    output n34698;
    output n34699;
    output n34700;
    output n34701;
    output n34702;
    input valid;
    output clk_c_enable_1373;
    input \op_i_23__N_1130[14]_adj_70 ;
    output n31508;
    input \op_i_23__N_1130[15]_adj_71 ;
    output n31506;
    input \op_r_23__N_1082[14]_adj_72 ;
    output n31459;
    input \op_r_23__N_1082[15]_adj_73 ;
    output n31457;
    input \op_i_23__N_1130[13]_adj_74 ;
    output n31510;
    input \op_r_23__N_1082[12]_adj_75 ;
    output n31463;
    input \op_r_23__N_1082[13]_adj_76 ;
    output n31461;
    input \op_i_23__N_1130[12]_adj_77 ;
    output n31512;
    input \op_r_23__N_1082[28] ;
    output n31431;
    input \op_r_23__N_1082[10]_adj_78 ;
    output n31467;
    input \op_r_23__N_1082[11]_adj_79 ;
    output n31465;
    input \op_i_23__N_1130[10]_adj_80 ;
    output n31516;
    input \op_i_23__N_1130[11]_adj_81 ;
    output n31514;
    input \op_r_23__N_1082[8]_adj_82 ;
    output n31471;
    input \op_r_23__N_1082[9]_adj_83 ;
    output n31469;
    input \op_i_23__N_1130[8]_adj_84 ;
    output n31520;
    input \op_i_23__N_1130[9]_adj_85 ;
    output n31518;
    input \op_i_23__N_1130[29] ;
    output n31478;
    input \op_i_23__N_1130[28] ;
    output n31480;
    
    
    wire n18419, n18420, n18421, n18422, n18423, n18424, n18425, 
        n18426, n18427, n18428, n18429, n18430, n18431, n18432, 
        n18433, n18434, n18435, n18436, n18437, n18438, n18439, 
        n18440, n18441, n18442, n18443, n18444, n18445, n18446, 
        n18447, n18448, n18449, n18450, n18451, n18452, n18453, 
        n18454, n18455, n18456, n18457, n18458, n18459, n18460, 
        n18461, n18462, n18463, n18464, n18465, n18466, n18467, 
        n18468, n18469, n18470, n18471, n18472, n18473, n18474, 
        n18475, n18476, n18477, n18478, n18479, n18480, n18481, 
        n18482, n18483, n18484, n18485, n18486, n18487, n18488, 
        n18489, n18490, n18491, n18492, n18493, n18494, n18495, 
        n18496, n18497, n18498, n18499, n18500, n18501, n18502, 
        n18503, n18504, n18505, n18506, n18507, n18508, n18509, 
        n18510, n18511, n18512, n18513, n18514, n18515, n18516, 
        n18517, n18518, n18519, n18520, n18521, n18522, n18523, 
        n18524, n18525, n18526, n18527, n18528, n18529, n18530, 
        n18531, n18532, n18533, n18534, n18535, n18536, n18537, 
        n18538, n18539, n18540, n18541, n18542, n18543, n18544, 
        n18545, n18546, n18547, n18548, n18549, n18550, n18551, 
        n18552, n18553, n18554, n18555, n18556, n18557, n18558, 
        n18559, n18560, n18561, n18562, n18563, n18564, n17544, 
        n17545, n17546, n17547, n17548, n17549, n17550, n17551, 
        n17552, n17553, n17554, n17555, n17556, n17557, n17558, 
        n17559, n17560, n17561, n17562, n17563, n17564, n17565, 
        n17566, n17567, n17568, n17569, n17570, n17571, n17572, 
        n17573, n17574, n17575, n17576, n17577, n17578, n17579, 
        n17580, n17581, n17582, n17583, n17584, n17585, n17586, 
        n17587, n17588, n17589, n17590, n17591, n17592, n17593, 
        n17594, n17595, n17596, n17597, n17598, n17599, n17600, 
        n17601, n17602, n17603, n17604, n17605, n17606, n17607, 
        n17608, n17609, n17610, n17611, n17612, n17613, n17614, 
        n17615, n17616, n17617, n17618, n17619, n17620, n17621, 
        n17622, n17623, n17624, n17625, n17626, n17627, n17628, 
        n17629, n17630, n17631, n17632, n17633, n17634, n17635, 
        n17636, n17637, n17638, n17639, n17640, n17641, n17642, 
        n17643, n17644, n17645, n17646, n17647, n17648, n17649, 
        n17650, n17651, n17652, n17653, n17654, n17655, n17656, 
        n17657, n17658, n17659, n17660, n17661, n17662, n17663, 
        n17664, n17665, n17666, n17667, n17668, n17669, n17670, 
        n17671, n17672, n17673, n17674, n17675, n17676, n17677, 
        n17678, n17679, n17680, n17681, n17682, n17683, n17684, 
        n17685, n17686, n17687, n17688, n17689, n17398, n17399, 
        n17400, n17401, n17402, n17403, n17404, n17405, n17406, 
        n17407, n17408, n17409, n17410, n17411, n17412, n17413, 
        n17414, n17415, n17416, n17417, n17418, n17419, n17420, 
        n17421, n17422, n17423, n17424, n17425, n17426, n17427, 
        n17428, n17429, n17430, n17431, n17432, n17433, n17434, 
        n17435, n17436, n17437, n17438, n17439, n17440, n17441, 
        n17442, n17443, n17444, n17445, n17446, n17447, n17448, 
        n17449, n17450, n17451, n17452, n17453, n17454, n17455, 
        n17456, n17457, n17458, n17459, n17460, n17461, n17462, 
        n17463, n17464, n17465, n17466, n17467, n17468, n17469, 
        n17470, n17471, n17472, n17473, n17474, n17475, n17476, 
        n17477, n17478, n17479, n17480, n17481, n17482, n17483, 
        n17484, n17485, n17486, n17487, n17488, n17489, n17490, 
        n17491, n17492, n17493, n17494, n17495, n17496, n17497, 
        n17498, n17499, n17500, n17501, n17502, n17503, n17504, 
        n17505, n17506, n17507, n17508, n17509, n17510, n17511, 
        n17512, n17513, n17514, n17515, n17516, n17517, n17518, 
        n17519, n17520, n17521, n17522, n17523, n17524, n17525, 
        n17526, n17527, n17528, n17529, n17530, n17531, n17532, 
        n17533, n17534, n17535, n17536, n17537, n17538, n17539, 
        n17540, n17541, n17542, n17543, n17690, n17691, n17692, 
        n17693, n17694, n17695, n17696, n17697, n17698, n17699, 
        n17700, n17701, n17702, n17703, n17704, n17705, n17706, 
        n17707, n17708, n17709, n17710, n17711, n17712, n17713, 
        n17714, n17715, n17716, n17717, n17718, n17719, n17720, 
        n17721, n17722, n17723, n17724, n17725, n17726, n17890, 
        n17891, n17892, n17893, n17894, n17895, n17896, n17897, 
        n17898, n17899, n17900, n17901, n17902, n17903, n17904, 
        n17905, n17906, n17907, n17908, n17909, n17910, n17911, 
        n17912, n17913, n17914, n17915, n17916, n17917, n17918, 
        n17919, n17920, n17921, n17922, n17923, n17924, n17925, 
        n17926, n17927, n17928, n17929, n17930, n17931, n17932, 
        n17933, n17934, n17935, n17936, n17937, n17938, n17939, 
        n17940, n17941, n17942, n17943, n17944, n17945, n17946, 
        n17947, n17948, n17949, n17950, n17951, n17952, n17953, 
        n17954, n17955, n17956, n17957, n17958, n17959, n17960, 
        n17961, n17962, n17963, n17964, n17965, n17966, n17967, 
        n17968, n17969, n17970, n17971, n17972, n17973, n17974, 
        n17975, n17976, n17977, n17978, n17979, n17980, n17981, 
        n17982, n17983, n17984, n17985, n17986, n17987, n17988, 
        n17989, n17990, n17991, n17992, n17993, n17994, n17995, 
        n17996, n17997, n17998, n17999, n18000, n18001, n18002, 
        n18003, n18004, n18005, n18006, n18007, n18008, n18009, 
        n18010, n18011, n18012, n18013, n18014, n18015, n18016, 
        n18017, n18018, n18019, n18020, n18021, n18022, n18023, 
        n18024, n18025, n18026, n18027, n18028, n18029, n18030, 
        n18031, n18032, n18033, n18034, n18035, n18036, n18037, 
        n18038, n18039, n18040, n18041, n18042, n18043, n18044, 
        n18045, n18046, n18047, n18048, n18049, n18050, n18051, 
        n18052, n18053, n18054, n18055, n18056, n18057, n18058, 
        n18059, n18060, n18061, n18062, n18063, n18064, n18065, 
        n18066, n18067, n18068, n18069, n18070, n18071, n18072, 
        n17744, n17745, n17746, n17747, n17748, n17749, n17750, 
        n17751, n17752, n17753, n17754, n17755, n17756, n17757, 
        n17758, n17759, n17760, n17761, n17762, n17763, n17764, 
        n17765, n17766, n17767, n17768, n17769, n17770, n17771, 
        n17772, n17773, n17774, n17775, n17776, n17777, n17778, 
        n17779, n17780, n17781, n17782, n17783, n17784, n17785, 
        n17786, n17787, n17788, n17789, n17790, n17791, n17792, 
        n17793, n17794, n17795, n17796, n17797, n17798, n17799, 
        n17800, n17801, n17802, n17803, n17804, n17805, n17806, 
        n17807, n17808, n17809, n17810, n17811, n17812, n17813, 
        n17814, n17815, n17816, n13687, n13688, n13689, n13690, 
        n13691, n13692, n13693, n13694, n13695, n13696, n13697, 
        n13698, n13699, n13700, n13701, n13702, n13703, n13704, 
        n13705, n13706, n13707, n13708, n13709, n13710, n13711, 
        n13712, n13713, n13714, n13715, n13716, n13717, n13718, 
        n13719, n13720, n13721, n13722, n13723, n13724, n13725, 
        n13726, n13727, n13728, n13729, n13730, n13731, n13732, 
        n13733, n13734, n13735, n13736, n13737, n13738, n13739, 
        n13740, n13741, n13742, n13743, n13744, n13745, n13746, 
        n13747, n13748, n13749, n13750, n13751, n13752, n13753, 
        n13754, n13755, n13756, n13757, n13758, n13759, n13760, 
        n13761, n13762, n13763, n13764, n13765, n13766, n13767, 
        n13768, n13769, n13770, n13771, n13772, n13773, n13774, 
        n13775, n13776, n13777, n13778, n13779, n13780, n13781, 
        n13782, n13783, n13784, n13785, n13786, n13787, n13788, 
        n13789, n13790, n13791, n13792, n13793, n13794, n13795, 
        n13796, n13797, n13798, n13799, n13800, n13801, n13802, 
        n13803, n13804, n13805, n13806, n13807, n13808, n13809, 
        n13810, n13811, n13812, n13813, n13814, n13815, n13816, 
        n13817, n13818, n13819, n13820, n13821, n13822, n13823, 
        n13824, n13825, n13826, n13827, n13828, n13829, n13830, 
        n13831, n13832, n13833, n13834, n13835, n13836, n13837, 
        n13838, n13839, n13840, n13841, n13842, n13843, n13844, 
        n13845, n13846, n13847, n13848, n13849, n13850, n13851, 
        n13852, n13853, n13854, n13855, n13856, n13857, n13858, 
        n13859, n13860, n13861, n13862, n13863, n13864, n13865, 
        n13866, n13867, n13868, n13869, n13541, n13542, n13543, 
        n13544, n13545, n13546, n13547, n13548, n13549, n13550, 
        n13551, n13552, n13553, n13554, n13555, n13556, n13557, 
        n13558, n13559, n13560, n13561, n13562, n13563, n13564, 
        n13565, n13566, n13567, n13568, n13569, n13570, n13571, 
        n13572, n13573, n13574, n13575, n13576, n13577, n13578, 
        n13579, n13580, n13581, n13582, n13583, n13584, n13585, 
        n13586, n13587, n13588, n13589, n13590, n13591, n13592, 
        n13593, n13594, n13595, n13596, n13597, n13598, n13599, 
        n13600, n13601, n13602, n13603, n13604, n13605, n13606, 
        n13607, n13608, n13609, n13610, n13611, n13612, n13613, 
        n13614, n13615, n13616, n13617, n13618, n13619, n13620, 
        n13621, n13622, n13623, n13624, n13625, n13626, n13627, 
        n13628, n13629, n13630, n13631, n13632, n13633, n13634, 
        n13635, n13636, n13637, n13638, n13639, n13640, n13641, 
        n13642, n13643, n13644, n13645, n13646, n13647, n13648, 
        n13649, n13650, n13651, n13652, n13653, n13654, n13655, 
        n13656, n13657, n13658, n13659, n13660, n13661, n13662, 
        n13663, n13664, n13665, n13666, n13667, n13668, n13669, 
        n13670, n13671, n13672, n13673, n13674, n13675, n13676, 
        n13677, n13678, n13679, n13680, n13681, n13682, n13683, 
        n13684, n13685, n13686, n17817, n17818, n17819, n17820, 
        n17821, n17822, n17823, n17824, n17825, n17826, n17827, 
        n17828, n17829, n17830, n17831, n17832, n17833, n17834, 
        n17835, n17836, n17837, n17838, n17839, n17840, n17841, 
        n17842, n17843, n17844, n17845, n17846, n17847, n17848, 
        n17849, n17850, n17851, n17852, n17853, n17854, n17855, 
        n17856, n17857, n17858, n17859, n17860, n17861, n17862, 
        n17863, n17864, n17865, n17866, n17867, n17868, n17869, 
        n17870, n17871, n17872, n17873, n17874, n17875, n17876, 
        n17877, n17878, n17879, n17880, n17881, n17882, n17883, 
        n17884, n17885, n17886, n17887, n17888, n17889;
    
    LUT4 mux_391_i22_3_lut_4_lut (.A(op_r_23__N_1106[21]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[21]), .Z(n7431[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i22_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13684_3_lut_4_lut (.A(op_r_23__N_1106[21]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[29] ), .Z(n31429)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13684_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i19_3_lut_4_lut (.A(op_i_23__N_1154[18]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[18]), .Z(n7590[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i19_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13739_3_lut_4_lut (.A(op_i_23__N_1154[18]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[26] ), .Z(n31484)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13739_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i20_3_lut_4_lut (.A(op_i_23__N_1154[19]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[19]), .Z(n7590[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i20_3_lut_4_lut.init = 16'h8f80;
    ALU54B lat_alu_76 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18455), .SIGNEDIB(n18528), .SIGNEDCIN(GND_net), 
           .A35(n18454), .A34(n18453), .A33(n18452), .A32(n18451), .A31(n18450), 
           .A30(n18449), .A29(n18448), .A28(n18447), .A27(n18446), .A26(n18445), 
           .A25(n18444), .A24(n18443), .A23(n18442), .A22(n18441), .A21(n18440), 
           .A20(n18439), .A19(n18438), .A18(n18437), .A17(n18436), .A16(n18435), 
           .A15(n18434), .A14(n18433), .A13(n18432), .A12(n18431), .A11(n18430), 
           .A10(n18429), .A9(n18428), .A8(n18427), .A7(n18426), .A6(n18425), 
           .A5(n18424), .A4(n18423), .A3(n18422), .A2(n18421), .A1(n18420), 
           .A0(n18419), .B35(n18527), .B34(n18526), .B33(n18525), .B32(n18524), 
           .B31(n18523), .B30(n18522), .B29(n18521), .B28(n18520), .B27(n18519), 
           .B26(n18518), .B25(n18517), .B24(n18516), .B23(n18515), .B22(n18514), 
           .B21(n18513), .B20(n18512), .B19(n18511), .B18(n18510), .B17(n18509), 
           .B16(n18508), .B15(n18507), .B14(n18506), .B13(n18505), .B12(n18504), 
           .B11(n18503), .B10(n18502), .B9(n18501), .B8(n18500), .B7(n18499), 
           .B6(n18498), .B5(n18497), .B4(n18496), .B3(n18495), .B2(n18494), 
           .B1(n18493), .B0(n18492), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18491), .MA34(n18490), .MA33(n18489), .MA32(n18488), 
           .MA31(n18487), .MA30(n18486), .MA29(n18485), .MA28(n18484), 
           .MA27(n18483), .MA26(n18482), .MA25(n18481), .MA24(n18480), 
           .MA23(n18479), .MA22(n18478), .MA21(n18477), .MA20(n18476), 
           .MA19(n18475), .MA18(n18474), .MA17(n18473), .MA16(n18472), 
           .MA15(n18471), .MA14(n18470), .MA13(n18469), .MA12(n18468), 
           .MA11(n18467), .MA10(n18466), .MA9(n18465), .MA8(n18464), 
           .MA7(n18463), .MA6(n18462), .MA5(n18461), .MA4(n18460), .MA3(n18459), 
           .MA2(n18458), .MA1(n18457), .MA0(n18456), .MB35(n18564), 
           .MB34(n18563), .MB33(n18562), .MB32(n18561), .MB31(n18560), 
           .MB30(n18559), .MB29(n18558), .MB28(n18557), .MB27(n18556), 
           .MB26(n18555), .MB25(n18554), .MB24(n18553), .MB23(n18552), 
           .MB22(n18551), .MB21(n18550), .MB20(n18549), .MB19(n18548), 
           .MB18(n18547), .MB17(n18546), .MB16(n18545), .MB15(n18544), 
           .MB14(n18543), .MB13(n18542), .MB12(n18541), .MB11(n18540), 
           .MB10(n18539), .MB9(n18538), .MB8(n18537), .MB7(n18536), 
           .MB6(n18535), .MB5(n18534), .MB4(n18533), .MB3(n18532), .MB2(n18531), 
           .MB1(n18530), .MB0(n18529), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R30(n65), .R29(n66), 
           .R28(n67), .R27(n68), .R26(n69), .R25(n70), .R24(n71), 
           .R23(n72), .R22(n73), .R21(n74), .R20(n75), .R19(n76), 
           .R18(n77), .R17(n78), .R16(n79), .R15(n80), .R14(n81), 
           .R13(n82), .R12(n83), .R11(n84), .R10(n85), .R9(n86), .R8(n87), 
           .R7(n88), .R6(n89), .R5(\op_i_23__N_1310[5] ), .R4(\op_i_23__N_1310[4] ), 
           .R3(\op_i_23__N_1310[3] ), .R2(\op_i_23__N_1310[2] ), .R1(\op_i_23__N_1310[1] ), 
           .R0(\op_i_23__N_1310[0] ));
    defparam lat_alu_76.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_76.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_76.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_76.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_76.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_76.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_76.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_76.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_76.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_76.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_76.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_76.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_76.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_76.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_76.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_76.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_76.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_76.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_76.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_76.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_76.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_76.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_76.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_76.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_76.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_76.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_76.REG_FLAG_CLK = "NONE";
    defparam lat_alu_76.REG_FLAG_CE = "CE0";
    defparam lat_alu_76.REG_FLAG_RST = "RST0";
    defparam lat_alu_76.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_76.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_76.MASK01 = "0x00000000000000";
    defparam lat_alu_76.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_76.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_76.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_76.CLK0_DIV = "ENABLED";
    defparam lat_alu_76.CLK1_DIV = "ENABLED";
    defparam lat_alu_76.CLK2_DIV = "ENABLED";
    defparam lat_alu_76.CLK3_DIV = "ENABLED";
    defparam lat_alu_76.MCPAT = "0x00000000000000";
    defparam lat_alu_76.MASKPAT = "0x00000000000000";
    defparam lat_alu_76.RNDPAT = "0x00000000000000";
    defparam lat_alu_76.GSR = "DISABLED";
    defparam lat_alu_76.RESETMODE = "SYNC";
    defparam lat_alu_76.MULT9_MODE = "DISABLED";
    defparam lat_alu_76.LEGACY = "DISABLED";
    MULT18X18D lat_mult_75 (.A17(\rom8_w_i[12] ), .A16(\rom8_w_i[12] ), 
            .A15(\rom8_w_i[12] ), .A14(\rom8_w_i[12] ), .A13(\rom8_w_i[12] ), 
            .A12(\rom8_w_i[12] ), .A11(\rom8_w_i[12] ), .A10(\rom8_w_i[12] ), 
            .A9(\rom8_w_i[12] ), .A8(\rom8_w_i[12] ), .A7(\rom8_w_i[12] ), 
            .A6(\rom8_w_i[12] ), .A5(\rom8_w_i[12] ), .A4(\rom8_w_i[12] ), 
            .A3(\rom8_w_i[12] ), .A2(\rom8_w_i[12] ), .A1(\rom8_w_i[12] ), 
            .A0(\rom8_w_i[12] ), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(GND_net), .B7(GND_net), 
            .B6(GND_net), .B5(n11153), .B4(n11152), .B3(n11151), .B2(n11150), 
            .B1(n11149), .B0(n11148), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n18509), .ROA16(n18508), .ROA15(n18507), .ROA14(n18506), 
            .ROA13(n18505), .ROA12(n18504), .ROA11(n18503), .ROA10(n18502), 
            .ROA9(n18501), .ROA8(n18500), .ROA7(n18499), .ROA6(n18498), 
            .ROA5(n18497), .ROA4(n18496), .ROA3(n18495), .ROA2(n18494), 
            .ROA1(n18493), .ROA0(n18492), .ROB17(n18527), .ROB16(n18526), 
            .ROB15(n18525), .ROB14(n18524), .ROB13(n18523), .ROB12(n18522), 
            .ROB11(n18521), .ROB10(n18520), .ROB9(n18519), .ROB8(n18518), 
            .ROB7(n18517), .ROB6(n18516), .ROB5(n18515), .ROB4(n18514), 
            .ROB3(n18513), .ROB2(n18512), .ROB1(n18511), .ROB0(n18510), 
            .P35(n18564), .P34(n18563), .P33(n18562), .P32(n18561), 
            .P31(n18560), .P30(n18559), .P29(n18558), .P28(n18557), 
            .P27(n18556), .P26(n18555), .P25(n18554), .P24(n18553), 
            .P23(n18552), .P22(n18551), .P21(n18550), .P20(n18549), 
            .P19(n18548), .P18(n18547), .P17(n18546), .P16(n18545), 
            .P15(n18544), .P14(n18543), .P13(n18542), .P12(n18541), 
            .P11(n18540), .P10(n18539), .P9(n18538), .P8(n18537), .P7(n18536), 
            .P6(n18535), .P5(n18534), .P4(n18533), .P3(n18532), .P2(n18531), 
            .P1(n18530), .P0(n18529), .SIGNEDP(n18528));
    defparam lat_mult_75.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_75.REG_INPUTA_CE = "CE0";
    defparam lat_mult_75.REG_INPUTA_RST = "RST0";
    defparam lat_mult_75.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_75.REG_INPUTB_CE = "CE0";
    defparam lat_mult_75.REG_INPUTB_RST = "RST0";
    defparam lat_mult_75.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_75.REG_INPUTC_CE = "CE0";
    defparam lat_mult_75.REG_INPUTC_RST = "RST0";
    defparam lat_mult_75.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_75.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_75.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_75.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_75.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_75.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_75.CLK0_DIV = "ENABLED";
    defparam lat_mult_75.CLK1_DIV = "ENABLED";
    defparam lat_mult_75.CLK2_DIV = "ENABLED";
    defparam lat_mult_75.CLK3_DIV = "ENABLED";
    defparam lat_mult_75.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_75.GSR = "DISABLED";
    defparam lat_mult_75.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_75.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_75.MULT_BYPASS = "DISABLED";
    defparam lat_mult_75.RESETMODE = "SYNC";
    LUT4 i13737_3_lut_4_lut (.A(op_i_23__N_1154[19]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[27] ), .Z(n31482)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13737_3_lut_4_lut.init = 16'hf808;
    MULT18X18D mult_970_mult_2 (.A17(\rom8_w_i[12] ), .A16(\rom8_w_i[12] ), 
            .A15(\rom8_w_i[12] ), .A14(\rom8_w_i[12] ), .A13(\rom8_w_i[12] ), 
            .A12(\rom8_w_i[12] ), .A11(\rom8_w_i[12] ), .A10(\rom8_w_i[12] ), 
            .A9(\rom8_w_i[12] ), .A8(\rom8_w_i[12] ), .A7(\rom8_w_i[2] ), 
            .A6(\rom8_w_i[6] ), .A5(GND_net), .A4(\rom8_w_i[4] ), .A3(\rom8_w_i[3] ), 
            .A2(\rom8_w_i[2] ), .A1(\rom8_w_i[1] ), .A0(\rom8_w_i[0] ), 
            .B17(GND_net), .B16(GND_net), .B15(GND_net), .B14(GND_net), 
            .B13(GND_net), .B12(GND_net), .B11(GND_net), .B10(GND_net), 
            .B9(GND_net), .B8(GND_net), .B7(GND_net), .B6(GND_net), 
            .B5(n11153), .B4(n11152), .B3(n11151), .B2(n11150), .B1(n11149), 
            .B0(n11148), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18436), 
            .ROA16(n18435), .ROA15(n18434), .ROA14(n18433), .ROA13(n18432), 
            .ROA12(n18431), .ROA11(n18430), .ROA10(n18429), .ROA9(n18428), 
            .ROA8(n18427), .ROA7(n18426), .ROA6(n18425), .ROA5(n18424), 
            .ROA4(n18423), .ROA3(n18422), .ROA2(n18421), .ROA1(n18420), 
            .ROA0(n18419), .ROB17(n18454), .ROB16(n18453), .ROB15(n18452), 
            .ROB14(n18451), .ROB13(n18450), .ROB12(n18449), .ROB11(n18448), 
            .ROB10(n18447), .ROB9(n18446), .ROB8(n18445), .ROB7(n18444), 
            .ROB6(n18443), .ROB5(n18442), .ROB4(n18441), .ROB3(n18440), 
            .ROB2(n18439), .ROB1(n18438), .ROB0(n18437), .P35(n18491), 
            .P34(n18490), .P33(n18489), .P32(n18488), .P31(n18487), 
            .P30(n18486), .P29(n18485), .P28(n18484), .P27(n18483), 
            .P26(n18482), .P25(n18481), .P24(n18480), .P23(n18479), 
            .P22(n18478), .P21(n18477), .P20(n18476), .P19(n18475), 
            .P18(n18474), .P17(n18473), .P16(n18472), .P15(n18471), 
            .P14(n18470), .P13(n18469), .P12(n18468), .P11(n18467), 
            .P10(n18466), .P9(n18465), .P8(n18464), .P7(n18463), .P6(n18462), 
            .P5(n18461), .P4(n18460), .P3(n18459), .P2(n18458), .P1(n18457), 
            .P0(n18456), .SIGNEDP(n18455));
    defparam mult_970_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_970_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_970_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_970_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_970_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_970_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_970_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_970_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_970_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_970_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_970_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_970_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_970_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_970_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_970_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_970_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_970_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_970_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_970_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_970_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_970_mult_2.GSR = "DISABLED";
    defparam mult_970_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_970_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_970_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_970_mult_2.RESETMODE = "SYNC";
    LUT4 mux_391_i19_3_lut_4_lut (.A(op_r_23__N_1106[18]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[18]), .Z(n7431[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i19_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13690_3_lut_4_lut (.A(op_r_23__N_1106[18]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[26] ), .Z(n31435)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13690_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i20_3_lut_4_lut (.A(op_r_23__N_1106[19]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[19]), .Z(n7431[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13688_3_lut_4_lut (.A(op_r_23__N_1106[19]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[27] ), .Z(n31433)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13688_3_lut_4_lut.init = 16'hf808;
    MULT18X18D lat_mult_61 (.A17(shift_8_dout_i[17]), .A16(shift_8_dout_i[16]), 
            .A15(shift_8_dout_i[15]), .A14(shift_8_dout_i[14]), .A13(shift_8_dout_i[13]), 
            .A12(shift_8_dout_i[12]), .A11(shift_8_dout_i[11]), .A10(shift_8_dout_i[10]), 
            .A9(shift_8_dout_i[9]), .A8(shift_8_dout_i[8]), .A7(shift_8_dout_i[7]), 
            .A6(shift_8_dout_i[6]), .A5(shift_8_dout_i[5]), .A4(shift_8_dout_i[4]), 
            .A3(shift_8_dout_i[3]), .A2(shift_8_dout_i[2]), .A1(shift_8_dout_i[1]), 
            .A0(shift_8_dout_i[0]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n119), .B8(n119), .B7(n119), .B6(n119), .B5(n119), 
            .B4(n119), .B3(n119), .B2(n119), .B1(n119), .B0(n119), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17561), .ROA16(n17560), 
            .ROA15(n17559), .ROA14(n17558), .ROA13(n17557), .ROA12(n17556), 
            .ROA11(n17555), .ROA10(n17554), .ROA9(n17553), .ROA8(n17552), 
            .ROA7(n17551), .ROA6(n17550), .ROA5(n17549), .ROA4(n17548), 
            .ROA3(n17547), .ROA2(n17546), .ROA1(n17545), .ROA0(n17544), 
            .ROB17(n17579), .ROB16(n17578), .ROB15(n17577), .ROB14(n17576), 
            .ROB13(n17575), .ROB12(n17574), .ROB11(n17573), .ROB10(n17572), 
            .ROB9(n17571), .ROB8(n17570), .ROB7(n17569), .ROB6(n17568), 
            .ROB5(n17567), .ROB4(n17566), .ROB3(n17565), .ROB2(n17564), 
            .ROB1(n17563), .ROB0(n17562), .P35(n17616), .P34(n17615), 
            .P33(n17614), .P32(n17613), .P31(n17612), .P30(n17611), 
            .P29(n17610), .P28(n17609), .P27(n17608), .P26(n17607), 
            .P25(n17606), .P24(n17605), .P23(n17604), .P22(n17603), 
            .P21(n17602), .P20(n17601), .P19(n17600), .P18(n17599), 
            .P17(n17598), .P16(n17597), .P15(n17596), .P14(n17595), 
            .P13(n17594), .P12(n17593), .P11(n17592), .P10(n17591), 
            .P9(n17590), .P8(n17589), .P7(n17588), .P6(n17587), .P5(n17586), 
            .P4(n17585), .P3(n17584), .P2(n17583), .P1(n17582), .P0(n17581), 
            .SIGNEDP(n17580));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_61.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_61.REG_INPUTA_CE = "CE0";
    defparam lat_mult_61.REG_INPUTA_RST = "RST0";
    defparam lat_mult_61.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_61.REG_INPUTB_CE = "CE0";
    defparam lat_mult_61.REG_INPUTB_RST = "RST0";
    defparam lat_mult_61.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_61.REG_INPUTC_CE = "CE0";
    defparam lat_mult_61.REG_INPUTC_RST = "RST0";
    defparam lat_mult_61.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_61.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_61.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_61.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_61.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_61.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_61.CLK0_DIV = "ENABLED";
    defparam lat_mult_61.CLK1_DIV = "ENABLED";
    defparam lat_mult_61.CLK2_DIV = "ENABLED";
    defparam lat_mult_61.CLK3_DIV = "ENABLED";
    defparam lat_mult_61.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_61.GSR = "DISABLED";
    defparam lat_mult_61.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_61.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_61.MULT_BYPASS = "DISABLED";
    defparam lat_mult_61.RESETMODE = "SYNC";
    MULT18X18D lat_mult_62 (.A17(shift_8_dout_i[23]), .A16(shift_8_dout_i[23]), 
            .A15(shift_8_dout_i[23]), .A14(shift_8_dout_i[23]), .A13(shift_8_dout_i[23]), 
            .A12(shift_8_dout_i[23]), .A11(shift_8_dout_i[23]), .A10(shift_8_dout_i[23]), 
            .A9(shift_8_dout_i[23]), .A8(shift_8_dout_i[23]), .A7(shift_8_dout_i[23]), 
            .A6(shift_8_dout_i[23]), .A5(shift_8_dout_i[23]), .A4(shift_8_dout_i[22]), 
            .A3(shift_8_dout_i[21]), .A2(shift_8_dout_i[20]), .A1(shift_8_dout_i[19]), 
            .A0(shift_8_dout_i[18]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n119), .B8(n119), .B7(n119), .B6(n119), .B5(n119), 
            .B4(n119), .B3(n119), .B2(n119), .B1(n119), .B0(n119), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17634), .ROA16(n17633), 
            .ROA15(n17632), .ROA14(n17631), .ROA13(n17630), .ROA12(n17629), 
            .ROA11(n17628), .ROA10(n17627), .ROA9(n17626), .ROA8(n17625), 
            .ROA7(n17624), .ROA6(n17623), .ROA5(n17622), .ROA4(n17621), 
            .ROA3(n17620), .ROA2(n17619), .ROA1(n17618), .ROA0(n17617), 
            .ROB17(n17652), .ROB16(n17651), .ROB15(n17650), .ROB14(n17649), 
            .ROB13(n17648), .ROB12(n17647), .ROB11(n17646), .ROB10(n17645), 
            .ROB9(n17644), .ROB8(n17643), .ROB7(n17642), .ROB6(n17641), 
            .ROB5(n17640), .ROB4(n17639), .ROB3(n17638), .ROB2(n17637), 
            .ROB1(n17636), .ROB0(n17635), .P35(n17689), .P34(n17688), 
            .P33(n17687), .P32(n17686), .P31(n17685), .P30(n17684), 
            .P29(n17683), .P28(n17682), .P27(n17681), .P26(n17680), 
            .P25(n17679), .P24(n17678), .P23(n17677), .P22(n17676), 
            .P21(n17675), .P20(n17674), .P19(n17673), .P18(n17672), 
            .P17(n17671), .P16(n17670), .P15(n17669), .P14(n17668), 
            .P13(n17667), .P12(n17666), .P11(n17665), .P10(n17664), 
            .P9(n17663), .P8(n17662), .P7(n17661), .P6(n17660), .P5(n17659), 
            .P4(n17658), .P3(n17657), .P2(n17656), .P1(n17655), .P0(n17654), 
            .SIGNEDP(n17653));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_62.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_62.REG_INPUTA_CE = "CE0";
    defparam lat_mult_62.REG_INPUTA_RST = "RST0";
    defparam lat_mult_62.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_62.REG_INPUTB_CE = "CE0";
    defparam lat_mult_62.REG_INPUTB_RST = "RST0";
    defparam lat_mult_62.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_62.REG_INPUTC_CE = "CE0";
    defparam lat_mult_62.REG_INPUTC_RST = "RST0";
    defparam lat_mult_62.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_62.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_62.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_62.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_62.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_62.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_62.CLK0_DIV = "ENABLED";
    defparam lat_mult_62.CLK1_DIV = "ENABLED";
    defparam lat_mult_62.CLK2_DIV = "ENABLED";
    defparam lat_mult_62.CLK3_DIV = "ENABLED";
    defparam lat_mult_62.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_62.GSR = "DISABLED";
    defparam lat_mult_62.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_62.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_62.MULT_BYPASS = "DISABLED";
    defparam lat_mult_62.RESETMODE = "SYNC";
    ALU54B lat_alu_63 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n17434), .SIGNEDIB(n17507), .SIGNEDCIN(GND_net), 
           .A35(n17433), .A34(n17432), .A33(n17431), .A32(n17430), .A31(n17429), 
           .A30(n17428), .A29(n17427), .A28(n17426), .A27(n17425), .A26(n17424), 
           .A25(n17423), .A24(n17422), .A23(n17421), .A22(n17420), .A21(n17419), 
           .A20(n17418), .A19(n17417), .A18(n17416), .A17(n17415), .A16(n17414), 
           .A15(n17413), .A14(n17412), .A13(n17411), .A12(n17410), .A11(n17409), 
           .A10(n17408), .A9(n17407), .A8(n17406), .A7(n17405), .A6(n17404), 
           .A5(n17403), .A4(n17402), .A3(n17401), .A2(n17400), .A1(n17399), 
           .A0(n17398), .B35(n17506), .B34(n17505), .B33(n17504), .B32(n17503), 
           .B31(n17502), .B30(n17501), .B29(n17500), .B28(n17499), .B27(n17498), 
           .B26(n17497), .B25(n17496), .B24(n17495), .B23(n17494), .B22(n17493), 
           .B21(n17492), .B20(n17491), .B19(n17490), .B18(n17489), .B17(n17488), 
           .B16(n17487), .B15(n17486), .B14(n17485), .B13(n17484), .B12(n17483), 
           .B11(n17482), .B10(n17481), .B9(n17480), .B8(n17479), .B7(n17478), 
           .B6(n17477), .B5(n17476), .B4(n17475), .B3(n17474), .B2(n17473), 
           .B1(n17472), .B0(n17471), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n17470), .MA34(n17469), .MA33(n17468), .MA32(n17467), 
           .MA31(n17466), .MA30(n17465), .MA29(n17464), .MA28(n17463), 
           .MA27(n17462), .MA26(n17461), .MA25(n17460), .MA24(n17459), 
           .MA23(n17458), .MA22(n17457), .MA21(n17456), .MA20(n17455), 
           .MA19(n17454), .MA18(n17453), .MA17(n17452), .MA16(n17451), 
           .MA15(n17450), .MA14(n17449), .MA13(n17448), .MA12(n17447), 
           .MA11(n17446), .MA10(n17445), .MA9(n17444), .MA8(n17443), 
           .MA7(n17442), .MA6(n17441), .MA5(n17440), .MA4(n17439), .MA3(n17438), 
           .MA2(n17437), .MA1(n17436), .MA0(n17435), .MB35(n17543), 
           .MB34(n17542), .MB33(n17541), .MB32(n17540), .MB31(n17539), 
           .MB30(n17538), .MB29(n17537), .MB28(n17536), .MB27(n17535), 
           .MB26(n17534), .MB25(n17533), .MB24(n17532), .MB23(n17531), 
           .MB22(n17530), .MB21(n17529), .MB20(n17528), .MB19(n17527), 
           .MB18(n17526), .MB17(n17525), .MB16(n17524), .MB15(n17523), 
           .MB14(n17522), .MB13(n17521), .MB12(n17520), .MB11(n17519), 
           .MB10(n17518), .MB9(n17517), .MB8(n17516), .MB7(n17515), 
           .MB6(n17514), .MB5(n17513), .MB4(n17512), .MB3(n17511), .MB2(n17510), 
           .MB1(n17509), .MB0(n17508), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n17725), 
           .R52(n17724), .R51(n17723), .R50(n17722), .R49(n17721), .R48(n17720), 
           .R47(n17719), .R46(n17718), .R45(n17717), .R44(n17716), .R43(n17715), 
           .R42(n17714), .R41(n17713), .R40(n17712), .R39(n17711), .R38(n17710), 
           .R37(n17709), .R36(n17708), .R35(n17707), .R34(n17706), .R33(n17705), 
           .R32(n17704), .R31(n17703), .R30(n17702), .R29(n17701), .R28(n17700), 
           .R27(n17699), .R26(n17698), .R25(n17697), .R24(n17696), .R23(n17695), 
           .R22(n17694), .R21(n17693), .R20(n17692), .R19(n17691), .R18(n17690), 
           .R17(\op_r_23__N_1268[17] ), .R16(\op_r_23__N_1268[16] ), .R15(\op_r_23__N_1268[15] ), 
           .R14(\op_r_23__N_1268[14] ), .R13(\op_r_23__N_1268[13] ), .R12(\op_r_23__N_1268[12] ), 
           .R11(\op_r_23__N_1268[11] ), .R10(\op_r_23__N_1268[10] ), .R9(\op_r_23__N_1268[9] ), 
           .R8(\op_r_23__N_1268[8] ), .R7(\op_r_23__N_1268[7] ), .R6(\op_r_23__N_1268[6] ), 
           .R5(\op_r_23__N_1268[5] ), .R4(\op_r_23__N_1268[4] ), .R3(\op_r_23__N_1268[3] ), 
           .R2(\op_r_23__N_1268[2] ), .R1(\op_r_23__N_1268[1] ), .R0(\op_r_23__N_1268[0] ), 
           .SIGNEDR(n17726));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_63.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_63.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_63.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_63.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_63.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_63.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_63.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_63.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_63.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_63.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_63.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_63.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_63.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_63.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_63.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_63.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_63.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_63.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_63.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_63.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_63.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_63.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_63.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_63.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_63.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_63.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_63.REG_FLAG_CLK = "NONE";
    defparam lat_alu_63.REG_FLAG_CE = "CE0";
    defparam lat_alu_63.REG_FLAG_RST = "RST0";
    defparam lat_alu_63.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_63.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_63.MASK01 = "0x00000000000000";
    defparam lat_alu_63.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_63.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_63.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_63.CLK0_DIV = "ENABLED";
    defparam lat_alu_63.CLK1_DIV = "ENABLED";
    defparam lat_alu_63.CLK2_DIV = "ENABLED";
    defparam lat_alu_63.CLK3_DIV = "ENABLED";
    defparam lat_alu_63.MCPAT = "0x00000000000000";
    defparam lat_alu_63.MASKPAT = "0x00000000000000";
    defparam lat_alu_63.RNDPAT = "0x00000000000000";
    defparam lat_alu_63.GSR = "DISABLED";
    defparam lat_alu_63.RESETMODE = "SYNC";
    defparam lat_alu_63.MULT9_MODE = "DISABLED";
    defparam lat_alu_63.LEGACY = "DISABLED";
    ALU54B lat_alu_64 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n17580), .SIGNEDIB(n17653), .SIGNEDCIN(n17726), .A35(n17579), 
           .A34(n17578), .A33(n17577), .A32(n17576), .A31(n17575), .A30(n17574), 
           .A29(n17573), .A28(n17572), .A27(n17571), .A26(n17570), .A25(n17569), 
           .A24(n17568), .A23(n17567), .A22(n17566), .A21(n17565), .A20(n17564), 
           .A19(n17563), .A18(n17562), .A17(n17561), .A16(n17560), .A15(n17559), 
           .A14(n17558), .A13(n17557), .A12(n17556), .A11(n17555), .A10(n17554), 
           .A9(n17553), .A8(n17552), .A7(n17551), .A6(n17550), .A5(n17549), 
           .A4(n17548), .A3(n17547), .A2(n17546), .A1(n17545), .A0(n17544), 
           .B35(n17652), .B34(n17651), .B33(n17650), .B32(n17649), .B31(n17648), 
           .B30(n17647), .B29(n17646), .B28(n17645), .B27(n17644), .B26(n17643), 
           .B25(n17642), .B24(n17641), .B23(n17640), .B22(n17639), .B21(n17638), 
           .B20(n17637), .B19(n17636), .B18(n17635), .B17(n17634), .B16(n17633), 
           .B15(n17632), .B14(n17631), .B13(n17630), .B12(n17629), .B11(n17628), 
           .B10(n17627), .B9(n17626), .B8(n17625), .B7(n17624), .B6(n17623), 
           .B5(n17622), .B4(n17621), .B3(n17620), .B2(n17619), .B1(n17618), 
           .B0(n17617), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n17616), .MA34(n17615), .MA33(n17614), .MA32(n17613), 
           .MA31(n17612), .MA30(n17611), .MA29(n17610), .MA28(n17609), 
           .MA27(n17608), .MA26(n17607), .MA25(n17606), .MA24(n17605), 
           .MA23(n17604), .MA22(n17603), .MA21(n17602), .MA20(n17601), 
           .MA19(n17600), .MA18(n17599), .MA17(n17598), .MA16(n17597), 
           .MA15(n17596), .MA14(n17595), .MA13(n17594), .MA12(n17593), 
           .MA11(n17592), .MA10(n17591), .MA9(n17590), .MA8(n17589), 
           .MA7(n17588), .MA6(n17587), .MA5(n17586), .MA4(n17585), .MA3(n17584), 
           .MA2(n17583), .MA1(n17582), .MA0(n17581), .MB35(n17689), 
           .MB34(n17688), .MB33(n17687), .MB32(n17686), .MB31(n17685), 
           .MB30(n17684), .MB29(n17683), .MB28(n17682), .MB27(n17681), 
           .MB26(n17680), .MB25(n17679), .MB24(n17678), .MB23(n17677), 
           .MB22(n17676), .MB21(n17675), .MB20(n17674), .MB19(n17673), 
           .MB18(n17672), .MB17(n17671), .MB16(n17670), .MB15(n17669), 
           .MB14(n17668), .MB13(n17667), .MB12(n17666), .MB11(n17665), 
           .MB10(n17664), .MB9(n17663), .MB8(n17662), .MB7(n17661), 
           .MB6(n17660), .MB5(n17659), .MB4(n17658), .MB3(n17657), .MB2(n17656), 
           .MB1(n17655), .MB0(n17654), .CIN53(n17725), .CIN52(n17724), 
           .CIN51(n17723), .CIN50(n17722), .CIN49(n17721), .CIN48(n17720), 
           .CIN47(n17719), .CIN46(n17718), .CIN45(n17717), .CIN44(n17716), 
           .CIN43(n17715), .CIN42(n17714), .CIN41(n17713), .CIN40(n17712), 
           .CIN39(n17711), .CIN38(n17710), .CIN37(n17709), .CIN36(n17708), 
           .CIN35(n17707), .CIN34(n17706), .CIN33(n17705), .CIN32(n17704), 
           .CIN31(n17703), .CIN30(n17702), .CIN29(n17701), .CIN28(n17700), 
           .CIN27(n17699), .CIN26(n17698), .CIN25(n17697), .CIN24(n17696), 
           .CIN23(n17695), .CIN22(n17694), .CIN21(n17693), .CIN20(n17692), 
           .CIN19(n17691), .CIN18(n17690), .CIN17(\op_r_23__N_1268[17] ), 
           .CIN16(\op_r_23__N_1268[16] ), .CIN15(\op_r_23__N_1268[15] ), 
           .CIN14(\op_r_23__N_1268[14] ), .CIN13(\op_r_23__N_1268[13] ), 
           .CIN12(\op_r_23__N_1268[12] ), .CIN11(\op_r_23__N_1268[11] ), 
           .CIN10(\op_r_23__N_1268[10] ), .CIN9(\op_r_23__N_1268[9] ), .CIN8(\op_r_23__N_1268[8] ), 
           .CIN7(\op_r_23__N_1268[7] ), .CIN6(\op_r_23__N_1268[6] ), .CIN5(\op_r_23__N_1268[5] ), 
           .CIN4(\op_r_23__N_1268[4] ), .CIN3(\op_r_23__N_1268[3] ), .CIN2(\op_r_23__N_1268[2] ), 
           .CIN1(\op_r_23__N_1268[1] ), .CIN0(\op_r_23__N_1268[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1268[31] ), 
           .R12(\op_r_23__N_1268[30] ), .R11(\op_r_23__N_1268[29] ), .R10(\op_r_23__N_1268[28] ), 
           .R9(\op_r_23__N_1268[27] ), .R8(\op_r_23__N_1268[26] ), .R7(\op_r_23__N_1268[25] ), 
           .R6(\op_r_23__N_1268[24] ), .R5(\op_r_23__N_1268[23] ), .R4(\op_r_23__N_1268[22] ), 
           .R3(\op_r_23__N_1268[21] ), .R2(\op_r_23__N_1268[20] ), .R1(\op_r_23__N_1268[19] ), 
           .R0(\op_r_23__N_1268[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_64.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_64.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_64.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_64.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_64.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_64.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_64.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_64.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_64.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_64.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_64.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_64.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_64.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_64.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_64.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_64.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_64.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_64.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_64.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_64.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_64.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_64.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_64.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_64.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_64.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_64.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_64.REG_FLAG_CLK = "NONE";
    defparam lat_alu_64.REG_FLAG_CE = "CE0";
    defparam lat_alu_64.REG_FLAG_RST = "RST0";
    defparam lat_alu_64.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_64.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_64.MASK01 = "0x00000000000000";
    defparam lat_alu_64.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_64.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_64.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_64.CLK0_DIV = "ENABLED";
    defparam lat_alu_64.CLK1_DIV = "ENABLED";
    defparam lat_alu_64.CLK2_DIV = "ENABLED";
    defparam lat_alu_64.CLK3_DIV = "ENABLED";
    defparam lat_alu_64.MCPAT = "0x00000000000000";
    defparam lat_alu_64.MASKPAT = "0x00000000000000";
    defparam lat_alu_64.RNDPAT = "0x00000000000000";
    defparam lat_alu_64.GSR = "DISABLED";
    defparam lat_alu_64.RESETMODE = "SYNC";
    defparam lat_alu_64.MULT9_MODE = "DISABLED";
    defparam lat_alu_64.LEGACY = "DISABLED";
    ALU54B lat_alu_69 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n17926), .SIGNEDIB(n17999), .SIGNEDCIN(n18072), .A35(n17925), 
           .A34(n17924), .A33(n17923), .A32(n17922), .A31(n17921), .A30(n17920), 
           .A29(n17919), .A28(n17918), .A27(n17917), .A26(n17916), .A25(n17915), 
           .A24(n17914), .A23(n17913), .A22(n17912), .A21(n17911), .A20(n17910), 
           .A19(n17909), .A18(n17908), .A17(n17907), .A16(n17906), .A15(n17905), 
           .A14(n17904), .A13(n17903), .A12(n17902), .A11(n17901), .A10(n17900), 
           .A9(n17899), .A8(n17898), .A7(n17897), .A6(n17896), .A5(n17895), 
           .A4(n17894), .A3(n17893), .A2(n17892), .A1(n17891), .A0(n17890), 
           .B35(n17998), .B34(n17997), .B33(n17996), .B32(n17995), .B31(n17994), 
           .B30(n17993), .B29(n17992), .B28(n17991), .B27(n17990), .B26(n17989), 
           .B25(n17988), .B24(n17987), .B23(n17986), .B22(n17985), .B21(n17984), 
           .B20(n17983), .B19(n17982), .B18(n17981), .B17(n17980), .B16(n17979), 
           .B15(n17978), .B14(n17977), .B13(n17976), .B12(n17975), .B11(n17974), 
           .B10(n17973), .B9(n17972), .B8(n17971), .B7(n17970), .B6(n17969), 
           .B5(n17968), .B4(n17967), .B3(n17966), .B2(n17965), .B1(n17964), 
           .B0(n17963), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n17962), .MA34(n17961), .MA33(n17960), .MA32(n17959), 
           .MA31(n17958), .MA30(n17957), .MA29(n17956), .MA28(n17955), 
           .MA27(n17954), .MA26(n17953), .MA25(n17952), .MA24(n17951), 
           .MA23(n17950), .MA22(n17949), .MA21(n17948), .MA20(n17947), 
           .MA19(n17946), .MA18(n17945), .MA17(n17944), .MA16(n17943), 
           .MA15(n17942), .MA14(n17941), .MA13(n17940), .MA12(n17939), 
           .MA11(n17938), .MA10(n17937), .MA9(n17936), .MA8(n17935), 
           .MA7(n17934), .MA6(n17933), .MA5(n17932), .MA4(n17931), .MA3(n17930), 
           .MA2(n17929), .MA1(n17928), .MA0(n17927), .MB35(n18035), 
           .MB34(n18034), .MB33(n18033), .MB32(n18032), .MB31(n18031), 
           .MB30(n18030), .MB29(n18029), .MB28(n18028), .MB27(n18027), 
           .MB26(n18026), .MB25(n18025), .MB24(n18024), .MB23(n18023), 
           .MB22(n18022), .MB21(n18021), .MB20(n18020), .MB19(n18019), 
           .MB18(n18018), .MB17(n18017), .MB16(n18016), .MB15(n18015), 
           .MB14(n18014), .MB13(n18013), .MB12(n18012), .MB11(n18011), 
           .MB10(n18010), .MB9(n18009), .MB8(n18008), .MB7(n18007), 
           .MB6(n18006), .MB5(n18005), .MB4(n18004), .MB3(n18003), .MB2(n18002), 
           .MB1(n18001), .MB0(n18000), .CIN53(n18071), .CIN52(n18070), 
           .CIN51(n18069), .CIN50(n18068), .CIN49(n18067), .CIN48(n18066), 
           .CIN47(n18065), .CIN46(n18064), .CIN45(n18063), .CIN44(n18062), 
           .CIN43(n18061), .CIN42(n18060), .CIN41(n18059), .CIN40(n18058), 
           .CIN39(n18057), .CIN38(n18056), .CIN37(n18055), .CIN36(n18054), 
           .CIN35(n18053), .CIN34(n18052), .CIN33(n18051), .CIN32(n18050), 
           .CIN31(n18049), .CIN30(n18048), .CIN29(n18047), .CIN28(n18046), 
           .CIN27(n18045), .CIN26(n18044), .CIN25(n18043), .CIN24(n18042), 
           .CIN23(n18041), .CIN22(n18040), .CIN21(n18039), .CIN20(n18038), 
           .CIN19(n18037), .CIN18(n18036), .CIN17(\op_r_23__N_1226[17] ), 
           .CIN16(\op_r_23__N_1226[16] ), .CIN15(\op_r_23__N_1226[15] ), 
           .CIN14(\op_r_23__N_1226[14] ), .CIN13(\op_r_23__N_1226[13] ), 
           .CIN12(\op_r_23__N_1226[12] ), .CIN11(\op_r_23__N_1226[11] ), 
           .CIN10(\op_r_23__N_1226[10] ), .CIN9(\op_r_23__N_1226[9] ), .CIN8(\op_r_23__N_1226[8] ), 
           .CIN7(\op_r_23__N_1226[7] ), .CIN6(\op_r_23__N_1226[6] ), .CIN5(\op_r_23__N_1226[5] ), 
           .CIN4(\op_r_23__N_1226[4] ), .CIN3(\op_r_23__N_1226[3] ), .CIN2(\op_r_23__N_1226[2] ), 
           .CIN1(\op_r_23__N_1226[1] ), .CIN0(\op_r_23__N_1226[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1226[31] ), 
           .R12(\op_r_23__N_1226[30] ), .R11(\op_r_23__N_1226[29] ), .R10(\op_r_23__N_1226[28] ), 
           .R9(\op_r_23__N_1226[27] ), .R8(\op_r_23__N_1226[26] ), .R7(\op_r_23__N_1226[25] ), 
           .R6(\op_r_23__N_1226[24] ), .R5(\op_r_23__N_1226[23] ), .R4(\op_r_23__N_1226[22] ), 
           .R3(\op_r_23__N_1226[21] ), .R2(\op_r_23__N_1226[20] ), .R1(\op_r_23__N_1226[19] ), 
           .R0(\op_r_23__N_1226[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_69.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_69.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_69.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_69.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_69.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_69.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_69.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_69.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_69.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_69.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_69.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_69.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_69.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_69.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_69.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_69.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_69.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_69.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_69.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_69.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_69.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_69.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_69.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_69.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_69.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_69.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_69.REG_FLAG_CLK = "NONE";
    defparam lat_alu_69.REG_FLAG_CE = "CE0";
    defparam lat_alu_69.REG_FLAG_RST = "RST0";
    defparam lat_alu_69.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_69.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_69.MASK01 = "0x00000000000000";
    defparam lat_alu_69.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_69.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_69.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_69.CLK0_DIV = "ENABLED";
    defparam lat_alu_69.CLK1_DIV = "ENABLED";
    defparam lat_alu_69.CLK2_DIV = "ENABLED";
    defparam lat_alu_69.CLK3_DIV = "ENABLED";
    defparam lat_alu_69.MCPAT = "0x00000000000000";
    defparam lat_alu_69.MASKPAT = "0x00000000000000";
    defparam lat_alu_69.RNDPAT = "0x00000000000000";
    defparam lat_alu_69.GSR = "DISABLED";
    defparam lat_alu_69.RESETMODE = "SYNC";
    defparam lat_alu_69.MULT9_MODE = "DISABLED";
    defparam lat_alu_69.LEGACY = "DISABLED";
    LUT4 mux_403_i17_3_lut_4_lut (.A(op_i_23__N_1154[16]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[16]), .Z(n7590[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13743_3_lut_4_lut (.A(op_i_23__N_1154[16]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[24] ), .Z(n31488)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13743_3_lut_4_lut.init = 16'hf808;
    MULT18X18D mult_10_mult_2 (.A17(\rom8_w_r[10] ), .A16(\rom8_w_r[10] ), 
            .A15(\rom8_w_r[10] ), .A14(\rom8_w_r[10] ), .A13(\rom8_w_r[10] ), 
            .A12(\rom8_w_r[10] ), .A11(\rom8_w_r[10] ), .A10(\rom8_w_r[10] ), 
            .A9(\rom8_w_r[10] ), .A8(\rom8_w_r[8] ), .A7(\rom8_w_r[7] ), 
            .A6(\rom8_w_r[6] ), .A5(\rom8_w_r[5] ), .A4(\rom8_w_r[4] ), 
            .A3(\rom8_w_r[3] ), .A2(\rom8_w_r[7] ), .A1(\rom8_w_r[1] ), 
            .A0(\rom8_w_r[0] ), .B17(n12287), .B16(n12286), .B15(n12285), 
            .B14(n12284), .B13(n12283), .B12(n12282), .B11(n12281), 
            .B10(n12280), .B9(n12279), .B8(n12278), .B7(n12277), .B6(n12276), 
            .B5(n12275), .B4(n12274), .B3(n12273), .B2(n12272), .B1(n12271), 
            .B0(n12270), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17761), 
            .ROA16(n17760), .ROA15(n17759), .ROA14(n17758), .ROA13(n17757), 
            .ROA12(n17756), .ROA11(n17755), .ROA10(n17754), .ROA9(n17753), 
            .ROA8(n17752), .ROA7(n17751), .ROA6(n17750), .ROA5(n17749), 
            .ROA4(n17748), .ROA3(n17747), .ROA2(n17746), .ROA1(n17745), 
            .ROA0(n17744), .ROB17(n17779), .ROB16(n17778), .ROB15(n17777), 
            .ROB14(n17776), .ROB13(n17775), .ROB12(n17774), .ROB11(n17773), 
            .ROB10(n17772), .ROB9(n17771), .ROB8(n17770), .ROB7(n17769), 
            .ROB6(n17768), .ROB5(n17767), .ROB4(n17766), .ROB3(n17765), 
            .ROB2(n17764), .ROB1(n17763), .ROB0(n17762), .P35(n17816), 
            .P34(n17815), .P33(n17814), .P32(n17813), .P31(n17812), 
            .P30(n17811), .P29(n17810), .P28(n17809), .P27(n17808), 
            .P26(n17807), .P25(n17806), .P24(n17805), .P23(n17804), 
            .P22(n17803), .P21(n17802), .P20(n17801), .P19(n17800), 
            .P18(n17799), .P17(n17798), .P16(n17797), .P15(n17796), 
            .P14(n17795), .P13(n17794), .P12(n17793), .P11(n17792), 
            .P10(n17791), .P9(n17790), .P8(n17789), .P7(n17788), .P6(n17787), 
            .P5(n17786), .P4(n17785), .P3(n17784), .P2(n17783), .P1(n17782), 
            .P0(n17781), .SIGNEDP(n17780));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam mult_10_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_10_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_10_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_10_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_10_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_10_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_10_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_10_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_10_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_10_mult_2.GSR = "DISABLED";
    defparam mult_10_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_10_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_10_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_10_mult_2.RESETMODE = "SYNC";
    LUT4 mux_403_i18_3_lut_4_lut (.A(op_i_23__N_1154[17]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[17]), .Z(n7590[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i18_3_lut_4_lut.init = 16'h8f80;
    ALU54B lat_alu_9 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n13723), .SIGNEDIB(n13796), .SIGNEDCIN(n13869), .A35(n13722), 
           .A34(n13721), .A33(n13720), .A32(n13719), .A31(n13718), .A30(n13717), 
           .A29(n13716), .A28(n13715), .A27(n13714), .A26(n13713), .A25(n13712), 
           .A24(n13711), .A23(n13710), .A22(n13709), .A21(n13708), .A20(n13707), 
           .A19(n13706), .A18(n13705), .A17(n13704), .A16(n13703), .A15(n13702), 
           .A14(n13701), .A13(n13700), .A12(n13699), .A11(n13698), .A10(n13697), 
           .A9(n13696), .A8(n13695), .A7(n13694), .A6(n13693), .A5(n13692), 
           .A4(n13691), .A3(n13690), .A2(n13689), .A1(n13688), .A0(n13687), 
           .B35(n13795), .B34(n13794), .B33(n13793), .B32(n13792), .B31(n13791), 
           .B30(n13790), .B29(n13789), .B28(n13788), .B27(n13787), .B26(n13786), 
           .B25(n13785), .B24(n13784), .B23(n13783), .B22(n13782), .B21(n13781), 
           .B20(n13780), .B19(n13779), .B18(n13778), .B17(n13777), .B16(n13776), 
           .B15(n13775), .B14(n13774), .B13(n13773), .B12(n13772), .B11(n13771), 
           .B10(n13770), .B9(n13769), .B8(n13768), .B7(n13767), .B6(n13766), 
           .B5(n13765), .B4(n13764), .B3(n13763), .B2(n13762), .B1(n13761), 
           .B0(n13760), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n13759), .MA34(n13758), .MA33(n13757), .MA32(n13756), 
           .MA31(n13755), .MA30(n13754), .MA29(n13753), .MA28(n13752), 
           .MA27(n13751), .MA26(n13750), .MA25(n13749), .MA24(n13748), 
           .MA23(n13747), .MA22(n13746), .MA21(n13745), .MA20(n13744), 
           .MA19(n13743), .MA18(n13742), .MA17(n13741), .MA16(n13740), 
           .MA15(n13739), .MA14(n13738), .MA13(n13737), .MA12(n13736), 
           .MA11(n13735), .MA10(n13734), .MA9(n13733), .MA8(n13732), 
           .MA7(n13731), .MA6(n13730), .MA5(n13729), .MA4(n13728), .MA3(n13727), 
           .MA2(n13726), .MA1(n13725), .MA0(n13724), .MB35(n13832), 
           .MB34(n13831), .MB33(n13830), .MB32(n13829), .MB31(n13828), 
           .MB30(n13827), .MB29(n13826), .MB28(n13825), .MB27(n13824), 
           .MB26(n13823), .MB25(n13822), .MB24(n13821), .MB23(n13820), 
           .MB22(n13819), .MB21(n13818), .MB20(n13817), .MB19(n13816), 
           .MB18(n13815), .MB17(n13814), .MB16(n13813), .MB15(n13812), 
           .MB14(n13811), .MB13(n13810), .MB12(n13809), .MB11(n13808), 
           .MB10(n13807), .MB9(n13806), .MB8(n13805), .MB7(n13804), 
           .MB6(n13803), .MB5(n13802), .MB4(n13801), .MB3(n13800), .MB2(n13799), 
           .MB1(n13798), .MB0(n13797), .CIN53(n13868), .CIN52(n13867), 
           .CIN51(n13866), .CIN50(n13865), .CIN49(n13864), .CIN48(n13863), 
           .CIN47(n13862), .CIN46(n13861), .CIN45(n13860), .CIN44(n13859), 
           .CIN43(n13858), .CIN42(n13857), .CIN41(n13856), .CIN40(n13855), 
           .CIN39(n13854), .CIN38(n13853), .CIN37(n13852), .CIN36(n13851), 
           .CIN35(n13850), .CIN34(n13849), .CIN33(n13848), .CIN32(n13847), 
           .CIN31(n13846), .CIN30(n13845), .CIN29(n13844), .CIN28(n13843), 
           .CIN27(n13842), .CIN26(n13841), .CIN25(n13840), .CIN24(n13839), 
           .CIN23(n13838), .CIN22(n13837), .CIN21(n13836), .CIN20(n13835), 
           .CIN19(n13834), .CIN18(n13833), .CIN17(n8704), .CIN16(n8705), 
           .CIN15(n8706), .CIN14(n8707), .CIN13(n8708), .CIN12(n8709), 
           .CIN11(n8710), .CIN10(n8711), .CIN9(n8712), .CIN8(n8713), 
           .CIN7(n8714), .CIN6(n8715), .CIN5(n8716), .CIN4(n8717), .CIN3(n8718), 
           .CIN2(n8719), .CIN1(n8720), .CIN0(n8721), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R7(n8696), .R6(n8697), .R5(n8698), 
           .R4(n8699), .R3(n8700), .R2(n8701), .R1(n8702), .R0(n8703));
    defparam lat_alu_9.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_9.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_9.REG_FLAG_CLK = "NONE";
    defparam lat_alu_9.REG_FLAG_CE = "CE0";
    defparam lat_alu_9.REG_FLAG_RST = "RST0";
    defparam lat_alu_9.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASK01 = "0x00000000000000";
    defparam lat_alu_9.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_9.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_9.CLK0_DIV = "ENABLED";
    defparam lat_alu_9.CLK1_DIV = "ENABLED";
    defparam lat_alu_9.CLK2_DIV = "ENABLED";
    defparam lat_alu_9.CLK3_DIV = "ENABLED";
    defparam lat_alu_9.MCPAT = "0x00000000000000";
    defparam lat_alu_9.MASKPAT = "0x00000000000000";
    defparam lat_alu_9.RNDPAT = "0x00000000000000";
    defparam lat_alu_9.GSR = "DISABLED";
    defparam lat_alu_9.RESETMODE = "SYNC";
    defparam lat_alu_9.MULT9_MODE = "DISABLED";
    defparam lat_alu_9.LEGACY = "DISABLED";
    ALU54B lat_alu_8 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n13577), .SIGNEDIB(n13650), .SIGNEDCIN(GND_net), 
           .A35(n13576), .A34(n13575), .A33(n13574), .A32(n13573), .A31(n13572), 
           .A30(n13571), .A29(n13570), .A28(n13569), .A27(n13568), .A26(n13567), 
           .A25(n13566), .A24(n13565), .A23(n13564), .A22(n13563), .A21(n13562), 
           .A20(n13561), .A19(n13560), .A18(n13559), .A17(n13558), .A16(n13557), 
           .A15(n13556), .A14(n13555), .A13(n13554), .A12(n13553), .A11(n13552), 
           .A10(n13551), .A9(n13550), .A8(n13549), .A7(n13548), .A6(n13547), 
           .A5(n13546), .A4(n13545), .A3(n13544), .A2(n13543), .A1(n13542), 
           .A0(n13541), .B35(n13649), .B34(n13648), .B33(n13647), .B32(n13646), 
           .B31(n13645), .B30(n13644), .B29(n13643), .B28(n13642), .B27(n13641), 
           .B26(n13640), .B25(n13639), .B24(n13638), .B23(n13637), .B22(n13636), 
           .B21(n13635), .B20(n13634), .B19(n13633), .B18(n13632), .B17(n13631), 
           .B16(n13630), .B15(n13629), .B14(n13628), .B13(n13627), .B12(n13626), 
           .B11(n13625), .B10(n13624), .B9(n13623), .B8(n13622), .B7(n13621), 
           .B6(n13620), .B5(n13619), .B4(n13618), .B3(n13617), .B2(n13616), 
           .B1(n13615), .B0(n13614), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n13613), .MA34(n13612), .MA33(n13611), .MA32(n13610), 
           .MA31(n13609), .MA30(n13608), .MA29(n13607), .MA28(n13606), 
           .MA27(n13605), .MA26(n13604), .MA25(n13603), .MA24(n13602), 
           .MA23(n13601), .MA22(n13600), .MA21(n13599), .MA20(n13598), 
           .MA19(n13597), .MA18(n13596), .MA17(n13595), .MA16(n13594), 
           .MA15(n13593), .MA14(n13592), .MA13(n13591), .MA12(n13590), 
           .MA11(n13589), .MA10(n13588), .MA9(n13587), .MA8(n13586), 
           .MA7(n13585), .MA6(n13584), .MA5(n13583), .MA4(n13582), .MA3(n13581), 
           .MA2(n13580), .MA1(n13579), .MA0(n13578), .MB35(n13686), 
           .MB34(n13685), .MB33(n13684), .MB32(n13683), .MB31(n13682), 
           .MB30(n13681), .MB29(n13680), .MB28(n13679), .MB27(n13678), 
           .MB26(n13677), .MB25(n13676), .MB24(n13675), .MB23(n13674), 
           .MB22(n13673), .MB21(n13672), .MB20(n13671), .MB19(n13670), 
           .MB18(n13669), .MB17(n13668), .MB16(n13667), .MB15(n13666), 
           .MB14(n13665), .MB13(n13664), .MB12(n13663), .MB11(n13662), 
           .MB10(n13661), .MB9(n13660), .MB8(n13659), .MB7(n13658), 
           .MB6(n13657), .MB5(n13656), .MB4(n13655), .MB3(n13654), .MB2(n13653), 
           .MB1(n13652), .MB0(n13651), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n13868), 
           .R52(n13867), .R51(n13866), .R50(n13865), .R49(n13864), .R48(n13863), 
           .R47(n13862), .R46(n13861), .R45(n13860), .R44(n13859), .R43(n13858), 
           .R42(n13857), .R41(n13856), .R40(n13855), .R39(n13854), .R38(n13853), 
           .R37(n13852), .R36(n13851), .R35(n13850), .R34(n13849), .R33(n13848), 
           .R32(n13847), .R31(n13846), .R30(n13845), .R29(n13844), .R28(n13843), 
           .R27(n13842), .R26(n13841), .R25(n13840), .R24(n13839), .R23(n13838), 
           .R22(n13837), .R21(n13836), .R20(n13835), .R19(n13834), .R18(n13833), 
           .R17(n8704), .R16(n8705), .R15(n8706), .R14(n8707), .R13(n8708), 
           .R12(n8709), .R11(n8710), .R10(n8711), .R9(n8712), .R8(n8713), 
           .R7(n8714), .R6(n8715), .R5(n8716), .R4(n8717), .R3(n8718), 
           .R2(n8719), .R1(n8720), .R0(n8721), .SIGNEDR(n13869));
    defparam lat_alu_8.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_8.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_8.REG_FLAG_CLK = "NONE";
    defparam lat_alu_8.REG_FLAG_CE = "CE0";
    defparam lat_alu_8.REG_FLAG_RST = "RST0";
    defparam lat_alu_8.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASK01 = "0x00000000000000";
    defparam lat_alu_8.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_8.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_8.CLK0_DIV = "ENABLED";
    defparam lat_alu_8.CLK1_DIV = "ENABLED";
    defparam lat_alu_8.CLK2_DIV = "ENABLED";
    defparam lat_alu_8.CLK3_DIV = "ENABLED";
    defparam lat_alu_8.MCPAT = "0x00000000000000";
    defparam lat_alu_8.MASKPAT = "0x00000000000000";
    defparam lat_alu_8.RNDPAT = "0x00000000000000";
    defparam lat_alu_8.GSR = "DISABLED";
    defparam lat_alu_8.RESETMODE = "SYNC";
    defparam lat_alu_8.MULT9_MODE = "DISABLED";
    defparam lat_alu_8.LEGACY = "DISABLED";
    MULT18X18D lat_mult_7 (.A17(\rom8_w_i[12] ), .A16(\rom8_w_i[12] ), .A15(\rom8_w_i[12] ), 
            .A14(\rom8_w_i[12] ), .A13(\rom8_w_i[12] ), .A12(\rom8_w_i[12] ), 
            .A11(\rom8_w_i[12] ), .A10(\rom8_w_i[12] ), .A9(\rom8_w_i[12] ), 
            .A8(\rom8_w_i[12] ), .A7(\rom8_w_i[12] ), .A6(\rom8_w_i[12] ), 
            .A5(\rom8_w_i[12] ), .A4(\rom8_w_i[12] ), .A3(\rom8_w_i[12] ), 
            .A2(\rom8_w_i[12] ), .A1(\rom8_w_i[12] ), .A0(\rom8_w_i[12] ), 
            .B17(n319), .B16(n319), .B15(n319), .B14(n319), .B13(n319), 
            .B12(n319), .B11(n319), .B10(n319), .B9(n319), .B8(n319), 
            .B7(n319), .B6(n319), .B5(n319), .B4(n319), .B3(n319), 
            .B2(n319), .B1(n319), .B0(n319), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n13777), .ROA16(n13776), .ROA15(n13775), .ROA14(n13774), 
            .ROA13(n13773), .ROA12(n13772), .ROA11(n13771), .ROA10(n13770), 
            .ROA9(n13769), .ROA8(n13768), .ROA7(n13767), .ROA6(n13766), 
            .ROA5(n13765), .ROA4(n13764), .ROA3(n13763), .ROA2(n13762), 
            .ROA1(n13761), .ROA0(n13760), .ROB17(n13795), .ROB16(n13794), 
            .ROB15(n13793), .ROB14(n13792), .ROB13(n13791), .ROB12(n13790), 
            .ROB11(n13789), .ROB10(n13788), .ROB9(n13787), .ROB8(n13786), 
            .ROB7(n13785), .ROB6(n13784), .ROB5(n13783), .ROB4(n13782), 
            .ROB3(n13781), .ROB2(n13780), .ROB1(n13779), .ROB0(n13778), 
            .P35(n13832), .P34(n13831), .P33(n13830), .P32(n13829), 
            .P31(n13828), .P30(n13827), .P29(n13826), .P28(n13825), 
            .P27(n13824), .P26(n13823), .P25(n13822), .P24(n13821), 
            .P23(n13820), .P22(n13819), .P21(n13818), .P20(n13817), 
            .P19(n13816), .P18(n13815), .P17(n13814), .P16(n13813), 
            .P15(n13812), .P14(n13811), .P13(n13810), .P12(n13809), 
            .P11(n13808), .P10(n13807), .P9(n13806), .P8(n13805), .P7(n13804), 
            .P6(n13803), .P5(n13802), .P4(n13801), .P3(n13800), .P2(n13799), 
            .P1(n13798), .P0(n13797), .SIGNEDP(n13796));
    defparam lat_mult_7.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTA_CE = "CE0";
    defparam lat_mult_7.REG_INPUTA_RST = "RST0";
    defparam lat_mult_7.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTB_CE = "CE0";
    defparam lat_mult_7.REG_INPUTB_RST = "RST0";
    defparam lat_mult_7.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTC_CE = "CE0";
    defparam lat_mult_7.REG_INPUTC_RST = "RST0";
    defparam lat_mult_7.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_7.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_7.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_7.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_7.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_7.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_7.CLK0_DIV = "ENABLED";
    defparam lat_mult_7.CLK1_DIV = "ENABLED";
    defparam lat_mult_7.CLK2_DIV = "ENABLED";
    defparam lat_mult_7.CLK3_DIV = "ENABLED";
    defparam lat_mult_7.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_7.GSR = "DISABLED";
    defparam lat_mult_7.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_7.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_7.MULT_BYPASS = "DISABLED";
    defparam lat_mult_7.RESETMODE = "SYNC";
    MULT18X18D lat_mult_6 (.A17(\rom8_w_i[12] ), .A16(\rom8_w_i[12] ), .A15(\rom8_w_i[12] ), 
            .A14(\rom8_w_i[12] ), .A13(\rom8_w_i[12] ), .A12(\rom8_w_i[12] ), 
            .A11(\rom8_w_i[12] ), .A10(\rom8_w_i[12] ), .A9(\rom8_w_i[12] ), 
            .A8(\rom8_w_i[12] ), .A7(\rom8_w_i[2] ), .A6(\rom8_w_i[6] ), 
            .A5(GND_net), .A4(\rom8_w_i[4] ), .A3(\rom8_w_i[3] ), .A2(\rom8_w_i[2] ), 
            .A1(\rom8_w_i[1] ), .A0(\rom8_w_i[0] ), .B17(n319), .B16(n319), 
            .B15(n319), .B14(n319), .B13(n319), .B12(n319), .B11(n319), 
            .B10(n319), .B9(n319), .B8(n319), .B7(n319), .B6(n319), 
            .B5(n319), .B4(n319), .B3(n319), .B2(n319), .B1(n319), 
            .B0(n319), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n13704), 
            .ROA16(n13703), .ROA15(n13702), .ROA14(n13701), .ROA13(n13700), 
            .ROA12(n13699), .ROA11(n13698), .ROA10(n13697), .ROA9(n13696), 
            .ROA8(n13695), .ROA7(n13694), .ROA6(n13693), .ROA5(n13692), 
            .ROA4(n13691), .ROA3(n13690), .ROA2(n13689), .ROA1(n13688), 
            .ROA0(n13687), .ROB17(n13722), .ROB16(n13721), .ROB15(n13720), 
            .ROB14(n13719), .ROB13(n13718), .ROB12(n13717), .ROB11(n13716), 
            .ROB10(n13715), .ROB9(n13714), .ROB8(n13713), .ROB7(n13712), 
            .ROB6(n13711), .ROB5(n13710), .ROB4(n13709), .ROB3(n13708), 
            .ROB2(n13707), .ROB1(n13706), .ROB0(n13705), .P35(n13759), 
            .P34(n13758), .P33(n13757), .P32(n13756), .P31(n13755), 
            .P30(n13754), .P29(n13753), .P28(n13752), .P27(n13751), 
            .P26(n13750), .P25(n13749), .P24(n13748), .P23(n13747), 
            .P22(n13746), .P21(n13745), .P20(n13744), .P19(n13743), 
            .P18(n13742), .P17(n13741), .P16(n13740), .P15(n13739), 
            .P14(n13738), .P13(n13737), .P12(n13736), .P11(n13735), 
            .P10(n13734), .P9(n13733), .P8(n13732), .P7(n13731), .P6(n13730), 
            .P5(n13729), .P4(n13728), .P3(n13727), .P2(n13726), .P1(n13725), 
            .P0(n13724), .SIGNEDP(n13723));
    defparam lat_mult_6.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTA_CE = "CE0";
    defparam lat_mult_6.REG_INPUTA_RST = "RST0";
    defparam lat_mult_6.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTB_CE = "CE0";
    defparam lat_mult_6.REG_INPUTB_RST = "RST0";
    defparam lat_mult_6.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTC_CE = "CE0";
    defparam lat_mult_6.REG_INPUTC_RST = "RST0";
    defparam lat_mult_6.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_6.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_6.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_6.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_6.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_6.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_6.CLK0_DIV = "ENABLED";
    defparam lat_mult_6.CLK1_DIV = "ENABLED";
    defparam lat_mult_6.CLK2_DIV = "ENABLED";
    defparam lat_mult_6.CLK3_DIV = "ENABLED";
    defparam lat_mult_6.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_6.GSR = "DISABLED";
    defparam lat_mult_6.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_6.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_6.MULT_BYPASS = "DISABLED";
    defparam lat_mult_6.RESETMODE = "SYNC";
    MULT18X18D lat_mult_5 (.A17(\rom8_w_i[12] ), .A16(\rom8_w_i[12] ), .A15(\rom8_w_i[12] ), 
            .A14(\rom8_w_i[12] ), .A13(\rom8_w_i[12] ), .A12(\rom8_w_i[12] ), 
            .A11(\rom8_w_i[12] ), .A10(\rom8_w_i[12] ), .A9(\rom8_w_i[12] ), 
            .A8(\rom8_w_i[12] ), .A7(\rom8_w_i[12] ), .A6(\rom8_w_i[12] ), 
            .A5(\rom8_w_i[12] ), .A4(\rom8_w_i[12] ), .A3(\rom8_w_i[12] ), 
            .A2(\rom8_w_i[12] ), .A1(\rom8_w_i[12] ), .A0(\rom8_w_i[12] ), 
            .B17(n11171), .B16(n11170), .B15(n11169), .B14(n11168), 
            .B13(n11167), .B12(n11166), .B11(n11165), .B10(n11164), 
            .B9(n11163), .B8(n11162), .B7(n11161), .B6(n11160), .B5(n11159), 
            .B4(n11158), .B3(n11157), .B2(n11156), .B1(n11155), .B0(n11154), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n13631), .ROA16(n13630), 
            .ROA15(n13629), .ROA14(n13628), .ROA13(n13627), .ROA12(n13626), 
            .ROA11(n13625), .ROA10(n13624), .ROA9(n13623), .ROA8(n13622), 
            .ROA7(n13621), .ROA6(n13620), .ROA5(n13619), .ROA4(n13618), 
            .ROA3(n13617), .ROA2(n13616), .ROA1(n13615), .ROA0(n13614), 
            .ROB17(n13649), .ROB16(n13648), .ROB15(n13647), .ROB14(n13646), 
            .ROB13(n13645), .ROB12(n13644), .ROB11(n13643), .ROB10(n13642), 
            .ROB9(n13641), .ROB8(n13640), .ROB7(n13639), .ROB6(n13638), 
            .ROB5(n13637), .ROB4(n13636), .ROB3(n13635), .ROB2(n13634), 
            .ROB1(n13633), .ROB0(n13632), .P35(n13686), .P34(n13685), 
            .P33(n13684), .P32(n13683), .P31(n13682), .P30(n13681), 
            .P29(n13680), .P28(n13679), .P27(n13678), .P26(n13677), 
            .P25(n13676), .P24(n13675), .P23(n13674), .P22(n13673), 
            .P21(n13672), .P20(n13671), .P19(n13670), .P18(n13669), 
            .P17(n13668), .P16(n13667), .P15(n13666), .P14(n13665), 
            .P13(n13664), .P12(n13663), .P11(n13662), .P10(n13661), 
            .P9(n13660), .P8(n13659), .P7(n13658), .P6(n13657), .P5(n13656), 
            .P4(n13655), .P3(n13654), .P2(n13653), .P1(n13652), .P0(n13651), 
            .SIGNEDP(n13650));
    defparam lat_mult_5.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTA_CE = "CE0";
    defparam lat_mult_5.REG_INPUTA_RST = "RST0";
    defparam lat_mult_5.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTB_CE = "CE0";
    defparam lat_mult_5.REG_INPUTB_RST = "RST0";
    defparam lat_mult_5.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTC_CE = "CE0";
    defparam lat_mult_5.REG_INPUTC_RST = "RST0";
    defparam lat_mult_5.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_5.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_5.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_5.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_5.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_5.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_5.CLK0_DIV = "ENABLED";
    defparam lat_mult_5.CLK1_DIV = "ENABLED";
    defparam lat_mult_5.CLK2_DIV = "ENABLED";
    defparam lat_mult_5.CLK3_DIV = "ENABLED";
    defparam lat_mult_5.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_5.GSR = "DISABLED";
    defparam lat_mult_5.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_5.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_5.MULT_BYPASS = "DISABLED";
    defparam lat_mult_5.RESETMODE = "SYNC";
    MULT18X18D mult_969 (.A17(\rom8_w_i[12] ), .A16(\rom8_w_i[12] ), .A15(\rom8_w_i[12] ), 
            .A14(\rom8_w_i[12] ), .A13(\rom8_w_i[12] ), .A12(\rom8_w_i[12] ), 
            .A11(\rom8_w_i[12] ), .A10(\rom8_w_i[12] ), .A9(\rom8_w_i[12] ), 
            .A8(\rom8_w_i[12] ), .A7(\rom8_w_i[2] ), .A6(\rom8_w_i[6] ), 
            .A5(GND_net), .A4(\rom8_w_i[4] ), .A3(\rom8_w_i[3] ), .A2(\rom8_w_i[2] ), 
            .A1(\rom8_w_i[1] ), .A0(\rom8_w_i[0] ), .B17(n11171), .B16(n11170), 
            .B15(n11169), .B14(n11168), .B13(n11167), .B12(n11166), 
            .B11(n11165), .B10(n11164), .B9(n11163), .B8(n11162), .B7(n11161), 
            .B6(n11160), .B5(n11159), .B4(n11158), .B3(n11157), .B2(n11156), 
            .B1(n11155), .B0(n11154), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n13558), .ROA16(n13557), .ROA15(n13556), .ROA14(n13555), 
            .ROA13(n13554), .ROA12(n13553), .ROA11(n13552), .ROA10(n13551), 
            .ROA9(n13550), .ROA8(n13549), .ROA7(n13548), .ROA6(n13547), 
            .ROA5(n13546), .ROA4(n13545), .ROA3(n13544), .ROA2(n13543), 
            .ROA1(n13542), .ROA0(n13541), .ROB17(n13576), .ROB16(n13575), 
            .ROB15(n13574), .ROB14(n13573), .ROB13(n13572), .ROB12(n13571), 
            .ROB11(n13570), .ROB10(n13569), .ROB9(n13568), .ROB8(n13567), 
            .ROB7(n13566), .ROB6(n13565), .ROB5(n13564), .ROB4(n13563), 
            .ROB3(n13562), .ROB2(n13561), .ROB1(n13560), .ROB0(n13559), 
            .P35(n13613), .P34(n13612), .P33(n13611), .P32(n13610), 
            .P31(n13609), .P30(n13608), .P29(n13607), .P28(n13606), 
            .P27(n13605), .P26(n13604), .P25(n13603), .P24(n13602), 
            .P23(n13601), .P22(n13600), .P21(n13599), .P20(n13598), 
            .P19(n13597), .P18(n13596), .P17(n13595), .P16(n13594), 
            .P15(n13593), .P14(n13592), .P13(n13591), .P12(n13590), 
            .P11(n13589), .P10(n13588), .P9(n13587), .P8(n13586), .P7(n13585), 
            .P6(n13584), .P5(n13583), .P4(n13582), .P3(n13581), .P2(n13580), 
            .P1(n13579), .P0(n13578), .SIGNEDP(n13577));
    defparam mult_969.REG_INPUTA_CLK = "NONE";
    defparam mult_969.REG_INPUTA_CE = "CE0";
    defparam mult_969.REG_INPUTA_RST = "RST0";
    defparam mult_969.REG_INPUTB_CLK = "NONE";
    defparam mult_969.REG_INPUTB_CE = "CE0";
    defparam mult_969.REG_INPUTB_RST = "RST0";
    defparam mult_969.REG_INPUTC_CLK = "NONE";
    defparam mult_969.REG_INPUTC_CE = "CE0";
    defparam mult_969.REG_INPUTC_RST = "RST0";
    defparam mult_969.REG_PIPELINE_CLK = "NONE";
    defparam mult_969.REG_PIPELINE_CE = "CE0";
    defparam mult_969.REG_PIPELINE_RST = "RST0";
    defparam mult_969.REG_OUTPUT_CLK = "NONE";
    defparam mult_969.REG_OUTPUT_CE = "CE0";
    defparam mult_969.REG_OUTPUT_RST = "RST0";
    defparam mult_969.CLK0_DIV = "ENABLED";
    defparam mult_969.CLK1_DIV = "ENABLED";
    defparam mult_969.CLK2_DIV = "ENABLED";
    defparam mult_969.CLK3_DIV = "ENABLED";
    defparam mult_969.HIGHSPEED_CLK = "NONE";
    defparam mult_969.GSR = "DISABLED";
    defparam mult_969.CAS_MATCH_REG = "FALSE";
    defparam mult_969.SOURCEB_MODE = "B_SHIFT";
    defparam mult_969.MULT_BYPASS = "DISABLED";
    defparam mult_969.RESETMODE = "SYNC";
    MULT18X18D mult_8 (.A17(shift_8_dout_i[17]), .A16(shift_8_dout_i[16]), 
            .A15(shift_8_dout_i[15]), .A14(shift_8_dout_i[14]), .A13(shift_8_dout_i[13]), 
            .A12(shift_8_dout_i[12]), .A11(shift_8_dout_i[11]), .A10(shift_8_dout_i[10]), 
            .A9(shift_8_dout_i[9]), .A8(shift_8_dout_i[8]), .A7(shift_8_dout_i[7]), 
            .A6(shift_8_dout_i[6]), .A5(shift_8_dout_i[5]), .A4(shift_8_dout_i[4]), 
            .A3(shift_8_dout_i[3]), .A2(shift_8_dout_i[2]), .A1(shift_8_dout_i[1]), 
            .A0(shift_8_dout_i[0]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n12453), .B8(n12452), .B7(n12451), .B6(n12450), .B5(n12449), 
            .B4(n12448), .B3(n12447), .B2(n12446), .B1(n12445), .B0(n12444), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17415), .ROA16(n17414), 
            .ROA15(n17413), .ROA14(n17412), .ROA13(n17411), .ROA12(n17410), 
            .ROA11(n17409), .ROA10(n17408), .ROA9(n17407), .ROA8(n17406), 
            .ROA7(n17405), .ROA6(n17404), .ROA5(n17403), .ROA4(n17402), 
            .ROA3(n17401), .ROA2(n17400), .ROA1(n17399), .ROA0(n17398), 
            .ROB17(n17433), .ROB16(n17432), .ROB15(n17431), .ROB14(n17430), 
            .ROB13(n17429), .ROB12(n17428), .ROB11(n17427), .ROB10(n17426), 
            .ROB9(n17425), .ROB8(n17424), .ROB7(n17423), .ROB6(n17422), 
            .ROB5(n17421), .ROB4(n17420), .ROB3(n17419), .ROB2(n17418), 
            .ROB1(n17417), .ROB0(n17416), .P35(n17470), .P34(n17469), 
            .P33(n17468), .P32(n17467), .P31(n17466), .P30(n17465), 
            .P29(n17464), .P28(n17463), .P27(n17462), .P26(n17461), 
            .P25(n17460), .P24(n17459), .P23(n17458), .P22(n17457), 
            .P21(n17456), .P20(n17455), .P19(n17454), .P18(n17453), 
            .P17(n17452), .P16(n17451), .P15(n17450), .P14(n17449), 
            .P13(n17448), .P12(n17447), .P11(n17446), .P10(n17445), 
            .P9(n17444), .P8(n17443), .P7(n17442), .P6(n17441), .P5(n17440), 
            .P4(n17439), .P3(n17438), .P2(n17437), .P1(n17436), .P0(n17435), 
            .SIGNEDP(n17434));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam mult_8.REG_INPUTA_CLK = "NONE";
    defparam mult_8.REG_INPUTA_CE = "CE0";
    defparam mult_8.REG_INPUTA_RST = "RST0";
    defparam mult_8.REG_INPUTB_CLK = "NONE";
    defparam mult_8.REG_INPUTB_CE = "CE0";
    defparam mult_8.REG_INPUTB_RST = "RST0";
    defparam mult_8.REG_INPUTC_CLK = "NONE";
    defparam mult_8.REG_INPUTC_CE = "CE0";
    defparam mult_8.REG_INPUTC_RST = "RST0";
    defparam mult_8.REG_PIPELINE_CLK = "NONE";
    defparam mult_8.REG_PIPELINE_CE = "CE0";
    defparam mult_8.REG_PIPELINE_RST = "RST0";
    defparam mult_8.REG_OUTPUT_CLK = "NONE";
    defparam mult_8.REG_OUTPUT_CE = "CE0";
    defparam mult_8.REG_OUTPUT_RST = "RST0";
    defparam mult_8.CLK0_DIV = "ENABLED";
    defparam mult_8.CLK1_DIV = "ENABLED";
    defparam mult_8.CLK2_DIV = "ENABLED";
    defparam mult_8.CLK3_DIV = "ENABLED";
    defparam mult_8.HIGHSPEED_CLK = "NONE";
    defparam mult_8.GSR = "DISABLED";
    defparam mult_8.CAS_MATCH_REG = "FALSE";
    defparam mult_8.SOURCEB_MODE = "B_SHIFT";
    defparam mult_8.MULT_BYPASS = "DISABLED";
    defparam mult_8.RESETMODE = "SYNC";
    MULT18X18D lat_mult_60 (.A17(shift_8_dout_i[23]), .A16(shift_8_dout_i[23]), 
            .A15(shift_8_dout_i[23]), .A14(shift_8_dout_i[23]), .A13(shift_8_dout_i[23]), 
            .A12(shift_8_dout_i[23]), .A11(shift_8_dout_i[23]), .A10(shift_8_dout_i[23]), 
            .A9(shift_8_dout_i[23]), .A8(shift_8_dout_i[23]), .A7(shift_8_dout_i[23]), 
            .A6(shift_8_dout_i[23]), .A5(shift_8_dout_i[23]), .A4(shift_8_dout_i[22]), 
            .A3(shift_8_dout_i[21]), .A2(shift_8_dout_i[20]), .A1(shift_8_dout_i[19]), 
            .A0(shift_8_dout_i[18]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n12453), .B8(n12452), .B7(n12451), .B6(n12450), .B5(n12449), 
            .B4(n12448), .B3(n12447), .B2(n12446), .B1(n12445), .B0(n12444), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17488), .ROA16(n17487), 
            .ROA15(n17486), .ROA14(n17485), .ROA13(n17484), .ROA12(n17483), 
            .ROA11(n17482), .ROA10(n17481), .ROA9(n17480), .ROA8(n17479), 
            .ROA7(n17478), .ROA6(n17477), .ROA5(n17476), .ROA4(n17475), 
            .ROA3(n17474), .ROA2(n17473), .ROA1(n17472), .ROA0(n17471), 
            .ROB17(n17506), .ROB16(n17505), .ROB15(n17504), .ROB14(n17503), 
            .ROB13(n17502), .ROB12(n17501), .ROB11(n17500), .ROB10(n17499), 
            .ROB9(n17498), .ROB8(n17497), .ROB7(n17496), .ROB6(n17495), 
            .ROB5(n17494), .ROB4(n17493), .ROB3(n17492), .ROB2(n17491), 
            .ROB1(n17490), .ROB0(n17489), .P35(n17543), .P34(n17542), 
            .P33(n17541), .P32(n17540), .P31(n17539), .P30(n17538), 
            .P29(n17537), .P28(n17536), .P27(n17535), .P26(n17534), 
            .P25(n17533), .P24(n17532), .P23(n17531), .P22(n17530), 
            .P21(n17529), .P20(n17528), .P19(n17527), .P18(n17526), 
            .P17(n17525), .P16(n17524), .P15(n17523), .P14(n17522), 
            .P13(n17521), .P12(n17520), .P11(n17519), .P10(n17518), 
            .P9(n17517), .P8(n17516), .P7(n17515), .P6(n17514), .P5(n17513), 
            .P4(n17512), .P3(n17511), .P2(n17510), .P1(n17509), .P0(n17508), 
            .SIGNEDP(n17507));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_60.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_60.REG_INPUTA_CE = "CE0";
    defparam lat_mult_60.REG_INPUTA_RST = "RST0";
    defparam lat_mult_60.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_60.REG_INPUTB_CE = "CE0";
    defparam lat_mult_60.REG_INPUTB_RST = "RST0";
    defparam lat_mult_60.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_60.REG_INPUTC_CE = "CE0";
    defparam lat_mult_60.REG_INPUTC_RST = "RST0";
    defparam lat_mult_60.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_60.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_60.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_60.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_60.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_60.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_60.CLK0_DIV = "ENABLED";
    defparam lat_mult_60.CLK1_DIV = "ENABLED";
    defparam lat_mult_60.CLK2_DIV = "ENABLED";
    defparam lat_mult_60.CLK3_DIV = "ENABLED";
    defparam lat_mult_60.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_60.GSR = "DISABLED";
    defparam lat_mult_60.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_60.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_60.MULT_BYPASS = "DISABLED";
    defparam lat_mult_60.RESETMODE = "SYNC";
    MULT18X18D lat_mult_65 (.A17(\rom8_w_r[10] ), .A16(\rom8_w_r[10] ), 
            .A15(\rom8_w_r[10] ), .A14(\rom8_w_r[10] ), .A13(\rom8_w_r[10] ), 
            .A12(\rom8_w_r[10] ), .A11(\rom8_w_r[10] ), .A10(\rom8_w_r[10] ), 
            .A9(\rom8_w_r[10] ), .A8(\rom8_w_r[10] ), .A7(\rom8_w_r[10] ), 
            .A6(\rom8_w_r[10] ), .A5(\rom8_w_r[10] ), .A4(\rom8_w_r[10] ), 
            .A3(\rom8_w_r[10] ), .A2(\rom8_w_r[10] ), .A1(\rom8_w_r[10] ), 
            .A0(\rom8_w_r[10] ), .B17(n12287), .B16(n12286), .B15(n12285), 
            .B14(n12284), .B13(n12283), .B12(n12282), .B11(n12281), 
            .B10(n12280), .B9(n12279), .B8(n12278), .B7(n12277), .B6(n12276), 
            .B5(n12275), .B4(n12274), .B3(n12273), .B2(n12272), .B1(n12271), 
            .B0(n12270), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17834), 
            .ROA16(n17833), .ROA15(n17832), .ROA14(n17831), .ROA13(n17830), 
            .ROA12(n17829), .ROA11(n17828), .ROA10(n17827), .ROA9(n17826), 
            .ROA8(n17825), .ROA7(n17824), .ROA6(n17823), .ROA5(n17822), 
            .ROA4(n17821), .ROA3(n17820), .ROA2(n17819), .ROA1(n17818), 
            .ROA0(n17817), .ROB17(n17852), .ROB16(n17851), .ROB15(n17850), 
            .ROB14(n17849), .ROB13(n17848), .ROB12(n17847), .ROB11(n17846), 
            .ROB10(n17845), .ROB9(n17844), .ROB8(n17843), .ROB7(n17842), 
            .ROB6(n17841), .ROB5(n17840), .ROB4(n17839), .ROB3(n17838), 
            .ROB2(n17837), .ROB1(n17836), .ROB0(n17835), .P35(n17889), 
            .P34(n17888), .P33(n17887), .P32(n17886), .P31(n17885), 
            .P30(n17884), .P29(n17883), .P28(n17882), .P27(n17881), 
            .P26(n17880), .P25(n17879), .P24(n17878), .P23(n17877), 
            .P22(n17876), .P21(n17875), .P20(n17874), .P19(n17873), 
            .P18(n17872), .P17(n17871), .P16(n17870), .P15(n17869), 
            .P14(n17868), .P13(n17867), .P12(n17866), .P11(n17865), 
            .P10(n17864), .P9(n17863), .P8(n17862), .P7(n17861), .P6(n17860), 
            .P5(n17859), .P4(n17858), .P3(n17857), .P2(n17856), .P1(n17855), 
            .P0(n17854), .SIGNEDP(n17853));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_65.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_65.REG_INPUTA_CE = "CE0";
    defparam lat_mult_65.REG_INPUTA_RST = "RST0";
    defparam lat_mult_65.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_65.REG_INPUTB_CE = "CE0";
    defparam lat_mult_65.REG_INPUTB_RST = "RST0";
    defparam lat_mult_65.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_65.REG_INPUTC_CE = "CE0";
    defparam lat_mult_65.REG_INPUTC_RST = "RST0";
    defparam lat_mult_65.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_65.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_65.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_65.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_65.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_65.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_65.CLK0_DIV = "ENABLED";
    defparam lat_mult_65.CLK1_DIV = "ENABLED";
    defparam lat_mult_65.CLK2_DIV = "ENABLED";
    defparam lat_mult_65.CLK3_DIV = "ENABLED";
    defparam lat_mult_65.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_65.GSR = "DISABLED";
    defparam lat_mult_65.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_65.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_65.MULT_BYPASS = "DISABLED";
    defparam lat_mult_65.RESETMODE = "SYNC";
    MULT18X18D lat_mult_66 (.A17(\rom8_w_r[10] ), .A16(\rom8_w_r[10] ), 
            .A15(\rom8_w_r[10] ), .A14(\rom8_w_r[10] ), .A13(\rom8_w_r[10] ), 
            .A12(\rom8_w_r[10] ), .A11(\rom8_w_r[10] ), .A10(\rom8_w_r[10] ), 
            .A9(\rom8_w_r[10] ), .A8(\rom8_w_r[8] ), .A7(\rom8_w_r[7] ), 
            .A6(\rom8_w_r[6] ), .A5(\rom8_w_r[5] ), .A4(\rom8_w_r[4] ), 
            .A3(\rom8_w_r[3] ), .A2(\rom8_w_r[7] ), .A1(\rom8_w_r[1] ), 
            .A0(\rom8_w_r[0] ), .B17(n12294), .B16(n12294), .B15(n12294), 
            .B14(n12294), .B13(n12294), .B12(n12294), .B11(n12294), 
            .B10(n12294), .B9(n12294), .B8(n12294), .B7(n12294), .B6(n12294), 
            .B5(n12293), .B4(n12292), .B3(n12291), .B2(n12290), .B1(n12289), 
            .B0(n12288), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17907), 
            .ROA16(n17906), .ROA15(n17905), .ROA14(n17904), .ROA13(n17903), 
            .ROA12(n17902), .ROA11(n17901), .ROA10(n17900), .ROA9(n17899), 
            .ROA8(n17898), .ROA7(n17897), .ROA6(n17896), .ROA5(n17895), 
            .ROA4(n17894), .ROA3(n17893), .ROA2(n17892), .ROA1(n17891), 
            .ROA0(n17890), .ROB17(n17925), .ROB16(n17924), .ROB15(n17923), 
            .ROB14(n17922), .ROB13(n17921), .ROB12(n17920), .ROB11(n17919), 
            .ROB10(n17918), .ROB9(n17917), .ROB8(n17916), .ROB7(n17915), 
            .ROB6(n17914), .ROB5(n17913), .ROB4(n17912), .ROB3(n17911), 
            .ROB2(n17910), .ROB1(n17909), .ROB0(n17908), .P35(n17962), 
            .P34(n17961), .P33(n17960), .P32(n17959), .P31(n17958), 
            .P30(n17957), .P29(n17956), .P28(n17955), .P27(n17954), 
            .P26(n17953), .P25(n17952), .P24(n17951), .P23(n17950), 
            .P22(n17949), .P21(n17948), .P20(n17947), .P19(n17946), 
            .P18(n17945), .P17(n17944), .P16(n17943), .P15(n17942), 
            .P14(n17941), .P13(n17940), .P12(n17939), .P11(n17938), 
            .P10(n17937), .P9(n17936), .P8(n17935), .P7(n17934), .P6(n17933), 
            .P5(n17932), .P4(n17931), .P3(n17930), .P2(n17929), .P1(n17928), 
            .P0(n17927), .SIGNEDP(n17926));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_66.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_66.REG_INPUTA_CE = "CE0";
    defparam lat_mult_66.REG_INPUTA_RST = "RST0";
    defparam lat_mult_66.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_66.REG_INPUTB_CE = "CE0";
    defparam lat_mult_66.REG_INPUTB_RST = "RST0";
    defparam lat_mult_66.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_66.REG_INPUTC_CE = "CE0";
    defparam lat_mult_66.REG_INPUTC_RST = "RST0";
    defparam lat_mult_66.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_66.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_66.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_66.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_66.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_66.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_66.CLK0_DIV = "ENABLED";
    defparam lat_mult_66.CLK1_DIV = "ENABLED";
    defparam lat_mult_66.CLK2_DIV = "ENABLED";
    defparam lat_mult_66.CLK3_DIV = "ENABLED";
    defparam lat_mult_66.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_66.GSR = "DISABLED";
    defparam lat_mult_66.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_66.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_66.MULT_BYPASS = "DISABLED";
    defparam lat_mult_66.RESETMODE = "SYNC";
    MULT18X18D lat_mult_67 (.A17(\rom8_w_r[10] ), .A16(\rom8_w_r[10] ), 
            .A15(\rom8_w_r[10] ), .A14(\rom8_w_r[10] ), .A13(\rom8_w_r[10] ), 
            .A12(\rom8_w_r[10] ), .A11(\rom8_w_r[10] ), .A10(\rom8_w_r[10] ), 
            .A9(\rom8_w_r[10] ), .A8(\rom8_w_r[10] ), .A7(\rom8_w_r[10] ), 
            .A6(\rom8_w_r[10] ), .A5(\rom8_w_r[10] ), .A4(\rom8_w_r[10] ), 
            .A3(\rom8_w_r[10] ), .A2(\rom8_w_r[10] ), .A1(\rom8_w_r[10] ), 
            .A0(\rom8_w_r[10] ), .B17(n12294), .B16(n12294), .B15(n12294), 
            .B14(n12294), .B13(n12294), .B12(n12294), .B11(n12294), 
            .B10(n12294), .B9(n12294), .B8(n12294), .B7(n12294), .B6(n12294), 
            .B5(n12293), .B4(n12292), .B3(n12291), .B2(n12290), .B1(n12289), 
            .B0(n12288), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17980), 
            .ROA16(n17979), .ROA15(n17978), .ROA14(n17977), .ROA13(n17976), 
            .ROA12(n17975), .ROA11(n17974), .ROA10(n17973), .ROA9(n17972), 
            .ROA8(n17971), .ROA7(n17970), .ROA6(n17969), .ROA5(n17968), 
            .ROA4(n17967), .ROA3(n17966), .ROA2(n17965), .ROA1(n17964), 
            .ROA0(n17963), .ROB17(n17998), .ROB16(n17997), .ROB15(n17996), 
            .ROB14(n17995), .ROB13(n17994), .ROB12(n17993), .ROB11(n17992), 
            .ROB10(n17991), .ROB9(n17990), .ROB8(n17989), .ROB7(n17988), 
            .ROB6(n17987), .ROB5(n17986), .ROB4(n17985), .ROB3(n17984), 
            .ROB2(n17983), .ROB1(n17982), .ROB0(n17981), .P35(n18035), 
            .P34(n18034), .P33(n18033), .P32(n18032), .P31(n18031), 
            .P30(n18030), .P29(n18029), .P28(n18028), .P27(n18027), 
            .P26(n18026), .P25(n18025), .P24(n18024), .P23(n18023), 
            .P22(n18022), .P21(n18021), .P20(n18020), .P19(n18019), 
            .P18(n18018), .P17(n18017), .P16(n18016), .P15(n18015), 
            .P14(n18014), .P13(n18013), .P12(n18012), .P11(n18011), 
            .P10(n18010), .P9(n18009), .P8(n18008), .P7(n18007), .P6(n18006), 
            .P5(n18005), .P4(n18004), .P3(n18003), .P2(n18002), .P1(n18001), 
            .P0(n18000), .SIGNEDP(n17999));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_67.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_67.REG_INPUTA_CE = "CE0";
    defparam lat_mult_67.REG_INPUTA_RST = "RST0";
    defparam lat_mult_67.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_67.REG_INPUTB_CE = "CE0";
    defparam lat_mult_67.REG_INPUTB_RST = "RST0";
    defparam lat_mult_67.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_67.REG_INPUTC_CE = "CE0";
    defparam lat_mult_67.REG_INPUTC_RST = "RST0";
    defparam lat_mult_67.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_67.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_67.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_67.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_67.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_67.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_67.CLK0_DIV = "ENABLED";
    defparam lat_mult_67.CLK1_DIV = "ENABLED";
    defparam lat_mult_67.CLK2_DIV = "ENABLED";
    defparam lat_mult_67.CLK3_DIV = "ENABLED";
    defparam lat_mult_67.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_67.GSR = "DISABLED";
    defparam lat_mult_67.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_67.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_67.MULT_BYPASS = "DISABLED";
    defparam lat_mult_67.RESETMODE = "SYNC";
    ALU54B lat_alu_68 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n17780), .SIGNEDIB(n17853), .SIGNEDCIN(GND_net), 
           .A35(n17779), .A34(n17778), .A33(n17777), .A32(n17776), .A31(n17775), 
           .A30(n17774), .A29(n17773), .A28(n17772), .A27(n17771), .A26(n17770), 
           .A25(n17769), .A24(n17768), .A23(n17767), .A22(n17766), .A21(n17765), 
           .A20(n17764), .A19(n17763), .A18(n17762), .A17(n17761), .A16(n17760), 
           .A15(n17759), .A14(n17758), .A13(n17757), .A12(n17756), .A11(n17755), 
           .A10(n17754), .A9(n17753), .A8(n17752), .A7(n17751), .A6(n17750), 
           .A5(n17749), .A4(n17748), .A3(n17747), .A2(n17746), .A1(n17745), 
           .A0(n17744), .B35(n17852), .B34(n17851), .B33(n17850), .B32(n17849), 
           .B31(n17848), .B30(n17847), .B29(n17846), .B28(n17845), .B27(n17844), 
           .B26(n17843), .B25(n17842), .B24(n17841), .B23(n17840), .B22(n17839), 
           .B21(n17838), .B20(n17837), .B19(n17836), .B18(n17835), .B17(n17834), 
           .B16(n17833), .B15(n17832), .B14(n17831), .B13(n17830), .B12(n17829), 
           .B11(n17828), .B10(n17827), .B9(n17826), .B8(n17825), .B7(n17824), 
           .B6(n17823), .B5(n17822), .B4(n17821), .B3(n17820), .B2(n17819), 
           .B1(n17818), .B0(n17817), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n17816), .MA34(n17815), .MA33(n17814), .MA32(n17813), 
           .MA31(n17812), .MA30(n17811), .MA29(n17810), .MA28(n17809), 
           .MA27(n17808), .MA26(n17807), .MA25(n17806), .MA24(n17805), 
           .MA23(n17804), .MA22(n17803), .MA21(n17802), .MA20(n17801), 
           .MA19(n17800), .MA18(n17799), .MA17(n17798), .MA16(n17797), 
           .MA15(n17796), .MA14(n17795), .MA13(n17794), .MA12(n17793), 
           .MA11(n17792), .MA10(n17791), .MA9(n17790), .MA8(n17789), 
           .MA7(n17788), .MA6(n17787), .MA5(n17786), .MA4(n17785), .MA3(n17784), 
           .MA2(n17783), .MA1(n17782), .MA0(n17781), .MB35(n17889), 
           .MB34(n17888), .MB33(n17887), .MB32(n17886), .MB31(n17885), 
           .MB30(n17884), .MB29(n17883), .MB28(n17882), .MB27(n17881), 
           .MB26(n17880), .MB25(n17879), .MB24(n17878), .MB23(n17877), 
           .MB22(n17876), .MB21(n17875), .MB20(n17874), .MB19(n17873), 
           .MB18(n17872), .MB17(n17871), .MB16(n17870), .MB15(n17869), 
           .MB14(n17868), .MB13(n17867), .MB12(n17866), .MB11(n17865), 
           .MB10(n17864), .MB9(n17863), .MB8(n17862), .MB7(n17861), 
           .MB6(n17860), .MB5(n17859), .MB4(n17858), .MB3(n17857), .MB2(n17856), 
           .MB1(n17855), .MB0(n17854), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n18071), 
           .R52(n18070), .R51(n18069), .R50(n18068), .R49(n18067), .R48(n18066), 
           .R47(n18065), .R46(n18064), .R45(n18063), .R44(n18062), .R43(n18061), 
           .R42(n18060), .R41(n18059), .R40(n18058), .R39(n18057), .R38(n18056), 
           .R37(n18055), .R36(n18054), .R35(n18053), .R34(n18052), .R33(n18051), 
           .R32(n18050), .R31(n18049), .R30(n18048), .R29(n18047), .R28(n18046), 
           .R27(n18045), .R26(n18044), .R25(n18043), .R24(n18042), .R23(n18041), 
           .R22(n18040), .R21(n18039), .R20(n18038), .R19(n18037), .R18(n18036), 
           .R17(\op_r_23__N_1226[17] ), .R16(\op_r_23__N_1226[16] ), .R15(\op_r_23__N_1226[15] ), 
           .R14(\op_r_23__N_1226[14] ), .R13(\op_r_23__N_1226[13] ), .R12(\op_r_23__N_1226[12] ), 
           .R11(\op_r_23__N_1226[11] ), .R10(\op_r_23__N_1226[10] ), .R9(\op_r_23__N_1226[9] ), 
           .R8(\op_r_23__N_1226[8] ), .R7(\op_r_23__N_1226[7] ), .R6(\op_r_23__N_1226[6] ), 
           .R5(\op_r_23__N_1226[5] ), .R4(\op_r_23__N_1226[4] ), .R3(\op_r_23__N_1226[3] ), 
           .R2(\op_r_23__N_1226[2] ), .R1(\op_r_23__N_1226[1] ), .R0(\op_r_23__N_1226[0] ), 
           .SIGNEDR(n18072));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_68.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_68.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_68.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_68.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_68.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_68.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_68.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_68.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_68.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_68.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_68.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_68.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_68.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_68.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_68.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_68.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_68.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_68.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_68.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_68.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_68.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_68.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_68.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_68.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_68.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_68.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_68.REG_FLAG_CLK = "NONE";
    defparam lat_alu_68.REG_FLAG_CE = "CE0";
    defparam lat_alu_68.REG_FLAG_RST = "RST0";
    defparam lat_alu_68.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_68.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_68.MASK01 = "0x00000000000000";
    defparam lat_alu_68.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_68.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_68.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_68.CLK0_DIV = "ENABLED";
    defparam lat_alu_68.CLK1_DIV = "ENABLED";
    defparam lat_alu_68.CLK2_DIV = "ENABLED";
    defparam lat_alu_68.CLK3_DIV = "ENABLED";
    defparam lat_alu_68.MCPAT = "0x00000000000000";
    defparam lat_alu_68.MASKPAT = "0x00000000000000";
    defparam lat_alu_68.RNDPAT = "0x00000000000000";
    defparam lat_alu_68.GSR = "DISABLED";
    defparam lat_alu_68.RESETMODE = "SYNC";
    defparam lat_alu_68.MULT9_MODE = "DISABLED";
    defparam lat_alu_68.LEGACY = "DISABLED";
    LUT4 i13741_3_lut_4_lut (.A(op_i_23__N_1154[17]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[25] ), .Z(n31486)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13741_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i21_3_lut_4_lut (.A(op_r_23__N_1106[20]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[20]), .Z(n7431[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i21_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_391_i17_3_lut_4_lut (.A(op_r_23__N_1106[16]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[16]), .Z(n7431[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13694_3_lut_4_lut (.A(op_r_23__N_1106[16]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[24] ), .Z(n31439)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13694_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i18_3_lut_4_lut (.A(op_r_23__N_1106[17]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[17]), .Z(n7431[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i18_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13692_3_lut_4_lut (.A(op_r_23__N_1106[17]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[25] ), .Z(n31437)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13692_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i15_3_lut_4_lut (.A(op_i_23__N_1154[14]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[14]), .Z(n7590[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i15_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13747_3_lut_4_lut (.A(op_i_23__N_1154[14]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[22] ), .Z(n31492)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13747_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i16_3_lut_4_lut (.A(op_i_23__N_1154[15]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[15]), .Z(n7590[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i16_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13745_3_lut_4_lut (.A(op_i_23__N_1154[15]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[23] ), .Z(n31490)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13745_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i15_3_lut_4_lut (.A(op_r_23__N_1106[14]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[14]), .Z(n7431[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i15_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13698_3_lut_4_lut (.A(op_r_23__N_1106[14]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[22] ), .Z(n31443)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13698_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i16_3_lut_4_lut (.A(op_r_23__N_1106[15]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[15]), .Z(n7431[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i16_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13696_3_lut_4_lut (.A(op_r_23__N_1106[15]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[23] ), .Z(n31441)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13696_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i13_3_lut_4_lut (.A(op_i_23__N_1154[12]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[12]), .Z(n7590[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13751_3_lut_4_lut (.A(op_i_23__N_1154[12]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[20] ), .Z(n31496)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13751_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i14_3_lut_4_lut (.A(op_i_23__N_1154[13]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[13]), .Z(n7590[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i14_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13749_3_lut_4_lut (.A(op_i_23__N_1154[13]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[21] ), .Z(n31494)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13749_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i24_3_lut_4_lut (.A(op_i_23__N_1154[23]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[23]), .Z(n7590[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i24_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_391_i13_3_lut_4_lut (.A(op_r_23__N_1106[12]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[12]), .Z(n7431[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13702_3_lut_4_lut (.A(op_r_23__N_1106[12]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[20] ), .Z(n31447)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13702_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i14_3_lut_4_lut (.A(op_r_23__N_1106[13]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[13]), .Z(n7431[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i14_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13700_3_lut_4_lut (.A(op_r_23__N_1106[13]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[21] ), .Z(n31445)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13700_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i11_3_lut_4_lut (.A(op_i_23__N_1154[10]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[10]), .Z(n7590[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i11_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13755_3_lut_4_lut (.A(op_i_23__N_1154[10]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[18] ), .Z(n31500)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13755_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i12_3_lut_4_lut (.A(op_i_23__N_1154[11]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[11]), .Z(n7590[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i12_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13753_3_lut_4_lut (.A(op_i_23__N_1154[11]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[19] ), .Z(n31498)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13753_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i11_3_lut_4_lut (.A(op_r_23__N_1106[10]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[10]), .Z(n7431[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i11_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13706_3_lut_4_lut (.A(op_r_23__N_1106[10]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[18] ), .Z(n31451)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13706_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i12_3_lut_4_lut (.A(op_r_23__N_1106[11]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[11]), .Z(n7431[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i12_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13704_3_lut_4_lut (.A(op_r_23__N_1106[11]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[19] ), .Z(n31449)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13704_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i9_3_lut_4_lut (.A(op_i_23__N_1154[8]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[8]), .Z(n7590[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13759_3_lut_4_lut (.A(op_i_23__N_1154[8]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[16] ), .Z(n31504)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13759_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i10_3_lut_4_lut (.A(op_i_23__N_1154[9]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[9]), .Z(n7590[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13757_3_lut_4_lut (.A(op_i_23__N_1154[9]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[17] ), .Z(n31502)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13757_3_lut_4_lut.init = 16'hf808;
    LUT4 i13729_3_lut_4_lut (.A(op_i_23__N_1154[23]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[31] ), .Z(n31474)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13729_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i9_3_lut_4_lut (.A(op_r_23__N_1106[8]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[8]), .Z(n7431[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13710_3_lut_4_lut (.A(op_r_23__N_1106[8]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[16] ), .Z(n31455)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13710_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i10_3_lut_4_lut (.A(op_r_23__N_1106[9]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[9]), .Z(n7431[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_403_i23_3_lut_4_lut (.A(op_i_23__N_1154[22]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[22]), .Z(n7590[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i23_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13708_3_lut_4_lut (.A(op_r_23__N_1106[9]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[17] ), .Z(n31453)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13708_3_lut_4_lut.init = 16'hf808;
    LUT4 i13682_3_lut_4_lut (.A(op_r_23__N_1106[22]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[30] ), .Z(n31427)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13682_3_lut_4_lut.init = 16'hf808;
    LUT4 i13731_3_lut_4_lut (.A(op_i_23__N_1154[22]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[30] ), .Z(n31476)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13731_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i24_3_lut_4_lut (.A(op_r_23__N_1106[23]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[23]), .Z(n7431[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i24_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13680_3_lut_4_lut (.A(op_r_23__N_1106[23]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[31] ), .Z(n31425)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13680_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i23_3_lut_4_lut (.A(op_r_23__N_1106[22]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[22]), .Z(n7431[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i23_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_395_i2_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[1] ), 
         .D(shift_8_dout_i[1]), .Z(n7507)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i1_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[0] ), 
         .D(shift_8_dout_i[0]), .Z(n7508)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i4_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[3] ), 
         .D(shift_8_dout_i[3]), .Z(n7505)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i3_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[2] ), 
         .D(shift_8_dout_i[2]), .Z(n7506)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i6_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[5] ), 
         .D(shift_8_dout_i[5]), .Z(n7503)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i5_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[4] ), 
         .D(shift_8_dout_i[4]), .Z(n7504)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i8_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[7] ), 
         .D(shift_8_dout_i[7]), .Z(n7501)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_395_i7_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_i[6] ), 
         .D(shift_8_dout_i[6]), .Z(n7502)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_395_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i2_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[1] ), 
         .D(\shift_8_dout_r[1] ), .Z(n7560)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i1_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[0] ), 
         .D(\shift_8_dout_r[0] ), .Z(n7561)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i4_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[3] ), 
         .D(\shift_8_dout_r[3] ), .Z(n7558)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i3_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[2] ), 
         .D(\shift_8_dout_r[2] ), .Z(n7559)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i6_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[5] ), 
         .D(\shift_8_dout_r[5] ), .Z(n7556)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i5_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[4] ), 
         .D(\shift_8_dout_r[4] ), .Z(n7557)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i8_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[7] ), 
         .D(\shift_8_dout_r[7] ), .Z(n7554)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_399_i7_3_lut_4_lut (.A(\rom8_state[0] ), .B(n34794), .C(\radix_no1_op_r[6] ), 
         .D(\shift_8_dout_r[6] ), .Z(n7555)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_399_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i13677_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[8] ), 
         .D(\radix_no1_op_i[0] ), .Z(n31422)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13677_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13675_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[9] ), 
         .D(\radix_no1_op_i[1] ), .Z(n31420)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13675_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13667_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[13] ), 
         .D(\radix_no1_op_i[5] ), .Z(n31412)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13667_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13673_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[10] ), 
         .D(\radix_no1_op_i[2] ), .Z(n31418)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13673_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13671_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[11] ), 
         .D(\radix_no1_op_i[3] ), .Z(n31416)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13671_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13665_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[14] ), 
         .D(\radix_no1_op_i[6] ), .Z(n31410)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13665_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13663_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[15] ), 
         .D(\radix_no1_op_i[7] ), .Z(n31408)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13663_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13669_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_i_23__N_1130[12] ), 
         .D(\radix_no1_op_i[4] ), .Z(n31414)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13669_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13861_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[14] ), 
         .D(\radix_no1_op_r[6] ), .Z(n31606)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13861_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13859_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[15] ), 
         .D(\radix_no1_op_r[7] ), .Z(n31604)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13859_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13865_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[12] ), 
         .D(\radix_no1_op_r[4] ), .Z(n31610)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13865_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13863_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[13] ), 
         .D(\radix_no1_op_r[5] ), .Z(n31608)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13863_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13869_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[10] ), 
         .D(\radix_no1_op_r[2] ), .Z(n31614)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13869_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13867_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[11] ), 
         .D(\radix_no1_op_r[3] ), .Z(n31612)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13867_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13873_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[8] ), 
         .D(\radix_no1_op_r[0] ), .Z(n31618)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13873_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13871_3_lut_4_lut (.A(n34794), .B(\rom8_state[0] ), .C(\op_r_23__N_1082[9] ), 
         .D(\radix_no1_op_r[1] ), .Z(n31616)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13871_3_lut_4_lut.init = 16'hfd20;
    LUT4 i12907_2_lut_rep_263_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[14]), 
         .Z(n34625)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12907_2_lut_rep_263_3_lut.init = 16'h6060;
    LUT4 i12887_2_lut_rep_258_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[17]), 
         .Z(n34620)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12887_2_lut_rep_258_3_lut.init = 16'h6060;
    LUT4 i12886_2_lut_rep_257_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[16]), 
         .Z(n34619)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12886_2_lut_rep_257_3_lut.init = 16'h6060;
    LUT4 i12910_2_lut_rep_252_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[17]), 
         .Z(n34614)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12910_2_lut_rep_252_3_lut.init = 16'h6060;
    LUT4 i12909_2_lut_rep_251_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[16]), 
         .Z(n34613)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12909_2_lut_rep_251_3_lut.init = 16'h6060;
    LUT4 i12889_2_lut_rep_246_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[19]), 
         .Z(n34608)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12889_2_lut_rep_246_3_lut.init = 16'h6060;
    LUT4 i12888_2_lut_rep_245_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[18]), 
         .Z(n34607)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12888_2_lut_rep_245_3_lut.init = 16'h6060;
    LUT4 i12912_2_lut_rep_244_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[19]), 
         .Z(n34606)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12912_2_lut_rep_244_3_lut.init = 16'h6060;
    LUT4 i12911_2_lut_rep_243_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[18]), 
         .Z(n34605)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12911_2_lut_rep_243_3_lut.init = 16'h6060;
    LUT4 i12891_2_lut_rep_238_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[21]), 
         .Z(n34600)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12891_2_lut_rep_238_3_lut.init = 16'h6060;
    LUT4 i12890_2_lut_rep_237_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[20]), 
         .Z(n34599)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12890_2_lut_rep_237_3_lut.init = 16'h6060;
    LUT4 i12913_2_lut_rep_236_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[20]), 
         .Z(n34598)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12913_2_lut_rep_236_3_lut.init = 16'h6060;
    LUT4 i12914_2_lut_rep_235_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[21]), 
         .Z(n34597)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12914_2_lut_rep_235_3_lut.init = 16'h6060;
    LUT4 i12893_2_lut_rep_230_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[23]), 
         .Z(n34592)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12893_2_lut_rep_230_3_lut.init = 16'h6060;
    LUT4 i12892_2_lut_rep_229_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[22]), 
         .Z(n34591)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12892_2_lut_rep_229_3_lut.init = 16'h6060;
    LUT4 i12915_2_lut_rep_228_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[22]), 
         .Z(n34590)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12915_2_lut_rep_228_3_lut.init = 16'h6060;
    LUT4 i12916_2_lut_rep_227_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[23]), 
         .Z(n34589)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12916_2_lut_rep_227_3_lut.init = 16'h6060;
    LUT4 i12908_2_lut_rep_264_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[15]), 
         .Z(n34626)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12908_2_lut_rep_264_3_lut.init = 16'h6060;
    LUT4 i12884_2_lut_rep_269_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[14]), 
         .Z(n34631)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12884_2_lut_rep_269_3_lut.init = 16'h6060;
    LUT4 i12885_2_lut_rep_270_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[15]), 
         .Z(n34632)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12885_2_lut_rep_270_3_lut.init = 16'h6060;
    LUT4 i12905_2_lut_rep_275_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[12]), 
         .Z(n34637)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12905_2_lut_rep_275_3_lut.init = 16'h6060;
    LUT4 i12906_2_lut_rep_276_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[13]), 
         .Z(n34638)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12906_2_lut_rep_276_3_lut.init = 16'h6060;
    LUT4 i12882_2_lut_rep_281_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[12]), 
         .Z(n34643)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12882_2_lut_rep_281_3_lut.init = 16'h6060;
    LUT4 i12883_2_lut_rep_282_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[13]), 
         .Z(n34644)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12883_2_lut_rep_282_3_lut.init = 16'h6060;
    LUT4 i12903_2_lut_rep_285_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[10]), 
         .Z(n34647)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12903_2_lut_rep_285_3_lut.init = 16'h6060;
    LUT4 i12904_2_lut_rep_286_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[11]), 
         .Z(n34648)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12904_2_lut_rep_286_3_lut.init = 16'h6060;
    LUT4 i12880_2_lut_rep_291_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[10]), 
         .Z(n34653)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12880_2_lut_rep_291_3_lut.init = 16'h6060;
    LUT4 i12881_2_lut_rep_292_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[11]), 
         .Z(n34654)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12881_2_lut_rep_292_3_lut.init = 16'h6060;
    LUT4 i12901_2_lut_rep_295_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[8]), 
         .Z(n34657)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12901_2_lut_rep_295_3_lut.init = 16'h6060;
    LUT4 i12902_2_lut_rep_296_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[9]), 
         .Z(n34658)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12902_2_lut_rep_296_3_lut.init = 16'h6060;
    LUT4 i12878_2_lut_rep_301_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[8]), 
         .Z(n34663)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12878_2_lut_rep_301_3_lut.init = 16'h6060;
    LUT4 i12879_2_lut_rep_302_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[9]), 
         .Z(n34664)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12879_2_lut_rep_302_3_lut.init = 16'h6060;
    LUT4 i12899_2_lut_rep_319_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[6]), 
         .Z(n34681)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12899_2_lut_rep_319_3_lut.init = 16'h6060;
    LUT4 i12900_2_lut_rep_320_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[7]), 
         .Z(n34682)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12900_2_lut_rep_320_3_lut.init = 16'h6060;
    LUT4 i12876_2_lut_rep_325_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[6]), 
         .Z(n34687)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12876_2_lut_rep_325_3_lut.init = 16'h6060;
    LUT4 i12877_2_lut_rep_326_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[7]), 
         .Z(n34688)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12877_2_lut_rep_326_3_lut.init = 16'h6060;
    LUT4 i12898_2_lut_rep_329_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[5]), 
         .Z(n34691)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12898_2_lut_rep_329_3_lut.init = 16'h6060;
    LUT4 i12874_2_lut_rep_330_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[4]), 
         .Z(n34692)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12874_2_lut_rep_330_3_lut.init = 16'h6060;
    LUT4 i12875_2_lut_rep_331_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[5]), 
         .Z(n34693)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12875_2_lut_rep_331_3_lut.init = 16'h6060;
    LUT4 i12897_2_lut_rep_332_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[4]), 
         .Z(n34694)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12897_2_lut_rep_332_3_lut.init = 16'h6060;
    LUT4 i12872_2_lut_rep_333_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[2]), 
         .Z(n34695)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12872_2_lut_rep_333_3_lut.init = 16'h6060;
    LUT4 i12873_2_lut_rep_334_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[3]), 
         .Z(n34696)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12873_2_lut_rep_334_3_lut.init = 16'h6060;
    LUT4 i12895_2_lut_rep_335_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[2]), 
         .Z(n34697)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12895_2_lut_rep_335_3_lut.init = 16'h6060;
    LUT4 i12896_2_lut_rep_336_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[3]), 
         .Z(n34698)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12896_2_lut_rep_336_3_lut.init = 16'h6060;
    LUT4 i12550_2_lut_rep_337_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[0]), 
         .Z(n34699)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12550_2_lut_rep_337_3_lut.init = 16'h6060;
    LUT4 i12871_2_lut_rep_338_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_r_23__N_1106[1]), 
         .Z(n34700)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12871_2_lut_rep_338_3_lut.init = 16'h6060;
    LUT4 i12551_2_lut_rep_339_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[0]), 
         .Z(n34701)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12551_2_lut_rep_339_3_lut.init = 16'h6060;
    LUT4 i12894_2_lut_rep_340_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(op_i_23__N_1154[1]), 
         .Z(n34702)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12894_2_lut_rep_340_3_lut.init = 16'h6060;
    LUT4 i206_2_lut_rep_385_3_lut (.A(\rom8_state[0] ), .B(n34794), .C(valid), 
         .Z(clk_c_enable_1373)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i206_2_lut_rep_385_3_lut.init = 16'hf6f6;
    LUT4 mux_403_i7_3_lut_4_lut (.A(op_i_23__N_1154[6]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[6]), .Z(n7590[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i7_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13763_3_lut_4_lut (.A(op_i_23__N_1154[6]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[14]_adj_70 ), .Z(n31508)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13763_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i8_3_lut_4_lut (.A(op_i_23__N_1154[7]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[7]), .Z(n7590[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13761_3_lut_4_lut (.A(op_i_23__N_1154[7]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[15]_adj_71 ), .Z(n31506)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13761_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i7_3_lut_4_lut (.A(op_r_23__N_1106[6]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[6]), .Z(n7431[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i7_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13714_3_lut_4_lut (.A(op_r_23__N_1106[6]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[14]_adj_72 ), .Z(n31459)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13714_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i8_3_lut_4_lut (.A(op_r_23__N_1106[7]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[7]), .Z(n7431[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13712_3_lut_4_lut (.A(op_r_23__N_1106[7]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[15]_adj_73 ), .Z(n31457)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13712_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i6_3_lut_4_lut (.A(op_i_23__N_1154[5]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[5]), .Z(n7590[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i6_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13765_3_lut_4_lut (.A(op_i_23__N_1154[5]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[13]_adj_74 ), .Z(n31510)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13765_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i5_3_lut_4_lut (.A(op_r_23__N_1106[4]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[4]), .Z(n7431[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i5_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13718_3_lut_4_lut (.A(op_r_23__N_1106[4]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[12]_adj_75 ), .Z(n31463)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13718_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i6_3_lut_4_lut (.A(op_r_23__N_1106[5]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[5]), .Z(n7431[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i6_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13716_3_lut_4_lut (.A(op_r_23__N_1106[5]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[13]_adj_76 ), .Z(n31461)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13716_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i5_3_lut_4_lut (.A(op_i_23__N_1154[4]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[4]), .Z(n7590[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i5_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13767_3_lut_4_lut (.A(op_i_23__N_1154[4]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[12]_adj_77 ), .Z(n31512)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13767_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i3_3_lut_4_lut (.A(op_r_23__N_1106[2]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[2]), .Z(n7431[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13686_3_lut_4_lut (.A(op_r_23__N_1106[20]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[28] ), .Z(n31431)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13686_3_lut_4_lut.init = 16'hf808;
    LUT4 i13722_3_lut_4_lut (.A(op_r_23__N_1106[2]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[10]_adj_78 ), .Z(n31467)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13722_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i4_3_lut_4_lut (.A(op_r_23__N_1106[3]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[3]), .Z(n7431[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13720_3_lut_4_lut (.A(op_r_23__N_1106[3]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[11]_adj_79 ), .Z(n31465)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13720_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i3_3_lut_4_lut (.A(op_i_23__N_1154[2]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[2]), .Z(n7590[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13771_3_lut_4_lut (.A(op_i_23__N_1154[2]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[10]_adj_80 ), .Z(n31516)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13771_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i4_3_lut_4_lut (.A(op_i_23__N_1154[3]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[3]), .Z(n7590[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13769_3_lut_4_lut (.A(op_i_23__N_1154[3]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[11]_adj_81 ), .Z(n31514)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13769_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i1_3_lut_4_lut (.A(op_r_23__N_1106[0]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[0]), .Z(n7431[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i1_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13726_3_lut_4_lut (.A(op_r_23__N_1106[0]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[8]_adj_82 ), .Z(n31471)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13726_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_391_i2_3_lut_4_lut (.A(op_r_23__N_1106[1]), .B(n34842), .C(n3), 
         .D(shift_4_dout_r[1]), .Z(n7431[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_391_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13724_3_lut_4_lut (.A(op_r_23__N_1106[1]), .B(n34842), .C(n6514), 
         .D(\op_r_23__N_1082[9]_adj_83 ), .Z(n31469)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13724_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i1_3_lut_4_lut (.A(op_i_23__N_1154[0]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[0]), .Z(n7590[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i1_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13775_3_lut_4_lut (.A(op_i_23__N_1154[0]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[8]_adj_84 ), .Z(n31520)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13775_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i2_3_lut_4_lut (.A(op_i_23__N_1154[1]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[1]), .Z(n7590[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13773_3_lut_4_lut (.A(op_i_23__N_1154[1]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[9]_adj_85 ), .Z(n31518)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13773_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i22_3_lut_4_lut (.A(op_i_23__N_1154[21]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[21]), .Z(n7590[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i22_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13733_3_lut_4_lut (.A(op_i_23__N_1154[21]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[29] ), .Z(n31478)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13733_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_403_i21_3_lut_4_lut (.A(op_i_23__N_1154[20]), .B(n34842), .C(n3), 
         .D(shift_4_dout_i[20]), .Z(n7590[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_403_i21_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13735_3_lut_4_lut (.A(op_i_23__N_1154[20]), .B(n34842), .C(n6514), 
         .D(\op_i_23__N_1130[28] ), .Z(n31480)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13735_3_lut_4_lut.init = 16'hf808;
    
endmodule
//
// Verilog Description of module radix2_U1
//

module radix2_U1 (shift_4_dout_i, n12300, n12301, n12302, n12303, 
            n12304, n12305, n12306, n12307, n12308, n12309, n119, 
            GND_net, VCC_net, \op_r_23__N_1268[0] , \op_r_23__N_1268[1] , 
            \op_r_23__N_1268[2] , \op_r_23__N_1268[3] , \op_r_23__N_1268[4] , 
            \op_r_23__N_1268[5] , \op_r_23__N_1268[6] , \op_r_23__N_1268[7] , 
            \op_r_23__N_1268[8] , \op_r_23__N_1268[9] , \op_r_23__N_1268[10] , 
            \op_r_23__N_1268[11] , \op_r_23__N_1268[12] , \op_r_23__N_1268[13] , 
            \op_r_23__N_1268[14] , \op_r_23__N_1268[15] , \op_r_23__N_1268[16] , 
            \op_r_23__N_1268[17] , \op_r_23__N_1226[0] , \op_r_23__N_1226[1] , 
            \op_r_23__N_1226[2] , \op_r_23__N_1226[3] , \op_r_23__N_1226[4] , 
            \op_r_23__N_1226[5] , \op_r_23__N_1226[6] , \op_r_23__N_1226[7] , 
            \op_r_23__N_1226[8] , \op_r_23__N_1226[9] , \op_r_23__N_1226[10] , 
            \op_r_23__N_1226[11] , \op_r_23__N_1226[12] , \op_r_23__N_1226[13] , 
            \op_r_23__N_1226[14] , \op_r_23__N_1226[15] , \op_r_23__N_1226[16] , 
            \op_r_23__N_1226[17] , \op_r_23__N_1226[18] , \op_r_23__N_1226[19] , 
            \op_r_23__N_1226[20] , \op_r_23__N_1226[21] , \op_r_23__N_1226[22] , 
            \op_r_23__N_1226[23] , \op_r_23__N_1226[24] , \op_r_23__N_1226[25] , 
            \op_r_23__N_1226[26] , \op_r_23__N_1226[27] , \op_r_23__N_1226[28] , 
            \op_r_23__N_1226[29] , \op_r_23__N_1226[30] , \op_r_23__N_1226[31] , 
            \op_r_23__N_1268[18] , \op_r_23__N_1268[19] , \op_r_23__N_1268[20] , 
            \op_r_23__N_1268[21] , \op_r_23__N_1268[22] , \op_r_23__N_1268[23] , 
            \op_r_23__N_1268[24] , \op_r_23__N_1268[25] , \op_r_23__N_1268[26] , 
            \op_r_23__N_1268[27] , \op_r_23__N_1268[28] , \op_r_23__N_1268[29] , 
            \op_r_23__N_1268[30] , \op_r_23__N_1268[31] , n8849, n8848, 
            n8847, n8846, n8845, n8844, n8843, n8842, n8841, n8840, 
            n8839, n8838, n8837, n8836, n8835, n8834, n8833, n8832, 
            n8831, n8830, n8829, n8828, n8827, n8826, n8825, n8824, 
            n34777, \rom4_w_r[1] , \rom4_w_r[5] , \rom4_w_r[8] , n12240, 
            n12241, n12242, n12243, n12244, n12245, n12246, n12247, 
            n12248, n12249, n12250, n12251, n12252, n12253, n12254, 
            n12255, n12256, n12257, \rom4_w_i[12] , n319, n10718, 
            n10719, n10720, n10721, n10722, n10723, n10724, n10725, 
            n10726, n10727, n10728, n10729, n10730, n10731, n10732, 
            n10733, n10734, n10735, n12258, n12259, n12260, n12261, 
            n12262, n12263, n12264, op_i_23__N_1154, n34841, n30179, 
            \delay_i_23__N_1202[18] , \dout_i_23__N_5777[18] , \delay_i_23__N_1202[2] , 
            \dout_i_23__N_5777[2] , \delay_i_23__N_1202[1] , \dout_i_23__N_5777[1] , 
            \delay_i_23__N_1202[0] , \dout_i_23__N_5777[0] , \rom4_state[0] , 
            n34799, op_r_23__N_1106, n34610, n34609, n34576, n34575, 
            n34690, n34612, valid, clk_c_enable_1396, n34621, n34665, 
            n34593, n34578, \delay_r_23__N_1178[0] , \dout_r_23__N_5681[0] , 
            n34624, n34579, n34587, n34588, n34666, n34594, n34622, 
            n34577, n34623, n34611, n34689, n34633, n34580, n34634, 
            n34581, n34635, n34582, n34636, n34583, n34645, n34584, 
            n34646, n34585, n34655, n34586, n34656, n34667, n34595, 
            n34668, n34596, n34673, n34601, n34674, n34602, n34679, 
            n34603, n34604, n34680) /* synthesis syn_module_defined=1 */ ;
    input [23:0]shift_4_dout_i;
    input n12300;
    input n12301;
    input n12302;
    input n12303;
    input n12304;
    input n12305;
    input n12306;
    input n12307;
    input n12308;
    input n12309;
    input n119;
    input GND_net;
    input VCC_net;
    output \op_r_23__N_1268[0] ;
    output \op_r_23__N_1268[1] ;
    output \op_r_23__N_1268[2] ;
    output \op_r_23__N_1268[3] ;
    output \op_r_23__N_1268[4] ;
    output \op_r_23__N_1268[5] ;
    output \op_r_23__N_1268[6] ;
    output \op_r_23__N_1268[7] ;
    output \op_r_23__N_1268[8] ;
    output \op_r_23__N_1268[9] ;
    output \op_r_23__N_1268[10] ;
    output \op_r_23__N_1268[11] ;
    output \op_r_23__N_1268[12] ;
    output \op_r_23__N_1268[13] ;
    output \op_r_23__N_1268[14] ;
    output \op_r_23__N_1268[15] ;
    output \op_r_23__N_1268[16] ;
    output \op_r_23__N_1268[17] ;
    output \op_r_23__N_1226[0] ;
    output \op_r_23__N_1226[1] ;
    output \op_r_23__N_1226[2] ;
    output \op_r_23__N_1226[3] ;
    output \op_r_23__N_1226[4] ;
    output \op_r_23__N_1226[5] ;
    output \op_r_23__N_1226[6] ;
    output \op_r_23__N_1226[7] ;
    output \op_r_23__N_1226[8] ;
    output \op_r_23__N_1226[9] ;
    output \op_r_23__N_1226[10] ;
    output \op_r_23__N_1226[11] ;
    output \op_r_23__N_1226[12] ;
    output \op_r_23__N_1226[13] ;
    output \op_r_23__N_1226[14] ;
    output \op_r_23__N_1226[15] ;
    output \op_r_23__N_1226[16] ;
    output \op_r_23__N_1226[17] ;
    output \op_r_23__N_1226[18] ;
    output \op_r_23__N_1226[19] ;
    output \op_r_23__N_1226[20] ;
    output \op_r_23__N_1226[21] ;
    output \op_r_23__N_1226[22] ;
    output \op_r_23__N_1226[23] ;
    output \op_r_23__N_1226[24] ;
    output \op_r_23__N_1226[25] ;
    output \op_r_23__N_1226[26] ;
    output \op_r_23__N_1226[27] ;
    output \op_r_23__N_1226[28] ;
    output \op_r_23__N_1226[29] ;
    output \op_r_23__N_1226[30] ;
    output \op_r_23__N_1226[31] ;
    output \op_r_23__N_1268[18] ;
    output \op_r_23__N_1268[19] ;
    output \op_r_23__N_1268[20] ;
    output \op_r_23__N_1268[21] ;
    output \op_r_23__N_1268[22] ;
    output \op_r_23__N_1268[23] ;
    output \op_r_23__N_1268[24] ;
    output \op_r_23__N_1268[25] ;
    output \op_r_23__N_1268[26] ;
    output \op_r_23__N_1268[27] ;
    output \op_r_23__N_1268[28] ;
    output \op_r_23__N_1268[29] ;
    output \op_r_23__N_1268[30] ;
    output \op_r_23__N_1268[31] ;
    output n8849;
    output n8848;
    output n8847;
    output n8846;
    output n8845;
    output n8844;
    output n8843;
    output n8842;
    output n8841;
    output n8840;
    output n8839;
    output n8838;
    output n8837;
    output n8836;
    output n8835;
    output n8834;
    output n8833;
    output n8832;
    output n8831;
    output n8830;
    output n8829;
    output n8828;
    output n8827;
    output n8826;
    output n8825;
    output n8824;
    input n34777;
    input \rom4_w_r[1] ;
    input \rom4_w_r[5] ;
    input \rom4_w_r[8] ;
    input n12240;
    input n12241;
    input n12242;
    input n12243;
    input n12244;
    input n12245;
    input n12246;
    input n12247;
    input n12248;
    input n12249;
    input n12250;
    input n12251;
    input n12252;
    input n12253;
    input n12254;
    input n12255;
    input n12256;
    input n12257;
    input \rom4_w_i[12] ;
    input n319;
    input n10718;
    input n10719;
    input n10720;
    input n10721;
    input n10722;
    input n10723;
    input n10724;
    input n10725;
    input n10726;
    input n10727;
    input n10728;
    input n10729;
    input n10730;
    input n10731;
    input n10732;
    input n10733;
    input n10734;
    input n10735;
    input n12258;
    input n12259;
    input n12260;
    input n12261;
    input n12262;
    input n12263;
    input n12264;
    input [23:0]op_i_23__N_1154;
    input n34841;
    input n30179;
    input \delay_i_23__N_1202[18] ;
    output \dout_i_23__N_5777[18] ;
    input \delay_i_23__N_1202[2] ;
    output \dout_i_23__N_5777[2] ;
    input \delay_i_23__N_1202[1] ;
    output \dout_i_23__N_5777[1] ;
    input \delay_i_23__N_1202[0] ;
    output \dout_i_23__N_5777[0] ;
    input \rom4_state[0] ;
    input n34799;
    input [23:0]op_r_23__N_1106;
    output n34610;
    output n34609;
    output n34576;
    output n34575;
    output n34690;
    output n34612;
    input valid;
    output clk_c_enable_1396;
    output n34621;
    output n34665;
    output n34593;
    output n34578;
    input \delay_r_23__N_1178[0] ;
    output \dout_r_23__N_5681[0] ;
    output n34624;
    output n34579;
    output n34587;
    output n34588;
    output n34666;
    output n34594;
    output n34622;
    output n34577;
    output n34623;
    output n34611;
    output n34689;
    output n34633;
    output n34580;
    output n34634;
    output n34581;
    output n34635;
    output n34582;
    output n34636;
    output n34583;
    output n34645;
    output n34584;
    output n34646;
    output n34585;
    output n34655;
    output n34586;
    output n34656;
    output n34667;
    output n34595;
    output n34668;
    output n34596;
    output n34673;
    output n34601;
    output n34674;
    output n34602;
    output n34679;
    output n34603;
    output n34604;
    output n34680;
    
    
    wire n17052, n17053, n17054, n17055, n17056, n17057, n17058, 
        n17059, n17060, n17061, n17062, n17063, n17064, n17065, 
        n17066, n17067, n17068, n17069, n17070, n17071, n17072, 
        n17073, n17074, n17075, n17076, n17077, n17078, n17079, 
        n17080, n17081, n17082, n17083, n17084, n17085, n17086, 
        n17087, n17088, n17089, n17090, n17091, n17092, n17093, 
        n17094, n17095, n17096, n17097, n17098, n17099, n17100, 
        n17101, n17102, n17103, n17104, n17105, n17106, n17107, 
        n17108, n17109, n17110, n17111, n17112, n17113, n17114, 
        n17115, n17116, n17117, n17118, n17119, n17120, n17121, 
        n17122, n17123, n17124, n17125, n17126, n17127, n17128, 
        n17129, n17130, n17131, n17132, n17133, n17134, n17135, 
        n17136, n17137, n17138, n17139, n17140, n17141, n17142, 
        n17143, n17144, n17145, n17146, n17147, n17148, n17149, 
        n17150, n17151, n17152, n17153, n17154, n17155, n17156, 
        n17157, n17158, n17159, n17160, n17161, n17162, n17163, 
        n17164, n17165, n17166, n17167, n17168, n17169, n17170, 
        n17171, n17172, n17173, n17174, n17175, n17176, n17177, 
        n17178, n17179, n17180, n17181, n17182, n17183, n17184, 
        n17185, n17186, n17187, n17188, n17189, n17190, n17191, 
        n17192, n17193, n17194, n17195, n17196, n17197, n17344, 
        n17345, n17346, n17347, n17348, n17349, n17350, n17351, 
        n17352, n17353, n17354, n17355, n17356, n17357, n17358, 
        n17359, n17360, n17361, n17362, n17363, n17364, n17365, 
        n17366, n17367, n17368, n17369, n17370, n17371, n17372, 
        n17373, n17374, n17375, n17376, n17377, n17378, n17379, 
        n17380, n16852, n16853, n16854, n16855, n16856, n16857, 
        n16858, n16859, n16860, n16861, n16862, n16863, n16864, 
        n16865, n16866, n16867, n16868, n16869, n16870, n16871, 
        n16872, n16873, n16874, n16875, n16876, n16877, n16878, 
        n16879, n16880, n16881, n16882, n16883, n16884, n16885, 
        n16886, n16887, n16888, n16889, n16890, n16891, n16892, 
        n16893, n16894, n16895, n16896, n16897, n16898, n16899, 
        n16900, n16901, n16902, n16903, n16904, n16905, n16906, 
        n16907, n16908, n16909, n16910, n16911, n16912, n16913, 
        n16914, n16915, n16916, n16917, n16918, n16919, n16920, 
        n16921, n16922, n16923, n16924, n16925, n16926, n16927, 
        n16928, n16929, n16930, n16931, n16932, n16933, n16934, 
        n16935, n16936, n16937, n16938, n16939, n16940, n16941, 
        n16942, n16943, n16944, n16945, n16946, n16947, n16948, 
        n16949, n16950, n16951, n16952, n16953, n16954, n16955, 
        n16956, n16957, n16958, n16959, n16960, n16961, n16962, 
        n16963, n16964, n16965, n16966, n16967, n16968, n16969, 
        n16970, n16971, n16972, n16973, n16974, n16975, n16976, 
        n16977, n16978, n16979, n16980, n16981, n16982, n16983, 
        n16984, n16985, n16986, n16987, n16988, n16989, n16990, 
        n16991, n16992, n16993, n16994, n16995, n16996, n16997, 
        n16998, n16999, n17000, n17001, n17002, n17003, n17004, 
        n17005, n17006, n17007, n17008, n17009, n17010, n17011, 
        n17012, n17013, n17014, n17015, n17016, n17017, n17018, 
        n17019, n17020, n17021, n17022, n17023, n17024, n17025, 
        n17026, n17027, n17028, n17029, n17030, n17031, n17032, 
        n17033, n17034, n17198, n17199, n17200, n17201, n17202, 
        n17203, n17204, n17205, n17206, n17207, n17208, n17209, 
        n17210, n17211, n17212, n17213, n17214, n17215, n17216, 
        n17217, n17218, n17219, n17220, n17221, n17222, n17223, 
        n17224, n17225, n17226, n17227, n17228, n17229, n17230, 
        n17231, n17232, n17233, n17234, n17235, n17236, n17237, 
        n17238, n17239, n17240, n17241, n17242, n17243, n17244, 
        n17245, n17246, n17247, n17248, n17249, n17250, n17251, 
        n17252, n17253, n17254, n17255, n17256, n17257, n17258, 
        n17259, n17260, n17261, n17262, n17263, n17264, n17265, 
        n17266, n17267, n17268, n17269, n17270, n17271, n17272, 
        n17273, n17274, n17275, n17276, n17277, n17278, n17279, 
        n17280, n17281, n17282, n17283, n17284, n17285, n17286, 
        n17287, n17288, n17289, n17290, n17291, n17292, n17293, 
        n17294, n17295, n17296, n17297, n17298, n17299, n17300, 
        n17301, n17302, n17303, n17304, n17305, n17306, n17307, 
        n17308, n17309, n17310, n17311, n17312, n17313, n17314, 
        n17315, n17316, n17317, n17318, n17319, n17320, n17321, 
        n17322, n17323, n17324, n17325, n17326, n17327, n17328, 
        n17329, n17330, n17331, n17332, n17333, n17334, n17335, 
        n17336, n17337, n17338, n17339, n17340, n17341, n17342, 
        n17343, n16706, n16707, n16708, n16709, n16710, n16711, 
        n16712, n16713, n16714, n16715, n16716, n16717, n16718, 
        n16719, n16720, n16721, n16722, n16723, n16724, n16725, 
        n16726, n16727, n16728, n16729, n16730, n16731, n16732, 
        n16733, n16734, n16735, n16736, n16737, n16738, n16739, 
        n16740, n16741, n16742, n16743, n16744, n16745, n16746, 
        n16747, n16748, n16749, n16750, n16751, n16752, n16753, 
        n16754, n16755, n16756, n16757, n16758, n16759, n16760, 
        n16761, n16762, n16763, n16764, n16765, n16766, n16767, 
        n16768, n16769, n16770, n16771, n16772, n16773, n16774, 
        n16775, n16776, n16777, n16778, n16779, n16780, n16781, 
        n16782, n16783, n16784, n16785, n16786, n16787, n16788, 
        n16789, n16790, n16791, n16792, n16793, n16794, n16795, 
        n16796, n16797, n16798, n16799, n16800, n16801, n16802, 
        n16803, n16804, n16805, n16806, n16807, n16808, n16809, 
        n16810, n16811, n16812, n16813, n16814, n16815, n16816, 
        n16817, n16818, n16819, n16820, n16821, n16822, n16823, 
        n16824, n16825, n16826, n16827, n16828, n16829, n16830, 
        n16831, n16832, n16833, n16834, n16835, n16836, n16837, 
        n16838, n16839, n16840, n16841, n16842, n16843, n16844, 
        n16845, n16846, n16847, n16848, n16849, n16850, n16851, 
        n14050, n14051, n14052, n14053, n14054, n14055, n14056, 
        n14057, n14058, n14059, n14060, n14061, n14062, n14063, 
        n14064, n14065, n14066, n14067, n14068, n14069, n14070, 
        n14071, n14072, n14073, n14074, n14075, n14076, n14077, 
        n14078, n14079, n14080, n14081, n14082, n14083, n14084, 
        n14085, n14086, n14087, n14088, n14089, n14090, n14091, 
        n14092, n14093, n14094, n14095, n14096, n14097, n14098, 
        n14099, n14100, n14101, n14102, n14103, n14104, n14105, 
        n14106, n14107, n14108, n14109, n14110, n14111, n14112, 
        n14113, n14114, n14115, n14116, n14117, n14118, n14119, 
        n14120, n14121, n14122, n14123, n14124, n14125, n14126, 
        n14127, n14128, n14129, n14130, n14131, n14132, n14133, 
        n14134, n14135, n14136, n14137, n14138, n14139, n14140, 
        n14141, n14142, n14143, n14144, n14145, n14146, n14147, 
        n14148, n14149, n14150, n14151, n14152, n14153, n14154, 
        n14155, n14156, n14157, n14158, n14159, n14160, n14161, 
        n14162, n14163, n14164, n14165, n14166, n14167, n14168, 
        n14169, n14170, n14171, n14172, n14173, n14174, n14175, 
        n14176, n14177, n14178, n14179, n14180, n14181, n14182, 
        n14183, n14184, n14185, n14186, n14187, n14188, n14189, 
        n14190, n14191, n14192, n14193, n14194, n14195, n14196, 
        n14197, n14198, n14199, n14200, n14201, n14202, n14203, 
        n14204, n14205, n14206, n14207, n14208, n14209, n14210, 
        n14211, n14212, n14213, n14214, n14215, n14216, n14217, 
        n14218, n14219, n14220, n14221, n14222, n14223, n14224, 
        n14225, n14226, n14227, n14228, n14229, n14230, n14231, 
        n14232, n13904, n13905, n13906, n13907, n13908, n13909, 
        n13910, n13911, n13912, n13913, n13914, n13915, n13916, 
        n13917, n13918, n13919, n13920, n13921, n13922, n13923, 
        n13924, n13925, n13926, n13927, n13928, n13929, n13930, 
        n13931, n13932, n13933, n13934, n13935, n13936, n13937, 
        n13938, n13939, n13940, n13941, n13942, n13943, n13944, 
        n13945, n13946, n13947, n13948, n13949, n13950, n13951, 
        n13952, n13953, n13954, n13955, n13956, n13957, n13958, 
        n13959, n13960, n13961, n13962, n13963, n13964, n13965, 
        n13966, n13967, n13968, n13969, n13970, n13971, n13972, 
        n13973, n13974, n13975, n13976, n13977, n13978, n13979, 
        n13980, n13981, n13982, n13983, n13984, n13985, n13986, 
        n13987, n13988, n13989, n13990, n13991, n13992, n13993, 
        n13994, n13995, n13996, n13997, n13998, n13999, n14000, 
        n14001, n14002, n14003, n14004, n14005, n14006, n14007, 
        n14008, n14009, n14010, n14011, n14012, n14013, n14014, 
        n14015, n14016, n14017, n14018, n14019, n14020, n14021, 
        n14022, n14023, n14024, n14025, n14026, n14027, n14028, 
        n14029, n14030, n14031, n14032, n14033, n14034, n14035, 
        n14036, n14037, n14038, n14039, n14040, n14041, n14042, 
        n14043, n14044, n14045, n14046, n14047, n14048, n14049;
    
    MULT18X18D mult_8 (.A17(shift_4_dout_i[17]), .A16(shift_4_dout_i[16]), 
            .A15(shift_4_dout_i[15]), .A14(shift_4_dout_i[14]), .A13(shift_4_dout_i[13]), 
            .A12(shift_4_dout_i[12]), .A11(shift_4_dout_i[11]), .A10(shift_4_dout_i[10]), 
            .A9(shift_4_dout_i[9]), .A8(shift_4_dout_i[8]), .A7(shift_4_dout_i[7]), 
            .A6(shift_4_dout_i[6]), .A5(shift_4_dout_i[5]), .A4(shift_4_dout_i[4]), 
            .A3(shift_4_dout_i[3]), .A2(shift_4_dout_i[2]), .A1(shift_4_dout_i[1]), 
            .A0(shift_4_dout_i[0]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n12309), .B8(n12308), .B7(n12307), .B6(n12306), .B5(n12305), 
            .B4(n12304), .B3(n12303), .B2(n12302), .B1(n12301), .B0(n12300), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17069), .ROA16(n17068), 
            .ROA15(n17067), .ROA14(n17066), .ROA13(n17065), .ROA12(n17064), 
            .ROA11(n17063), .ROA10(n17062), .ROA9(n17061), .ROA8(n17060), 
            .ROA7(n17059), .ROA6(n17058), .ROA5(n17057), .ROA4(n17056), 
            .ROA3(n17055), .ROA2(n17054), .ROA1(n17053), .ROA0(n17052), 
            .ROB17(n17087), .ROB16(n17086), .ROB15(n17085), .ROB14(n17084), 
            .ROB13(n17083), .ROB12(n17082), .ROB11(n17081), .ROB10(n17080), 
            .ROB9(n17079), .ROB8(n17078), .ROB7(n17077), .ROB6(n17076), 
            .ROB5(n17075), .ROB4(n17074), .ROB3(n17073), .ROB2(n17072), 
            .ROB1(n17071), .ROB0(n17070), .P35(n17124), .P34(n17123), 
            .P33(n17122), .P32(n17121), .P31(n17120), .P30(n17119), 
            .P29(n17118), .P28(n17117), .P27(n17116), .P26(n17115), 
            .P25(n17114), .P24(n17113), .P23(n17112), .P22(n17111), 
            .P21(n17110), .P20(n17109), .P19(n17108), .P18(n17107), 
            .P17(n17106), .P16(n17105), .P15(n17104), .P14(n17103), 
            .P13(n17102), .P12(n17101), .P11(n17100), .P10(n17099), 
            .P9(n17098), .P8(n17097), .P7(n17096), .P6(n17095), .P5(n17094), 
            .P4(n17093), .P3(n17092), .P2(n17091), .P1(n17090), .P0(n17089), 
            .SIGNEDP(n17088));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam mult_8.REG_INPUTA_CLK = "NONE";
    defparam mult_8.REG_INPUTA_CE = "CE0";
    defparam mult_8.REG_INPUTA_RST = "RST0";
    defparam mult_8.REG_INPUTB_CLK = "NONE";
    defparam mult_8.REG_INPUTB_CE = "CE0";
    defparam mult_8.REG_INPUTB_RST = "RST0";
    defparam mult_8.REG_INPUTC_CLK = "NONE";
    defparam mult_8.REG_INPUTC_CE = "CE0";
    defparam mult_8.REG_INPUTC_RST = "RST0";
    defparam mult_8.REG_PIPELINE_CLK = "NONE";
    defparam mult_8.REG_PIPELINE_CE = "CE0";
    defparam mult_8.REG_PIPELINE_RST = "RST0";
    defparam mult_8.REG_OUTPUT_CLK = "NONE";
    defparam mult_8.REG_OUTPUT_CE = "CE0";
    defparam mult_8.REG_OUTPUT_RST = "RST0";
    defparam mult_8.CLK0_DIV = "ENABLED";
    defparam mult_8.CLK1_DIV = "ENABLED";
    defparam mult_8.CLK2_DIV = "ENABLED";
    defparam mult_8.CLK3_DIV = "ENABLED";
    defparam mult_8.HIGHSPEED_CLK = "NONE";
    defparam mult_8.GSR = "DISABLED";
    defparam mult_8.CAS_MATCH_REG = "FALSE";
    defparam mult_8.SOURCEB_MODE = "B_SHIFT";
    defparam mult_8.MULT_BYPASS = "DISABLED";
    defparam mult_8.RESETMODE = "SYNC";
    ALU54B lat_alu_58 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n17088), .SIGNEDIB(n17161), .SIGNEDCIN(GND_net), 
           .A35(n17087), .A34(n17086), .A33(n17085), .A32(n17084), .A31(n17083), 
           .A30(n17082), .A29(n17081), .A28(n17080), .A27(n17079), .A26(n17078), 
           .A25(n17077), .A24(n17076), .A23(n17075), .A22(n17074), .A21(n17073), 
           .A20(n17072), .A19(n17071), .A18(n17070), .A17(n17069), .A16(n17068), 
           .A15(n17067), .A14(n17066), .A13(n17065), .A12(n17064), .A11(n17063), 
           .A10(n17062), .A9(n17061), .A8(n17060), .A7(n17059), .A6(n17058), 
           .A5(n17057), .A4(n17056), .A3(n17055), .A2(n17054), .A1(n17053), 
           .A0(n17052), .B35(n17160), .B34(n17159), .B33(n17158), .B32(n17157), 
           .B31(n17156), .B30(n17155), .B29(n17154), .B28(n17153), .B27(n17152), 
           .B26(n17151), .B25(n17150), .B24(n17149), .B23(n17148), .B22(n17147), 
           .B21(n17146), .B20(n17145), .B19(n17144), .B18(n17143), .B17(n17142), 
           .B16(n17141), .B15(n17140), .B14(n17139), .B13(n17138), .B12(n17137), 
           .B11(n17136), .B10(n17135), .B9(n17134), .B8(n17133), .B7(n17132), 
           .B6(n17131), .B5(n17130), .B4(n17129), .B3(n17128), .B2(n17127), 
           .B1(n17126), .B0(n17125), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n17124), .MA34(n17123), .MA33(n17122), .MA32(n17121), 
           .MA31(n17120), .MA30(n17119), .MA29(n17118), .MA28(n17117), 
           .MA27(n17116), .MA26(n17115), .MA25(n17114), .MA24(n17113), 
           .MA23(n17112), .MA22(n17111), .MA21(n17110), .MA20(n17109), 
           .MA19(n17108), .MA18(n17107), .MA17(n17106), .MA16(n17105), 
           .MA15(n17104), .MA14(n17103), .MA13(n17102), .MA12(n17101), 
           .MA11(n17100), .MA10(n17099), .MA9(n17098), .MA8(n17097), 
           .MA7(n17096), .MA6(n17095), .MA5(n17094), .MA4(n17093), .MA3(n17092), 
           .MA2(n17091), .MA1(n17090), .MA0(n17089), .MB35(n17197), 
           .MB34(n17196), .MB33(n17195), .MB32(n17194), .MB31(n17193), 
           .MB30(n17192), .MB29(n17191), .MB28(n17190), .MB27(n17189), 
           .MB26(n17188), .MB25(n17187), .MB24(n17186), .MB23(n17185), 
           .MB22(n17184), .MB21(n17183), .MB20(n17182), .MB19(n17181), 
           .MB18(n17180), .MB17(n17179), .MB16(n17178), .MB15(n17177), 
           .MB14(n17176), .MB13(n17175), .MB12(n17174), .MB11(n17173), 
           .MB10(n17172), .MB9(n17171), .MB8(n17170), .MB7(n17169), 
           .MB6(n17168), .MB5(n17167), .MB4(n17166), .MB3(n17165), .MB2(n17164), 
           .MB1(n17163), .MB0(n17162), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n17379), 
           .R52(n17378), .R51(n17377), .R50(n17376), .R49(n17375), .R48(n17374), 
           .R47(n17373), .R46(n17372), .R45(n17371), .R44(n17370), .R43(n17369), 
           .R42(n17368), .R41(n17367), .R40(n17366), .R39(n17365), .R38(n17364), 
           .R37(n17363), .R36(n17362), .R35(n17361), .R34(n17360), .R33(n17359), 
           .R32(n17358), .R31(n17357), .R30(n17356), .R29(n17355), .R28(n17354), 
           .R27(n17353), .R26(n17352), .R25(n17351), .R24(n17350), .R23(n17349), 
           .R22(n17348), .R21(n17347), .R20(n17346), .R19(n17345), .R18(n17344), 
           .R17(\op_r_23__N_1268[17] ), .R16(\op_r_23__N_1268[16] ), .R15(\op_r_23__N_1268[15] ), 
           .R14(\op_r_23__N_1268[14] ), .R13(\op_r_23__N_1268[13] ), .R12(\op_r_23__N_1268[12] ), 
           .R11(\op_r_23__N_1268[11] ), .R10(\op_r_23__N_1268[10] ), .R9(\op_r_23__N_1268[9] ), 
           .R8(\op_r_23__N_1268[8] ), .R7(\op_r_23__N_1268[7] ), .R6(\op_r_23__N_1268[6] ), 
           .R5(\op_r_23__N_1268[5] ), .R4(\op_r_23__N_1268[4] ), .R3(\op_r_23__N_1268[3] ), 
           .R2(\op_r_23__N_1268[2] ), .R1(\op_r_23__N_1268[1] ), .R0(\op_r_23__N_1268[0] ), 
           .SIGNEDR(n17380));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_58.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_58.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_58.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_58.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_58.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_58.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_58.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_58.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_58.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_58.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_58.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_58.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_58.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_58.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_58.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_58.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_58.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_58.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_58.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_58.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_58.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_58.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_58.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_58.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_58.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_58.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_58.REG_FLAG_CLK = "NONE";
    defparam lat_alu_58.REG_FLAG_CE = "CE0";
    defparam lat_alu_58.REG_FLAG_RST = "RST0";
    defparam lat_alu_58.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_58.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_58.MASK01 = "0x00000000000000";
    defparam lat_alu_58.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_58.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_58.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_58.CLK0_DIV = "ENABLED";
    defparam lat_alu_58.CLK1_DIV = "ENABLED";
    defparam lat_alu_58.CLK2_DIV = "ENABLED";
    defparam lat_alu_58.CLK3_DIV = "ENABLED";
    defparam lat_alu_58.MCPAT = "0x00000000000000";
    defparam lat_alu_58.MASKPAT = "0x00000000000000";
    defparam lat_alu_58.RNDPAT = "0x00000000000000";
    defparam lat_alu_58.GSR = "DISABLED";
    defparam lat_alu_58.RESETMODE = "SYNC";
    defparam lat_alu_58.MULT9_MODE = "DISABLED";
    defparam lat_alu_58.LEGACY = "DISABLED";
    ALU54B lat_alu_54 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n16888), .SIGNEDIB(n16961), .SIGNEDCIN(n17034), .A35(n16887), 
           .A34(n16886), .A33(n16885), .A32(n16884), .A31(n16883), .A30(n16882), 
           .A29(n16881), .A28(n16880), .A27(n16879), .A26(n16878), .A25(n16877), 
           .A24(n16876), .A23(n16875), .A22(n16874), .A21(n16873), .A20(n16872), 
           .A19(n16871), .A18(n16870), .A17(n16869), .A16(n16868), .A15(n16867), 
           .A14(n16866), .A13(n16865), .A12(n16864), .A11(n16863), .A10(n16862), 
           .A9(n16861), .A8(n16860), .A7(n16859), .A6(n16858), .A5(n16857), 
           .A4(n16856), .A3(n16855), .A2(n16854), .A1(n16853), .A0(n16852), 
           .B35(n16960), .B34(n16959), .B33(n16958), .B32(n16957), .B31(n16956), 
           .B30(n16955), .B29(n16954), .B28(n16953), .B27(n16952), .B26(n16951), 
           .B25(n16950), .B24(n16949), .B23(n16948), .B22(n16947), .B21(n16946), 
           .B20(n16945), .B19(n16944), .B18(n16943), .B17(n16942), .B16(n16941), 
           .B15(n16940), .B14(n16939), .B13(n16938), .B12(n16937), .B11(n16936), 
           .B10(n16935), .B9(n16934), .B8(n16933), .B7(n16932), .B6(n16931), 
           .B5(n16930), .B4(n16929), .B3(n16928), .B2(n16927), .B1(n16926), 
           .B0(n16925), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n16924), .MA34(n16923), .MA33(n16922), .MA32(n16921), 
           .MA31(n16920), .MA30(n16919), .MA29(n16918), .MA28(n16917), 
           .MA27(n16916), .MA26(n16915), .MA25(n16914), .MA24(n16913), 
           .MA23(n16912), .MA22(n16911), .MA21(n16910), .MA20(n16909), 
           .MA19(n16908), .MA18(n16907), .MA17(n16906), .MA16(n16905), 
           .MA15(n16904), .MA14(n16903), .MA13(n16902), .MA12(n16901), 
           .MA11(n16900), .MA10(n16899), .MA9(n16898), .MA8(n16897), 
           .MA7(n16896), .MA6(n16895), .MA5(n16894), .MA4(n16893), .MA3(n16892), 
           .MA2(n16891), .MA1(n16890), .MA0(n16889), .MB35(n16997), 
           .MB34(n16996), .MB33(n16995), .MB32(n16994), .MB31(n16993), 
           .MB30(n16992), .MB29(n16991), .MB28(n16990), .MB27(n16989), 
           .MB26(n16988), .MB25(n16987), .MB24(n16986), .MB23(n16985), 
           .MB22(n16984), .MB21(n16983), .MB20(n16982), .MB19(n16981), 
           .MB18(n16980), .MB17(n16979), .MB16(n16978), .MB15(n16977), 
           .MB14(n16976), .MB13(n16975), .MB12(n16974), .MB11(n16973), 
           .MB10(n16972), .MB9(n16971), .MB8(n16970), .MB7(n16969), 
           .MB6(n16968), .MB5(n16967), .MB4(n16966), .MB3(n16965), .MB2(n16964), 
           .MB1(n16963), .MB0(n16962), .CIN53(n17033), .CIN52(n17032), 
           .CIN51(n17031), .CIN50(n17030), .CIN49(n17029), .CIN48(n17028), 
           .CIN47(n17027), .CIN46(n17026), .CIN45(n17025), .CIN44(n17024), 
           .CIN43(n17023), .CIN42(n17022), .CIN41(n17021), .CIN40(n17020), 
           .CIN39(n17019), .CIN38(n17018), .CIN37(n17017), .CIN36(n17016), 
           .CIN35(n17015), .CIN34(n17014), .CIN33(n17013), .CIN32(n17012), 
           .CIN31(n17011), .CIN30(n17010), .CIN29(n17009), .CIN28(n17008), 
           .CIN27(n17007), .CIN26(n17006), .CIN25(n17005), .CIN24(n17004), 
           .CIN23(n17003), .CIN22(n17002), .CIN21(n17001), .CIN20(n17000), 
           .CIN19(n16999), .CIN18(n16998), .CIN17(\op_r_23__N_1226[17] ), 
           .CIN16(\op_r_23__N_1226[16] ), .CIN15(\op_r_23__N_1226[15] ), 
           .CIN14(\op_r_23__N_1226[14] ), .CIN13(\op_r_23__N_1226[13] ), 
           .CIN12(\op_r_23__N_1226[12] ), .CIN11(\op_r_23__N_1226[11] ), 
           .CIN10(\op_r_23__N_1226[10] ), .CIN9(\op_r_23__N_1226[9] ), .CIN8(\op_r_23__N_1226[8] ), 
           .CIN7(\op_r_23__N_1226[7] ), .CIN6(\op_r_23__N_1226[6] ), .CIN5(\op_r_23__N_1226[5] ), 
           .CIN4(\op_r_23__N_1226[4] ), .CIN3(\op_r_23__N_1226[3] ), .CIN2(\op_r_23__N_1226[2] ), 
           .CIN1(\op_r_23__N_1226[1] ), .CIN0(\op_r_23__N_1226[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1226[31] ), 
           .R12(\op_r_23__N_1226[30] ), .R11(\op_r_23__N_1226[29] ), .R10(\op_r_23__N_1226[28] ), 
           .R9(\op_r_23__N_1226[27] ), .R8(\op_r_23__N_1226[26] ), .R7(\op_r_23__N_1226[25] ), 
           .R6(\op_r_23__N_1226[24] ), .R5(\op_r_23__N_1226[23] ), .R4(\op_r_23__N_1226[22] ), 
           .R3(\op_r_23__N_1226[21] ), .R2(\op_r_23__N_1226[20] ), .R1(\op_r_23__N_1226[19] ), 
           .R0(\op_r_23__N_1226[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_54.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_54.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_54.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_54.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_54.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_54.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_54.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_54.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_54.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_54.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_54.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_54.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_54.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_54.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_54.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_54.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_54.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_54.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_54.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_54.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_54.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_54.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_54.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_54.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_54.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_54.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_54.REG_FLAG_CLK = "NONE";
    defparam lat_alu_54.REG_FLAG_CE = "CE0";
    defparam lat_alu_54.REG_FLAG_RST = "RST0";
    defparam lat_alu_54.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_54.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_54.MASK01 = "0x00000000000000";
    defparam lat_alu_54.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_54.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_54.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_54.CLK0_DIV = "ENABLED";
    defparam lat_alu_54.CLK1_DIV = "ENABLED";
    defparam lat_alu_54.CLK2_DIV = "ENABLED";
    defparam lat_alu_54.CLK3_DIV = "ENABLED";
    defparam lat_alu_54.MCPAT = "0x00000000000000";
    defparam lat_alu_54.MASKPAT = "0x00000000000000";
    defparam lat_alu_54.RNDPAT = "0x00000000000000";
    defparam lat_alu_54.GSR = "DISABLED";
    defparam lat_alu_54.RESETMODE = "SYNC";
    defparam lat_alu_54.MULT9_MODE = "DISABLED";
    defparam lat_alu_54.LEGACY = "DISABLED";
    ALU54B lat_alu_59 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n17234), .SIGNEDIB(n17307), .SIGNEDCIN(n17380), .A35(n17233), 
           .A34(n17232), .A33(n17231), .A32(n17230), .A31(n17229), .A30(n17228), 
           .A29(n17227), .A28(n17226), .A27(n17225), .A26(n17224), .A25(n17223), 
           .A24(n17222), .A23(n17221), .A22(n17220), .A21(n17219), .A20(n17218), 
           .A19(n17217), .A18(n17216), .A17(n17215), .A16(n17214), .A15(n17213), 
           .A14(n17212), .A13(n17211), .A12(n17210), .A11(n17209), .A10(n17208), 
           .A9(n17207), .A8(n17206), .A7(n17205), .A6(n17204), .A5(n17203), 
           .A4(n17202), .A3(n17201), .A2(n17200), .A1(n17199), .A0(n17198), 
           .B35(n17306), .B34(n17305), .B33(n17304), .B32(n17303), .B31(n17302), 
           .B30(n17301), .B29(n17300), .B28(n17299), .B27(n17298), .B26(n17297), 
           .B25(n17296), .B24(n17295), .B23(n17294), .B22(n17293), .B21(n17292), 
           .B20(n17291), .B19(n17290), .B18(n17289), .B17(n17288), .B16(n17287), 
           .B15(n17286), .B14(n17285), .B13(n17284), .B12(n17283), .B11(n17282), 
           .B10(n17281), .B9(n17280), .B8(n17279), .B7(n17278), .B6(n17277), 
           .B5(n17276), .B4(n17275), .B3(n17274), .B2(n17273), .B1(n17272), 
           .B0(n17271), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n17270), .MA34(n17269), .MA33(n17268), .MA32(n17267), 
           .MA31(n17266), .MA30(n17265), .MA29(n17264), .MA28(n17263), 
           .MA27(n17262), .MA26(n17261), .MA25(n17260), .MA24(n17259), 
           .MA23(n17258), .MA22(n17257), .MA21(n17256), .MA20(n17255), 
           .MA19(n17254), .MA18(n17253), .MA17(n17252), .MA16(n17251), 
           .MA15(n17250), .MA14(n17249), .MA13(n17248), .MA12(n17247), 
           .MA11(n17246), .MA10(n17245), .MA9(n17244), .MA8(n17243), 
           .MA7(n17242), .MA6(n17241), .MA5(n17240), .MA4(n17239), .MA3(n17238), 
           .MA2(n17237), .MA1(n17236), .MA0(n17235), .MB35(n17343), 
           .MB34(n17342), .MB33(n17341), .MB32(n17340), .MB31(n17339), 
           .MB30(n17338), .MB29(n17337), .MB28(n17336), .MB27(n17335), 
           .MB26(n17334), .MB25(n17333), .MB24(n17332), .MB23(n17331), 
           .MB22(n17330), .MB21(n17329), .MB20(n17328), .MB19(n17327), 
           .MB18(n17326), .MB17(n17325), .MB16(n17324), .MB15(n17323), 
           .MB14(n17322), .MB13(n17321), .MB12(n17320), .MB11(n17319), 
           .MB10(n17318), .MB9(n17317), .MB8(n17316), .MB7(n17315), 
           .MB6(n17314), .MB5(n17313), .MB4(n17312), .MB3(n17311), .MB2(n17310), 
           .MB1(n17309), .MB0(n17308), .CIN53(n17379), .CIN52(n17378), 
           .CIN51(n17377), .CIN50(n17376), .CIN49(n17375), .CIN48(n17374), 
           .CIN47(n17373), .CIN46(n17372), .CIN45(n17371), .CIN44(n17370), 
           .CIN43(n17369), .CIN42(n17368), .CIN41(n17367), .CIN40(n17366), 
           .CIN39(n17365), .CIN38(n17364), .CIN37(n17363), .CIN36(n17362), 
           .CIN35(n17361), .CIN34(n17360), .CIN33(n17359), .CIN32(n17358), 
           .CIN31(n17357), .CIN30(n17356), .CIN29(n17355), .CIN28(n17354), 
           .CIN27(n17353), .CIN26(n17352), .CIN25(n17351), .CIN24(n17350), 
           .CIN23(n17349), .CIN22(n17348), .CIN21(n17347), .CIN20(n17346), 
           .CIN19(n17345), .CIN18(n17344), .CIN17(\op_r_23__N_1268[17] ), 
           .CIN16(\op_r_23__N_1268[16] ), .CIN15(\op_r_23__N_1268[15] ), 
           .CIN14(\op_r_23__N_1268[14] ), .CIN13(\op_r_23__N_1268[13] ), 
           .CIN12(\op_r_23__N_1268[12] ), .CIN11(\op_r_23__N_1268[11] ), 
           .CIN10(\op_r_23__N_1268[10] ), .CIN9(\op_r_23__N_1268[9] ), .CIN8(\op_r_23__N_1268[8] ), 
           .CIN7(\op_r_23__N_1268[7] ), .CIN6(\op_r_23__N_1268[6] ), .CIN5(\op_r_23__N_1268[5] ), 
           .CIN4(\op_r_23__N_1268[4] ), .CIN3(\op_r_23__N_1268[3] ), .CIN2(\op_r_23__N_1268[2] ), 
           .CIN1(\op_r_23__N_1268[1] ), .CIN0(\op_r_23__N_1268[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1268[31] ), 
           .R12(\op_r_23__N_1268[30] ), .R11(\op_r_23__N_1268[29] ), .R10(\op_r_23__N_1268[28] ), 
           .R9(\op_r_23__N_1268[27] ), .R8(\op_r_23__N_1268[26] ), .R7(\op_r_23__N_1268[25] ), 
           .R6(\op_r_23__N_1268[24] ), .R5(\op_r_23__N_1268[23] ), .R4(\op_r_23__N_1268[22] ), 
           .R3(\op_r_23__N_1268[21] ), .R2(\op_r_23__N_1268[20] ), .R1(\op_r_23__N_1268[19] ), 
           .R0(\op_r_23__N_1268[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_59.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_59.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_59.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_59.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_59.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_59.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_59.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_59.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_59.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_59.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_59.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_59.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_59.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_59.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_59.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_59.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_59.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_59.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_59.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_59.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_59.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_59.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_59.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_59.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_59.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_59.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_59.REG_FLAG_CLK = "NONE";
    defparam lat_alu_59.REG_FLAG_CE = "CE0";
    defparam lat_alu_59.REG_FLAG_RST = "RST0";
    defparam lat_alu_59.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_59.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_59.MASK01 = "0x00000000000000";
    defparam lat_alu_59.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_59.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_59.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_59.CLK0_DIV = "ENABLED";
    defparam lat_alu_59.CLK1_DIV = "ENABLED";
    defparam lat_alu_59.CLK2_DIV = "ENABLED";
    defparam lat_alu_59.CLK3_DIV = "ENABLED";
    defparam lat_alu_59.MCPAT = "0x00000000000000";
    defparam lat_alu_59.MASKPAT = "0x00000000000000";
    defparam lat_alu_59.RNDPAT = "0x00000000000000";
    defparam lat_alu_59.GSR = "DISABLED";
    defparam lat_alu_59.RESETMODE = "SYNC";
    defparam lat_alu_59.MULT9_MODE = "DISABLED";
    defparam lat_alu_59.LEGACY = "DISABLED";
    ALU54B lat_alu_53 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n16742), .SIGNEDIB(n16815), .SIGNEDCIN(GND_net), 
           .A35(n16741), .A34(n16740), .A33(n16739), .A32(n16738), .A31(n16737), 
           .A30(n16736), .A29(n16735), .A28(n16734), .A27(n16733), .A26(n16732), 
           .A25(n16731), .A24(n16730), .A23(n16729), .A22(n16728), .A21(n16727), 
           .A20(n16726), .A19(n16725), .A18(n16724), .A17(n16723), .A16(n16722), 
           .A15(n16721), .A14(n16720), .A13(n16719), .A12(n16718), .A11(n16717), 
           .A10(n16716), .A9(n16715), .A8(n16714), .A7(n16713), .A6(n16712), 
           .A5(n16711), .A4(n16710), .A3(n16709), .A2(n16708), .A1(n16707), 
           .A0(n16706), .B35(n16814), .B34(n16813), .B33(n16812), .B32(n16811), 
           .B31(n16810), .B30(n16809), .B29(n16808), .B28(n16807), .B27(n16806), 
           .B26(n16805), .B25(n16804), .B24(n16803), .B23(n16802), .B22(n16801), 
           .B21(n16800), .B20(n16799), .B19(n16798), .B18(n16797), .B17(n16796), 
           .B16(n16795), .B15(n16794), .B14(n16793), .B13(n16792), .B12(n16791), 
           .B11(n16790), .B10(n16789), .B9(n16788), .B8(n16787), .B7(n16786), 
           .B6(n16785), .B5(n16784), .B4(n16783), .B3(n16782), .B2(n16781), 
           .B1(n16780), .B0(n16779), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n16778), .MA34(n16777), .MA33(n16776), .MA32(n16775), 
           .MA31(n16774), .MA30(n16773), .MA29(n16772), .MA28(n16771), 
           .MA27(n16770), .MA26(n16769), .MA25(n16768), .MA24(n16767), 
           .MA23(n16766), .MA22(n16765), .MA21(n16764), .MA20(n16763), 
           .MA19(n16762), .MA18(n16761), .MA17(n16760), .MA16(n16759), 
           .MA15(n16758), .MA14(n16757), .MA13(n16756), .MA12(n16755), 
           .MA11(n16754), .MA10(n16753), .MA9(n16752), .MA8(n16751), 
           .MA7(n16750), .MA6(n16749), .MA5(n16748), .MA4(n16747), .MA3(n16746), 
           .MA2(n16745), .MA1(n16744), .MA0(n16743), .MB35(n16851), 
           .MB34(n16850), .MB33(n16849), .MB32(n16848), .MB31(n16847), 
           .MB30(n16846), .MB29(n16845), .MB28(n16844), .MB27(n16843), 
           .MB26(n16842), .MB25(n16841), .MB24(n16840), .MB23(n16839), 
           .MB22(n16838), .MB21(n16837), .MB20(n16836), .MB19(n16835), 
           .MB18(n16834), .MB17(n16833), .MB16(n16832), .MB15(n16831), 
           .MB14(n16830), .MB13(n16829), .MB12(n16828), .MB11(n16827), 
           .MB10(n16826), .MB9(n16825), .MB8(n16824), .MB7(n16823), 
           .MB6(n16822), .MB5(n16821), .MB4(n16820), .MB3(n16819), .MB2(n16818), 
           .MB1(n16817), .MB0(n16816), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n17033), 
           .R52(n17032), .R51(n17031), .R50(n17030), .R49(n17029), .R48(n17028), 
           .R47(n17027), .R46(n17026), .R45(n17025), .R44(n17024), .R43(n17023), 
           .R42(n17022), .R41(n17021), .R40(n17020), .R39(n17019), .R38(n17018), 
           .R37(n17017), .R36(n17016), .R35(n17015), .R34(n17014), .R33(n17013), 
           .R32(n17012), .R31(n17011), .R30(n17010), .R29(n17009), .R28(n17008), 
           .R27(n17007), .R26(n17006), .R25(n17005), .R24(n17004), .R23(n17003), 
           .R22(n17002), .R21(n17001), .R20(n17000), .R19(n16999), .R18(n16998), 
           .R17(\op_r_23__N_1226[17] ), .R16(\op_r_23__N_1226[16] ), .R15(\op_r_23__N_1226[15] ), 
           .R14(\op_r_23__N_1226[14] ), .R13(\op_r_23__N_1226[13] ), .R12(\op_r_23__N_1226[12] ), 
           .R11(\op_r_23__N_1226[11] ), .R10(\op_r_23__N_1226[10] ), .R9(\op_r_23__N_1226[9] ), 
           .R8(\op_r_23__N_1226[8] ), .R7(\op_r_23__N_1226[7] ), .R6(\op_r_23__N_1226[6] ), 
           .R5(\op_r_23__N_1226[5] ), .R4(\op_r_23__N_1226[4] ), .R3(\op_r_23__N_1226[3] ), 
           .R2(\op_r_23__N_1226[2] ), .R1(\op_r_23__N_1226[1] ), .R0(\op_r_23__N_1226[0] ), 
           .SIGNEDR(n17034));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_53.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_53.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_53.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_53.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_53.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_53.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_53.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_53.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_53.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_53.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_53.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_53.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_53.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_53.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_53.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_53.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_53.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_53.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_53.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_53.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_53.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_53.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_53.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_53.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_53.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_53.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_53.REG_FLAG_CLK = "NONE";
    defparam lat_alu_53.REG_FLAG_CE = "CE0";
    defparam lat_alu_53.REG_FLAG_RST = "RST0";
    defparam lat_alu_53.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_53.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_53.MASK01 = "0x00000000000000";
    defparam lat_alu_53.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_53.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_53.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_53.CLK0_DIV = "ENABLED";
    defparam lat_alu_53.CLK1_DIV = "ENABLED";
    defparam lat_alu_53.CLK2_DIV = "ENABLED";
    defparam lat_alu_53.CLK3_DIV = "ENABLED";
    defparam lat_alu_53.MCPAT = "0x00000000000000";
    defparam lat_alu_53.MASKPAT = "0x00000000000000";
    defparam lat_alu_53.RNDPAT = "0x00000000000000";
    defparam lat_alu_53.GSR = "DISABLED";
    defparam lat_alu_53.RESETMODE = "SYNC";
    defparam lat_alu_53.MULT9_MODE = "DISABLED";
    defparam lat_alu_53.LEGACY = "DISABLED";
    ALU54B lat_alu_14 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n14086), .SIGNEDIB(n14159), .SIGNEDCIN(n14232), .A35(n14085), 
           .A34(n14084), .A33(n14083), .A32(n14082), .A31(n14081), .A30(n14080), 
           .A29(n14079), .A28(n14078), .A27(n14077), .A26(n14076), .A25(n14075), 
           .A24(n14074), .A23(n14073), .A22(n14072), .A21(n14071), .A20(n14070), 
           .A19(n14069), .A18(n14068), .A17(n14067), .A16(n14066), .A15(n14065), 
           .A14(n14064), .A13(n14063), .A12(n14062), .A11(n14061), .A10(n14060), 
           .A9(n14059), .A8(n14058), .A7(n14057), .A6(n14056), .A5(n14055), 
           .A4(n14054), .A3(n14053), .A2(n14052), .A1(n14051), .A0(n14050), 
           .B35(n14158), .B34(n14157), .B33(n14156), .B32(n14155), .B31(n14154), 
           .B30(n14153), .B29(n14152), .B28(n14151), .B27(n14150), .B26(n14149), 
           .B25(n14148), .B24(n14147), .B23(n14146), .B22(n14145), .B21(n14144), 
           .B20(n14143), .B19(n14142), .B18(n14141), .B17(n14140), .B16(n14139), 
           .B15(n14138), .B14(n14137), .B13(n14136), .B12(n14135), .B11(n14134), 
           .B10(n14133), .B9(n14132), .B8(n14131), .B7(n14130), .B6(n14129), 
           .B5(n14128), .B4(n14127), .B3(n14126), .B2(n14125), .B1(n14124), 
           .B0(n14123), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n14122), .MA34(n14121), .MA33(n14120), .MA32(n14119), 
           .MA31(n14118), .MA30(n14117), .MA29(n14116), .MA28(n14115), 
           .MA27(n14114), .MA26(n14113), .MA25(n14112), .MA24(n14111), 
           .MA23(n14110), .MA22(n14109), .MA21(n14108), .MA20(n14107), 
           .MA19(n14106), .MA18(n14105), .MA17(n14104), .MA16(n14103), 
           .MA15(n14102), .MA14(n14101), .MA13(n14100), .MA12(n14099), 
           .MA11(n14098), .MA10(n14097), .MA9(n14096), .MA8(n14095), 
           .MA7(n14094), .MA6(n14093), .MA5(n14092), .MA4(n14091), .MA3(n14090), 
           .MA2(n14089), .MA1(n14088), .MA0(n14087), .MB35(n14195), 
           .MB34(n14194), .MB33(n14193), .MB32(n14192), .MB31(n14191), 
           .MB30(n14190), .MB29(n14189), .MB28(n14188), .MB27(n14187), 
           .MB26(n14186), .MB25(n14185), .MB24(n14184), .MB23(n14183), 
           .MB22(n14182), .MB21(n14181), .MB20(n14180), .MB19(n14179), 
           .MB18(n14178), .MB17(n14177), .MB16(n14176), .MB15(n14175), 
           .MB14(n14174), .MB13(n14173), .MB12(n14172), .MB11(n14171), 
           .MB10(n14170), .MB9(n14169), .MB8(n14168), .MB7(n14167), 
           .MB6(n14166), .MB5(n14165), .MB4(n14164), .MB3(n14163), .MB2(n14162), 
           .MB1(n14161), .MB0(n14160), .CIN53(n14231), .CIN52(n14230), 
           .CIN51(n14229), .CIN50(n14228), .CIN49(n14227), .CIN48(n14226), 
           .CIN47(n14225), .CIN46(n14224), .CIN45(n14223), .CIN44(n14222), 
           .CIN43(n14221), .CIN42(n14220), .CIN41(n14219), .CIN40(n14218), 
           .CIN39(n14217), .CIN38(n14216), .CIN37(n14215), .CIN36(n14214), 
           .CIN35(n14213), .CIN34(n14212), .CIN33(n14211), .CIN32(n14210), 
           .CIN31(n14209), .CIN30(n14208), .CIN29(n14207), .CIN28(n14206), 
           .CIN27(n14205), .CIN26(n14204), .CIN25(n14203), .CIN24(n14202), 
           .CIN23(n14201), .CIN22(n14200), .CIN21(n14199), .CIN20(n14198), 
           .CIN19(n14197), .CIN18(n14196), .CIN17(n8832), .CIN16(n8833), 
           .CIN15(n8834), .CIN14(n8835), .CIN13(n8836), .CIN12(n8837), 
           .CIN11(n8838), .CIN10(n8839), .CIN9(n8840), .CIN8(n8841), 
           .CIN7(n8842), .CIN6(n8843), .CIN5(n8844), .CIN4(n8845), .CIN3(n8846), 
           .CIN2(n8847), .CIN1(n8848), .CIN0(n8849), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R7(n8824), .R6(n8825), .R5(n8826), 
           .R4(n8827), .R3(n8828), .R2(n8829), .R1(n8830), .R0(n8831));
    defparam lat_alu_14.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_14.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_14.REG_FLAG_CLK = "NONE";
    defparam lat_alu_14.REG_FLAG_CE = "CE0";
    defparam lat_alu_14.REG_FLAG_RST = "RST0";
    defparam lat_alu_14.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASK01 = "0x00000000000000";
    defparam lat_alu_14.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_14.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_14.CLK0_DIV = "ENABLED";
    defparam lat_alu_14.CLK1_DIV = "ENABLED";
    defparam lat_alu_14.CLK2_DIV = "ENABLED";
    defparam lat_alu_14.CLK3_DIV = "ENABLED";
    defparam lat_alu_14.MCPAT = "0x00000000000000";
    defparam lat_alu_14.MASKPAT = "0x00000000000000";
    defparam lat_alu_14.RNDPAT = "0x00000000000000";
    defparam lat_alu_14.GSR = "DISABLED";
    defparam lat_alu_14.RESETMODE = "SYNC";
    defparam lat_alu_14.MULT9_MODE = "DISABLED";
    defparam lat_alu_14.LEGACY = "DISABLED";
    ALU54B lat_alu_13 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n13940), .SIGNEDIB(n14013), .SIGNEDCIN(GND_net), 
           .A35(n13939), .A34(n13938), .A33(n13937), .A32(n13936), .A31(n13935), 
           .A30(n13934), .A29(n13933), .A28(n13932), .A27(n13931), .A26(n13930), 
           .A25(n13929), .A24(n13928), .A23(n13927), .A22(n13926), .A21(n13925), 
           .A20(n13924), .A19(n13923), .A18(n13922), .A17(n13921), .A16(n13920), 
           .A15(n13919), .A14(n13918), .A13(n13917), .A12(n13916), .A11(n13915), 
           .A10(n13914), .A9(n13913), .A8(n13912), .A7(n13911), .A6(n13910), 
           .A5(n13909), .A4(n13908), .A3(n13907), .A2(n13906), .A1(n13905), 
           .A0(n13904), .B35(n14012), .B34(n14011), .B33(n14010), .B32(n14009), 
           .B31(n14008), .B30(n14007), .B29(n14006), .B28(n14005), .B27(n14004), 
           .B26(n14003), .B25(n14002), .B24(n14001), .B23(n14000), .B22(n13999), 
           .B21(n13998), .B20(n13997), .B19(n13996), .B18(n13995), .B17(n13994), 
           .B16(n13993), .B15(n13992), .B14(n13991), .B13(n13990), .B12(n13989), 
           .B11(n13988), .B10(n13987), .B9(n13986), .B8(n13985), .B7(n13984), 
           .B6(n13983), .B5(n13982), .B4(n13981), .B3(n13980), .B2(n13979), 
           .B1(n13978), .B0(n13977), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n13976), .MA34(n13975), .MA33(n13974), .MA32(n13973), 
           .MA31(n13972), .MA30(n13971), .MA29(n13970), .MA28(n13969), 
           .MA27(n13968), .MA26(n13967), .MA25(n13966), .MA24(n13965), 
           .MA23(n13964), .MA22(n13963), .MA21(n13962), .MA20(n13961), 
           .MA19(n13960), .MA18(n13959), .MA17(n13958), .MA16(n13957), 
           .MA15(n13956), .MA14(n13955), .MA13(n13954), .MA12(n13953), 
           .MA11(n13952), .MA10(n13951), .MA9(n13950), .MA8(n13949), 
           .MA7(n13948), .MA6(n13947), .MA5(n13946), .MA4(n13945), .MA3(n13944), 
           .MA2(n13943), .MA1(n13942), .MA0(n13941), .MB35(n14049), 
           .MB34(n14048), .MB33(n14047), .MB32(n14046), .MB31(n14045), 
           .MB30(n14044), .MB29(n14043), .MB28(n14042), .MB27(n14041), 
           .MB26(n14040), .MB25(n14039), .MB24(n14038), .MB23(n14037), 
           .MB22(n14036), .MB21(n14035), .MB20(n14034), .MB19(n14033), 
           .MB18(n14032), .MB17(n14031), .MB16(n14030), .MB15(n14029), 
           .MB14(n14028), .MB13(n14027), .MB12(n14026), .MB11(n14025), 
           .MB10(n14024), .MB9(n14023), .MB8(n14022), .MB7(n14021), 
           .MB6(n14020), .MB5(n14019), .MB4(n14018), .MB3(n14017), .MB2(n14016), 
           .MB1(n14015), .MB0(n14014), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n14231), 
           .R52(n14230), .R51(n14229), .R50(n14228), .R49(n14227), .R48(n14226), 
           .R47(n14225), .R46(n14224), .R45(n14223), .R44(n14222), .R43(n14221), 
           .R42(n14220), .R41(n14219), .R40(n14218), .R39(n14217), .R38(n14216), 
           .R37(n14215), .R36(n14214), .R35(n14213), .R34(n14212), .R33(n14211), 
           .R32(n14210), .R31(n14209), .R30(n14208), .R29(n14207), .R28(n14206), 
           .R27(n14205), .R26(n14204), .R25(n14203), .R24(n14202), .R23(n14201), 
           .R22(n14200), .R21(n14199), .R20(n14198), .R19(n14197), .R18(n14196), 
           .R17(n8832), .R16(n8833), .R15(n8834), .R14(n8835), .R13(n8836), 
           .R12(n8837), .R11(n8838), .R10(n8839), .R9(n8840), .R8(n8841), 
           .R7(n8842), .R6(n8843), .R5(n8844), .R4(n8845), .R3(n8846), 
           .R2(n8847), .R1(n8848), .R0(n8849), .SIGNEDR(n14232));
    defparam lat_alu_13.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_13.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_13.REG_FLAG_CLK = "NONE";
    defparam lat_alu_13.REG_FLAG_CE = "CE0";
    defparam lat_alu_13.REG_FLAG_RST = "RST0";
    defparam lat_alu_13.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASK01 = "0x00000000000000";
    defparam lat_alu_13.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_13.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_13.CLK0_DIV = "ENABLED";
    defparam lat_alu_13.CLK1_DIV = "ENABLED";
    defparam lat_alu_13.CLK2_DIV = "ENABLED";
    defparam lat_alu_13.CLK3_DIV = "ENABLED";
    defparam lat_alu_13.MCPAT = "0x00000000000000";
    defparam lat_alu_13.MASKPAT = "0x00000000000000";
    defparam lat_alu_13.RNDPAT = "0x00000000000000";
    defparam lat_alu_13.GSR = "DISABLED";
    defparam lat_alu_13.RESETMODE = "SYNC";
    defparam lat_alu_13.MULT9_MODE = "DISABLED";
    defparam lat_alu_13.LEGACY = "DISABLED";
    MULT18X18D mult_10_mult_2 (.A17(\rom4_w_r[1] ), .A16(\rom4_w_r[1] ), 
            .A15(\rom4_w_r[1] ), .A14(\rom4_w_r[1] ), .A13(\rom4_w_r[1] ), 
            .A12(\rom4_w_r[1] ), .A11(\rom4_w_r[1] ), .A10(\rom4_w_r[1] ), 
            .A9(\rom4_w_r[1] ), .A8(\rom4_w_r[8] ), .A7(\rom4_w_r[5] ), 
            .A6(\rom4_w_r[1] ), .A5(\rom4_w_r[5] ), .A4(\rom4_w_r[5] ), 
            .A3(\rom4_w_r[1] ), .A2(\rom4_w_r[5] ), .A1(\rom4_w_r[1] ), 
            .A0(n34777), .B17(n12257), .B16(n12256), .B15(n12255), .B14(n12254), 
            .B13(n12253), .B12(n12252), .B11(n12251), .B10(n12250), 
            .B9(n12249), .B8(n12248), .B7(n12247), .B6(n12246), .B5(n12245), 
            .B4(n12244), .B3(n12243), .B2(n12242), .B1(n12241), .B0(n12240), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n16723), .ROA16(n16722), 
            .ROA15(n16721), .ROA14(n16720), .ROA13(n16719), .ROA12(n16718), 
            .ROA11(n16717), .ROA10(n16716), .ROA9(n16715), .ROA8(n16714), 
            .ROA7(n16713), .ROA6(n16712), .ROA5(n16711), .ROA4(n16710), 
            .ROA3(n16709), .ROA2(n16708), .ROA1(n16707), .ROA0(n16706), 
            .ROB17(n16741), .ROB16(n16740), .ROB15(n16739), .ROB14(n16738), 
            .ROB13(n16737), .ROB12(n16736), .ROB11(n16735), .ROB10(n16734), 
            .ROB9(n16733), .ROB8(n16732), .ROB7(n16731), .ROB6(n16730), 
            .ROB5(n16729), .ROB4(n16728), .ROB3(n16727), .ROB2(n16726), 
            .ROB1(n16725), .ROB0(n16724), .P35(n16778), .P34(n16777), 
            .P33(n16776), .P32(n16775), .P31(n16774), .P30(n16773), 
            .P29(n16772), .P28(n16771), .P27(n16770), .P26(n16769), 
            .P25(n16768), .P24(n16767), .P23(n16766), .P22(n16765), 
            .P21(n16764), .P20(n16763), .P19(n16762), .P18(n16761), 
            .P17(n16760), .P16(n16759), .P15(n16758), .P14(n16757), 
            .P13(n16756), .P12(n16755), .P11(n16754), .P10(n16753), 
            .P9(n16752), .P8(n16751), .P7(n16750), .P6(n16749), .P5(n16748), 
            .P4(n16747), .P3(n16746), .P2(n16745), .P1(n16744), .P0(n16743), 
            .SIGNEDP(n16742));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam mult_10_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_10_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_10_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_10_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_10_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_10_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_10_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_10_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_10_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_10_mult_2.GSR = "DISABLED";
    defparam mult_10_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_10_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_10_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_10_mult_2.RESETMODE = "SYNC";
    MULT18X18D lat_mult_12 (.A17(\rom4_w_i[12] ), .A16(\rom4_w_i[12] ), 
            .A15(\rom4_w_i[12] ), .A14(\rom4_w_i[12] ), .A13(\rom4_w_i[12] ), 
            .A12(\rom4_w_i[12] ), .A11(\rom4_w_i[12] ), .A10(\rom4_w_i[12] ), 
            .A9(\rom4_w_i[12] ), .A8(\rom4_w_i[12] ), .A7(\rom4_w_i[12] ), 
            .A6(\rom4_w_i[12] ), .A5(\rom4_w_i[12] ), .A4(\rom4_w_i[12] ), 
            .A3(\rom4_w_i[12] ), .A2(\rom4_w_i[12] ), .A1(\rom4_w_i[12] ), 
            .A0(\rom4_w_i[12] ), .B17(n319), .B16(n319), .B15(n319), 
            .B14(n319), .B13(n319), .B12(n319), .B11(n319), .B10(n319), 
            .B9(n319), .B8(n319), .B7(n319), .B6(n319), .B5(n319), 
            .B4(n319), .B3(n319), .B2(n319), .B1(n319), .B0(n319), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14140), .ROA16(n14139), 
            .ROA15(n14138), .ROA14(n14137), .ROA13(n14136), .ROA12(n14135), 
            .ROA11(n14134), .ROA10(n14133), .ROA9(n14132), .ROA8(n14131), 
            .ROA7(n14130), .ROA6(n14129), .ROA5(n14128), .ROA4(n14127), 
            .ROA3(n14126), .ROA2(n14125), .ROA1(n14124), .ROA0(n14123), 
            .ROB17(n14158), .ROB16(n14157), .ROB15(n14156), .ROB14(n14155), 
            .ROB13(n14154), .ROB12(n14153), .ROB11(n14152), .ROB10(n14151), 
            .ROB9(n14150), .ROB8(n14149), .ROB7(n14148), .ROB6(n14147), 
            .ROB5(n14146), .ROB4(n14145), .ROB3(n14144), .ROB2(n14143), 
            .ROB1(n14142), .ROB0(n14141), .P35(n14195), .P34(n14194), 
            .P33(n14193), .P32(n14192), .P31(n14191), .P30(n14190), 
            .P29(n14189), .P28(n14188), .P27(n14187), .P26(n14186), 
            .P25(n14185), .P24(n14184), .P23(n14183), .P22(n14182), 
            .P21(n14181), .P20(n14180), .P19(n14179), .P18(n14178), 
            .P17(n14177), .P16(n14176), .P15(n14175), .P14(n14174), 
            .P13(n14173), .P12(n14172), .P11(n14171), .P10(n14170), 
            .P9(n14169), .P8(n14168), .P7(n14167), .P6(n14166), .P5(n14165), 
            .P4(n14164), .P3(n14163), .P2(n14162), .P1(n14161), .P0(n14160), 
            .SIGNEDP(n14159));
    defparam lat_mult_12.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTA_CE = "CE0";
    defparam lat_mult_12.REG_INPUTA_RST = "RST0";
    defparam lat_mult_12.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTB_CE = "CE0";
    defparam lat_mult_12.REG_INPUTB_RST = "RST0";
    defparam lat_mult_12.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTC_CE = "CE0";
    defparam lat_mult_12.REG_INPUTC_RST = "RST0";
    defparam lat_mult_12.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_12.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_12.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_12.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_12.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_12.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_12.CLK0_DIV = "ENABLED";
    defparam lat_mult_12.CLK1_DIV = "ENABLED";
    defparam lat_mult_12.CLK2_DIV = "ENABLED";
    defparam lat_mult_12.CLK3_DIV = "ENABLED";
    defparam lat_mult_12.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_12.GSR = "DISABLED";
    defparam lat_mult_12.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_12.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_12.MULT_BYPASS = "DISABLED";
    defparam lat_mult_12.RESETMODE = "SYNC";
    MULT18X18D lat_mult_11 (.A17(\rom4_w_i[12] ), .A16(\rom4_w_i[12] ), 
            .A15(\rom4_w_i[12] ), .A14(\rom4_w_i[12] ), .A13(\rom4_w_i[12] ), 
            .A12(\rom4_w_i[12] ), .A11(\rom4_w_i[12] ), .A10(\rom4_w_i[12] ), 
            .A9(\rom4_w_i[12] ), .A8(\rom4_w_i[12] ), .A7(GND_net), .A6(n34777), 
            .A5(GND_net), .A4(GND_net), .A3(n34777), .A2(GND_net), .A1(n34777), 
            .A0(n34777), .B17(n319), .B16(n319), .B15(n319), .B14(n319), 
            .B13(n319), .B12(n319), .B11(n319), .B10(n319), .B9(n319), 
            .B8(n319), .B7(n319), .B6(n319), .B5(n319), .B4(n319), 
            .B3(n319), .B2(n319), .B1(n319), .B0(n319), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n14067), .ROA16(n14066), .ROA15(n14065), 
            .ROA14(n14064), .ROA13(n14063), .ROA12(n14062), .ROA11(n14061), 
            .ROA10(n14060), .ROA9(n14059), .ROA8(n14058), .ROA7(n14057), 
            .ROA6(n14056), .ROA5(n14055), .ROA4(n14054), .ROA3(n14053), 
            .ROA2(n14052), .ROA1(n14051), .ROA0(n14050), .ROB17(n14085), 
            .ROB16(n14084), .ROB15(n14083), .ROB14(n14082), .ROB13(n14081), 
            .ROB12(n14080), .ROB11(n14079), .ROB10(n14078), .ROB9(n14077), 
            .ROB8(n14076), .ROB7(n14075), .ROB6(n14074), .ROB5(n14073), 
            .ROB4(n14072), .ROB3(n14071), .ROB2(n14070), .ROB1(n14069), 
            .ROB0(n14068), .P35(n14122), .P34(n14121), .P33(n14120), 
            .P32(n14119), .P31(n14118), .P30(n14117), .P29(n14116), 
            .P28(n14115), .P27(n14114), .P26(n14113), .P25(n14112), 
            .P24(n14111), .P23(n14110), .P22(n14109), .P21(n14108), 
            .P20(n14107), .P19(n14106), .P18(n14105), .P17(n14104), 
            .P16(n14103), .P15(n14102), .P14(n14101), .P13(n14100), 
            .P12(n14099), .P11(n14098), .P10(n14097), .P9(n14096), .P8(n14095), 
            .P7(n14094), .P6(n14093), .P5(n14092), .P4(n14091), .P3(n14090), 
            .P2(n14089), .P1(n14088), .P0(n14087), .SIGNEDP(n14086));
    defparam lat_mult_11.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTA_CE = "CE0";
    defparam lat_mult_11.REG_INPUTA_RST = "RST0";
    defparam lat_mult_11.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTB_CE = "CE0";
    defparam lat_mult_11.REG_INPUTB_RST = "RST0";
    defparam lat_mult_11.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTC_CE = "CE0";
    defparam lat_mult_11.REG_INPUTC_RST = "RST0";
    defparam lat_mult_11.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_11.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_11.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_11.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_11.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_11.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_11.CLK0_DIV = "ENABLED";
    defparam lat_mult_11.CLK1_DIV = "ENABLED";
    defparam lat_mult_11.CLK2_DIV = "ENABLED";
    defparam lat_mult_11.CLK3_DIV = "ENABLED";
    defparam lat_mult_11.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_11.GSR = "DISABLED";
    defparam lat_mult_11.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_11.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_11.MULT_BYPASS = "DISABLED";
    defparam lat_mult_11.RESETMODE = "SYNC";
    MULT18X18D lat_mult_10 (.A17(\rom4_w_i[12] ), .A16(\rom4_w_i[12] ), 
            .A15(\rom4_w_i[12] ), .A14(\rom4_w_i[12] ), .A13(\rom4_w_i[12] ), 
            .A12(\rom4_w_i[12] ), .A11(\rom4_w_i[12] ), .A10(\rom4_w_i[12] ), 
            .A9(\rom4_w_i[12] ), .A8(\rom4_w_i[12] ), .A7(\rom4_w_i[12] ), 
            .A6(\rom4_w_i[12] ), .A5(\rom4_w_i[12] ), .A4(\rom4_w_i[12] ), 
            .A3(\rom4_w_i[12] ), .A2(\rom4_w_i[12] ), .A1(\rom4_w_i[12] ), 
            .A0(\rom4_w_i[12] ), .B17(n10735), .B16(n10734), .B15(n10733), 
            .B14(n10732), .B13(n10731), .B12(n10730), .B11(n10729), 
            .B10(n10728), .B9(n10727), .B8(n10726), .B7(n10725), .B6(n10724), 
            .B5(n10723), .B4(n10722), .B3(n10721), .B2(n10720), .B1(n10719), 
            .B0(n10718), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n13994), 
            .ROA16(n13993), .ROA15(n13992), .ROA14(n13991), .ROA13(n13990), 
            .ROA12(n13989), .ROA11(n13988), .ROA10(n13987), .ROA9(n13986), 
            .ROA8(n13985), .ROA7(n13984), .ROA6(n13983), .ROA5(n13982), 
            .ROA4(n13981), .ROA3(n13980), .ROA2(n13979), .ROA1(n13978), 
            .ROA0(n13977), .ROB17(n14012), .ROB16(n14011), .ROB15(n14010), 
            .ROB14(n14009), .ROB13(n14008), .ROB12(n14007), .ROB11(n14006), 
            .ROB10(n14005), .ROB9(n14004), .ROB8(n14003), .ROB7(n14002), 
            .ROB6(n14001), .ROB5(n14000), .ROB4(n13999), .ROB3(n13998), 
            .ROB2(n13997), .ROB1(n13996), .ROB0(n13995), .P35(n14049), 
            .P34(n14048), .P33(n14047), .P32(n14046), .P31(n14045), 
            .P30(n14044), .P29(n14043), .P28(n14042), .P27(n14041), 
            .P26(n14040), .P25(n14039), .P24(n14038), .P23(n14037), 
            .P22(n14036), .P21(n14035), .P20(n14034), .P19(n14033), 
            .P18(n14032), .P17(n14031), .P16(n14030), .P15(n14029), 
            .P14(n14028), .P13(n14027), .P12(n14026), .P11(n14025), 
            .P10(n14024), .P9(n14023), .P8(n14022), .P7(n14021), .P6(n14020), 
            .P5(n14019), .P4(n14018), .P3(n14017), .P2(n14016), .P1(n14015), 
            .P0(n14014), .SIGNEDP(n14013));
    defparam lat_mult_10.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTA_CE = "CE0";
    defparam lat_mult_10.REG_INPUTA_RST = "RST0";
    defparam lat_mult_10.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTB_CE = "CE0";
    defparam lat_mult_10.REG_INPUTB_RST = "RST0";
    defparam lat_mult_10.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTC_CE = "CE0";
    defparam lat_mult_10.REG_INPUTC_RST = "RST0";
    defparam lat_mult_10.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_10.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_10.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_10.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_10.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_10.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_10.CLK0_DIV = "ENABLED";
    defparam lat_mult_10.CLK1_DIV = "ENABLED";
    defparam lat_mult_10.CLK2_DIV = "ENABLED";
    defparam lat_mult_10.CLK3_DIV = "ENABLED";
    defparam lat_mult_10.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_10.GSR = "DISABLED";
    defparam lat_mult_10.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_10.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_10.MULT_BYPASS = "DISABLED";
    defparam lat_mult_10.RESETMODE = "SYNC";
    MULT18X18D mult_972 (.A17(\rom4_w_i[12] ), .A16(\rom4_w_i[12] ), .A15(\rom4_w_i[12] ), 
            .A14(\rom4_w_i[12] ), .A13(\rom4_w_i[12] ), .A12(\rom4_w_i[12] ), 
            .A11(\rom4_w_i[12] ), .A10(\rom4_w_i[12] ), .A9(\rom4_w_i[12] ), 
            .A8(\rom4_w_i[12] ), .A7(GND_net), .A6(n34777), .A5(GND_net), 
            .A4(GND_net), .A3(n34777), .A2(GND_net), .A1(n34777), .A0(n34777), 
            .B17(n10735), .B16(n10734), .B15(n10733), .B14(n10732), 
            .B13(n10731), .B12(n10730), .B11(n10729), .B10(n10728), 
            .B9(n10727), .B8(n10726), .B7(n10725), .B6(n10724), .B5(n10723), 
            .B4(n10722), .B3(n10721), .B2(n10720), .B1(n10719), .B0(n10718), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n13921), .ROA16(n13920), 
            .ROA15(n13919), .ROA14(n13918), .ROA13(n13917), .ROA12(n13916), 
            .ROA11(n13915), .ROA10(n13914), .ROA9(n13913), .ROA8(n13912), 
            .ROA7(n13911), .ROA6(n13910), .ROA5(n13909), .ROA4(n13908), 
            .ROA3(n13907), .ROA2(n13906), .ROA1(n13905), .ROA0(n13904), 
            .ROB17(n13939), .ROB16(n13938), .ROB15(n13937), .ROB14(n13936), 
            .ROB13(n13935), .ROB12(n13934), .ROB11(n13933), .ROB10(n13932), 
            .ROB9(n13931), .ROB8(n13930), .ROB7(n13929), .ROB6(n13928), 
            .ROB5(n13927), .ROB4(n13926), .ROB3(n13925), .ROB2(n13924), 
            .ROB1(n13923), .ROB0(n13922), .P35(n13976), .P34(n13975), 
            .P33(n13974), .P32(n13973), .P31(n13972), .P30(n13971), 
            .P29(n13970), .P28(n13969), .P27(n13968), .P26(n13967), 
            .P25(n13966), .P24(n13965), .P23(n13964), .P22(n13963), 
            .P21(n13962), .P20(n13961), .P19(n13960), .P18(n13959), 
            .P17(n13958), .P16(n13957), .P15(n13956), .P14(n13955), 
            .P13(n13954), .P12(n13953), .P11(n13952), .P10(n13951), 
            .P9(n13950), .P8(n13949), .P7(n13948), .P6(n13947), .P5(n13946), 
            .P4(n13945), .P3(n13944), .P2(n13943), .P1(n13942), .P0(n13941), 
            .SIGNEDP(n13940));
    defparam mult_972.REG_INPUTA_CLK = "NONE";
    defparam mult_972.REG_INPUTA_CE = "CE0";
    defparam mult_972.REG_INPUTA_RST = "RST0";
    defparam mult_972.REG_INPUTB_CLK = "NONE";
    defparam mult_972.REG_INPUTB_CE = "CE0";
    defparam mult_972.REG_INPUTB_RST = "RST0";
    defparam mult_972.REG_INPUTC_CLK = "NONE";
    defparam mult_972.REG_INPUTC_CE = "CE0";
    defparam mult_972.REG_INPUTC_RST = "RST0";
    defparam mult_972.REG_PIPELINE_CLK = "NONE";
    defparam mult_972.REG_PIPELINE_CE = "CE0";
    defparam mult_972.REG_PIPELINE_RST = "RST0";
    defparam mult_972.REG_OUTPUT_CLK = "NONE";
    defparam mult_972.REG_OUTPUT_CE = "CE0";
    defparam mult_972.REG_OUTPUT_RST = "RST0";
    defparam mult_972.CLK0_DIV = "ENABLED";
    defparam mult_972.CLK1_DIV = "ENABLED";
    defparam mult_972.CLK2_DIV = "ENABLED";
    defparam mult_972.CLK3_DIV = "ENABLED";
    defparam mult_972.HIGHSPEED_CLK = "NONE";
    defparam mult_972.GSR = "DISABLED";
    defparam mult_972.CAS_MATCH_REG = "FALSE";
    defparam mult_972.SOURCEB_MODE = "B_SHIFT";
    defparam mult_972.MULT_BYPASS = "DISABLED";
    defparam mult_972.RESETMODE = "SYNC";
    MULT18X18D lat_mult_52 (.A17(\rom4_w_r[1] ), .A16(\rom4_w_r[1] ), .A15(\rom4_w_r[1] ), 
            .A14(\rom4_w_r[1] ), .A13(\rom4_w_r[1] ), .A12(\rom4_w_r[1] ), 
            .A11(\rom4_w_r[1] ), .A10(\rom4_w_r[1] ), .A9(\rom4_w_r[1] ), 
            .A8(\rom4_w_r[1] ), .A7(\rom4_w_r[1] ), .A6(\rom4_w_r[1] ), 
            .A5(\rom4_w_r[1] ), .A4(\rom4_w_r[1] ), .A3(\rom4_w_r[1] ), 
            .A2(\rom4_w_r[1] ), .A1(\rom4_w_r[1] ), .A0(\rom4_w_r[1] ), 
            .B17(n12264), .B16(n12264), .B15(n12264), .B14(n12264), 
            .B13(n12264), .B12(n12264), .B11(n12264), .B10(n12264), 
            .B9(n12264), .B8(n12264), .B7(n12264), .B6(n12264), .B5(n12263), 
            .B4(n12262), .B3(n12261), .B2(n12260), .B1(n12259), .B0(n12258), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n16942), .ROA16(n16941), 
            .ROA15(n16940), .ROA14(n16939), .ROA13(n16938), .ROA12(n16937), 
            .ROA11(n16936), .ROA10(n16935), .ROA9(n16934), .ROA8(n16933), 
            .ROA7(n16932), .ROA6(n16931), .ROA5(n16930), .ROA4(n16929), 
            .ROA3(n16928), .ROA2(n16927), .ROA1(n16926), .ROA0(n16925), 
            .ROB17(n16960), .ROB16(n16959), .ROB15(n16958), .ROB14(n16957), 
            .ROB13(n16956), .ROB12(n16955), .ROB11(n16954), .ROB10(n16953), 
            .ROB9(n16952), .ROB8(n16951), .ROB7(n16950), .ROB6(n16949), 
            .ROB5(n16948), .ROB4(n16947), .ROB3(n16946), .ROB2(n16945), 
            .ROB1(n16944), .ROB0(n16943), .P35(n16997), .P34(n16996), 
            .P33(n16995), .P32(n16994), .P31(n16993), .P30(n16992), 
            .P29(n16991), .P28(n16990), .P27(n16989), .P26(n16988), 
            .P25(n16987), .P24(n16986), .P23(n16985), .P22(n16984), 
            .P21(n16983), .P20(n16982), .P19(n16981), .P18(n16980), 
            .P17(n16979), .P16(n16978), .P15(n16977), .P14(n16976), 
            .P13(n16975), .P12(n16974), .P11(n16973), .P10(n16972), 
            .P9(n16971), .P8(n16970), .P7(n16969), .P6(n16968), .P5(n16967), 
            .P4(n16966), .P3(n16965), .P2(n16964), .P1(n16963), .P0(n16962), 
            .SIGNEDP(n16961));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_52.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_52.REG_INPUTA_CE = "CE0";
    defparam lat_mult_52.REG_INPUTA_RST = "RST0";
    defparam lat_mult_52.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_52.REG_INPUTB_CE = "CE0";
    defparam lat_mult_52.REG_INPUTB_RST = "RST0";
    defparam lat_mult_52.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_52.REG_INPUTC_CE = "CE0";
    defparam lat_mult_52.REG_INPUTC_RST = "RST0";
    defparam lat_mult_52.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_52.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_52.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_52.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_52.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_52.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_52.CLK0_DIV = "ENABLED";
    defparam lat_mult_52.CLK1_DIV = "ENABLED";
    defparam lat_mult_52.CLK2_DIV = "ENABLED";
    defparam lat_mult_52.CLK3_DIV = "ENABLED";
    defparam lat_mult_52.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_52.GSR = "DISABLED";
    defparam lat_mult_52.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_52.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_52.MULT_BYPASS = "DISABLED";
    defparam lat_mult_52.RESETMODE = "SYNC";
    MULT18X18D lat_mult_57 (.A17(shift_4_dout_i[23]), .A16(shift_4_dout_i[23]), 
            .A15(shift_4_dout_i[23]), .A14(shift_4_dout_i[23]), .A13(shift_4_dout_i[23]), 
            .A12(shift_4_dout_i[23]), .A11(shift_4_dout_i[23]), .A10(shift_4_dout_i[23]), 
            .A9(shift_4_dout_i[23]), .A8(shift_4_dout_i[23]), .A7(shift_4_dout_i[23]), 
            .A6(shift_4_dout_i[23]), .A5(shift_4_dout_i[23]), .A4(shift_4_dout_i[22]), 
            .A3(shift_4_dout_i[21]), .A2(shift_4_dout_i[20]), .A1(shift_4_dout_i[19]), 
            .A0(shift_4_dout_i[18]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n119), .B8(n119), .B7(n119), .B6(n119), .B5(n119), 
            .B4(n119), .B3(n119), .B2(n119), .B1(n119), .B0(n119), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17288), .ROA16(n17287), 
            .ROA15(n17286), .ROA14(n17285), .ROA13(n17284), .ROA12(n17283), 
            .ROA11(n17282), .ROA10(n17281), .ROA9(n17280), .ROA8(n17279), 
            .ROA7(n17278), .ROA6(n17277), .ROA5(n17276), .ROA4(n17275), 
            .ROA3(n17274), .ROA2(n17273), .ROA1(n17272), .ROA0(n17271), 
            .ROB17(n17306), .ROB16(n17305), .ROB15(n17304), .ROB14(n17303), 
            .ROB13(n17302), .ROB12(n17301), .ROB11(n17300), .ROB10(n17299), 
            .ROB9(n17298), .ROB8(n17297), .ROB7(n17296), .ROB6(n17295), 
            .ROB5(n17294), .ROB4(n17293), .ROB3(n17292), .ROB2(n17291), 
            .ROB1(n17290), .ROB0(n17289), .P35(n17343), .P34(n17342), 
            .P33(n17341), .P32(n17340), .P31(n17339), .P30(n17338), 
            .P29(n17337), .P28(n17336), .P27(n17335), .P26(n17334), 
            .P25(n17333), .P24(n17332), .P23(n17331), .P22(n17330), 
            .P21(n17329), .P20(n17328), .P19(n17327), .P18(n17326), 
            .P17(n17325), .P16(n17324), .P15(n17323), .P14(n17322), 
            .P13(n17321), .P12(n17320), .P11(n17319), .P10(n17318), 
            .P9(n17317), .P8(n17316), .P7(n17315), .P6(n17314), .P5(n17313), 
            .P4(n17312), .P3(n17311), .P2(n17310), .P1(n17309), .P0(n17308), 
            .SIGNEDP(n17307));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_57.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_57.REG_INPUTA_CE = "CE0";
    defparam lat_mult_57.REG_INPUTA_RST = "RST0";
    defparam lat_mult_57.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_57.REG_INPUTB_CE = "CE0";
    defparam lat_mult_57.REG_INPUTB_RST = "RST0";
    defparam lat_mult_57.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_57.REG_INPUTC_CE = "CE0";
    defparam lat_mult_57.REG_INPUTC_RST = "RST0";
    defparam lat_mult_57.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_57.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_57.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_57.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_57.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_57.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_57.CLK0_DIV = "ENABLED";
    defparam lat_mult_57.CLK1_DIV = "ENABLED";
    defparam lat_mult_57.CLK2_DIV = "ENABLED";
    defparam lat_mult_57.CLK3_DIV = "ENABLED";
    defparam lat_mult_57.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_57.GSR = "DISABLED";
    defparam lat_mult_57.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_57.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_57.MULT_BYPASS = "DISABLED";
    defparam lat_mult_57.RESETMODE = "SYNC";
    MULT18X18D lat_mult_50 (.A17(\rom4_w_r[1] ), .A16(\rom4_w_r[1] ), .A15(\rom4_w_r[1] ), 
            .A14(\rom4_w_r[1] ), .A13(\rom4_w_r[1] ), .A12(\rom4_w_r[1] ), 
            .A11(\rom4_w_r[1] ), .A10(\rom4_w_r[1] ), .A9(\rom4_w_r[1] ), 
            .A8(\rom4_w_r[1] ), .A7(\rom4_w_r[1] ), .A6(\rom4_w_r[1] ), 
            .A5(\rom4_w_r[1] ), .A4(\rom4_w_r[1] ), .A3(\rom4_w_r[1] ), 
            .A2(\rom4_w_r[1] ), .A1(\rom4_w_r[1] ), .A0(\rom4_w_r[1] ), 
            .B17(n12257), .B16(n12256), .B15(n12255), .B14(n12254), 
            .B13(n12253), .B12(n12252), .B11(n12251), .B10(n12250), 
            .B9(n12249), .B8(n12248), .B7(n12247), .B6(n12246), .B5(n12245), 
            .B4(n12244), .B3(n12243), .B2(n12242), .B1(n12241), .B0(n12240), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n16796), .ROA16(n16795), 
            .ROA15(n16794), .ROA14(n16793), .ROA13(n16792), .ROA12(n16791), 
            .ROA11(n16790), .ROA10(n16789), .ROA9(n16788), .ROA8(n16787), 
            .ROA7(n16786), .ROA6(n16785), .ROA5(n16784), .ROA4(n16783), 
            .ROA3(n16782), .ROA2(n16781), .ROA1(n16780), .ROA0(n16779), 
            .ROB17(n16814), .ROB16(n16813), .ROB15(n16812), .ROB14(n16811), 
            .ROB13(n16810), .ROB12(n16809), .ROB11(n16808), .ROB10(n16807), 
            .ROB9(n16806), .ROB8(n16805), .ROB7(n16804), .ROB6(n16803), 
            .ROB5(n16802), .ROB4(n16801), .ROB3(n16800), .ROB2(n16799), 
            .ROB1(n16798), .ROB0(n16797), .P35(n16851), .P34(n16850), 
            .P33(n16849), .P32(n16848), .P31(n16847), .P30(n16846), 
            .P29(n16845), .P28(n16844), .P27(n16843), .P26(n16842), 
            .P25(n16841), .P24(n16840), .P23(n16839), .P22(n16838), 
            .P21(n16837), .P20(n16836), .P19(n16835), .P18(n16834), 
            .P17(n16833), .P16(n16832), .P15(n16831), .P14(n16830), 
            .P13(n16829), .P12(n16828), .P11(n16827), .P10(n16826), 
            .P9(n16825), .P8(n16824), .P7(n16823), .P6(n16822), .P5(n16821), 
            .P4(n16820), .P3(n16819), .P2(n16818), .P1(n16817), .P0(n16816), 
            .SIGNEDP(n16815));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_50.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_50.REG_INPUTA_CE = "CE0";
    defparam lat_mult_50.REG_INPUTA_RST = "RST0";
    defparam lat_mult_50.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_50.REG_INPUTB_CE = "CE0";
    defparam lat_mult_50.REG_INPUTB_RST = "RST0";
    defparam lat_mult_50.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_50.REG_INPUTC_CE = "CE0";
    defparam lat_mult_50.REG_INPUTC_RST = "RST0";
    defparam lat_mult_50.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_50.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_50.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_50.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_50.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_50.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_50.CLK0_DIV = "ENABLED";
    defparam lat_mult_50.CLK1_DIV = "ENABLED";
    defparam lat_mult_50.CLK2_DIV = "ENABLED";
    defparam lat_mult_50.CLK3_DIV = "ENABLED";
    defparam lat_mult_50.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_50.GSR = "DISABLED";
    defparam lat_mult_50.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_50.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_50.MULT_BYPASS = "DISABLED";
    defparam lat_mult_50.RESETMODE = "SYNC";
    MULT18X18D lat_mult_55 (.A17(shift_4_dout_i[23]), .A16(shift_4_dout_i[23]), 
            .A15(shift_4_dout_i[23]), .A14(shift_4_dout_i[23]), .A13(shift_4_dout_i[23]), 
            .A12(shift_4_dout_i[23]), .A11(shift_4_dout_i[23]), .A10(shift_4_dout_i[23]), 
            .A9(shift_4_dout_i[23]), .A8(shift_4_dout_i[23]), .A7(shift_4_dout_i[23]), 
            .A6(shift_4_dout_i[23]), .A5(shift_4_dout_i[23]), .A4(shift_4_dout_i[22]), 
            .A3(shift_4_dout_i[21]), .A2(shift_4_dout_i[20]), .A1(shift_4_dout_i[19]), 
            .A0(shift_4_dout_i[18]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n12309), .B8(n12308), .B7(n12307), .B6(n12306), .B5(n12305), 
            .B4(n12304), .B3(n12303), .B2(n12302), .B1(n12301), .B0(n12300), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17142), .ROA16(n17141), 
            .ROA15(n17140), .ROA14(n17139), .ROA13(n17138), .ROA12(n17137), 
            .ROA11(n17136), .ROA10(n17135), .ROA9(n17134), .ROA8(n17133), 
            .ROA7(n17132), .ROA6(n17131), .ROA5(n17130), .ROA4(n17129), 
            .ROA3(n17128), .ROA2(n17127), .ROA1(n17126), .ROA0(n17125), 
            .ROB17(n17160), .ROB16(n17159), .ROB15(n17158), .ROB14(n17157), 
            .ROB13(n17156), .ROB12(n17155), .ROB11(n17154), .ROB10(n17153), 
            .ROB9(n17152), .ROB8(n17151), .ROB7(n17150), .ROB6(n17149), 
            .ROB5(n17148), .ROB4(n17147), .ROB3(n17146), .ROB2(n17145), 
            .ROB1(n17144), .ROB0(n17143), .P35(n17197), .P34(n17196), 
            .P33(n17195), .P32(n17194), .P31(n17193), .P30(n17192), 
            .P29(n17191), .P28(n17190), .P27(n17189), .P26(n17188), 
            .P25(n17187), .P24(n17186), .P23(n17185), .P22(n17184), 
            .P21(n17183), .P20(n17182), .P19(n17181), .P18(n17180), 
            .P17(n17179), .P16(n17178), .P15(n17177), .P14(n17176), 
            .P13(n17175), .P12(n17174), .P11(n17173), .P10(n17172), 
            .P9(n17171), .P8(n17170), .P7(n17169), .P6(n17168), .P5(n17167), 
            .P4(n17166), .P3(n17165), .P2(n17164), .P1(n17163), .P0(n17162), 
            .SIGNEDP(n17161));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_55.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_55.REG_INPUTA_CE = "CE0";
    defparam lat_mult_55.REG_INPUTA_RST = "RST0";
    defparam lat_mult_55.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_55.REG_INPUTB_CE = "CE0";
    defparam lat_mult_55.REG_INPUTB_RST = "RST0";
    defparam lat_mult_55.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_55.REG_INPUTC_CE = "CE0";
    defparam lat_mult_55.REG_INPUTC_RST = "RST0";
    defparam lat_mult_55.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_55.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_55.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_55.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_55.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_55.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_55.CLK0_DIV = "ENABLED";
    defparam lat_mult_55.CLK1_DIV = "ENABLED";
    defparam lat_mult_55.CLK2_DIV = "ENABLED";
    defparam lat_mult_55.CLK3_DIV = "ENABLED";
    defparam lat_mult_55.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_55.GSR = "DISABLED";
    defparam lat_mult_55.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_55.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_55.MULT_BYPASS = "DISABLED";
    defparam lat_mult_55.RESETMODE = "SYNC";
    MULT18X18D lat_mult_51 (.A17(\rom4_w_r[1] ), .A16(\rom4_w_r[1] ), .A15(\rom4_w_r[1] ), 
            .A14(\rom4_w_r[1] ), .A13(\rom4_w_r[1] ), .A12(\rom4_w_r[1] ), 
            .A11(\rom4_w_r[1] ), .A10(\rom4_w_r[1] ), .A9(\rom4_w_r[1] ), 
            .A8(\rom4_w_r[8] ), .A7(\rom4_w_r[5] ), .A6(\rom4_w_r[1] ), 
            .A5(\rom4_w_r[5] ), .A4(\rom4_w_r[5] ), .A3(\rom4_w_r[1] ), 
            .A2(\rom4_w_r[5] ), .A1(\rom4_w_r[1] ), .A0(n34777), .B17(n12264), 
            .B16(n12264), .B15(n12264), .B14(n12264), .B13(n12264), 
            .B12(n12264), .B11(n12264), .B10(n12264), .B9(n12264), .B8(n12264), 
            .B7(n12264), .B6(n12264), .B5(n12263), .B4(n12262), .B3(n12261), 
            .B2(n12260), .B1(n12259), .B0(n12258), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n16869), .ROA16(n16868), .ROA15(n16867), .ROA14(n16866), 
            .ROA13(n16865), .ROA12(n16864), .ROA11(n16863), .ROA10(n16862), 
            .ROA9(n16861), .ROA8(n16860), .ROA7(n16859), .ROA6(n16858), 
            .ROA5(n16857), .ROA4(n16856), .ROA3(n16855), .ROA2(n16854), 
            .ROA1(n16853), .ROA0(n16852), .ROB17(n16887), .ROB16(n16886), 
            .ROB15(n16885), .ROB14(n16884), .ROB13(n16883), .ROB12(n16882), 
            .ROB11(n16881), .ROB10(n16880), .ROB9(n16879), .ROB8(n16878), 
            .ROB7(n16877), .ROB6(n16876), .ROB5(n16875), .ROB4(n16874), 
            .ROB3(n16873), .ROB2(n16872), .ROB1(n16871), .ROB0(n16870), 
            .P35(n16924), .P34(n16923), .P33(n16922), .P32(n16921), 
            .P31(n16920), .P30(n16919), .P29(n16918), .P28(n16917), 
            .P27(n16916), .P26(n16915), .P25(n16914), .P24(n16913), 
            .P23(n16912), .P22(n16911), .P21(n16910), .P20(n16909), 
            .P19(n16908), .P18(n16907), .P17(n16906), .P16(n16905), 
            .P15(n16904), .P14(n16903), .P13(n16902), .P12(n16901), 
            .P11(n16900), .P10(n16899), .P9(n16898), .P8(n16897), .P7(n16896), 
            .P6(n16895), .P5(n16894), .P4(n16893), .P3(n16892), .P2(n16891), 
            .P1(n16890), .P0(n16889), .SIGNEDP(n16888));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_51.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_51.REG_INPUTA_CE = "CE0";
    defparam lat_mult_51.REG_INPUTA_RST = "RST0";
    defparam lat_mult_51.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_51.REG_INPUTB_CE = "CE0";
    defparam lat_mult_51.REG_INPUTB_RST = "RST0";
    defparam lat_mult_51.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_51.REG_INPUTC_CE = "CE0";
    defparam lat_mult_51.REG_INPUTC_RST = "RST0";
    defparam lat_mult_51.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_51.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_51.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_51.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_51.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_51.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_51.CLK0_DIV = "ENABLED";
    defparam lat_mult_51.CLK1_DIV = "ENABLED";
    defparam lat_mult_51.CLK2_DIV = "ENABLED";
    defparam lat_mult_51.CLK3_DIV = "ENABLED";
    defparam lat_mult_51.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_51.GSR = "DISABLED";
    defparam lat_mult_51.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_51.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_51.MULT_BYPASS = "DISABLED";
    defparam lat_mult_51.RESETMODE = "SYNC";
    MULT18X18D lat_mult_56 (.A17(shift_4_dout_i[17]), .A16(shift_4_dout_i[16]), 
            .A15(shift_4_dout_i[15]), .A14(shift_4_dout_i[14]), .A13(shift_4_dout_i[13]), 
            .A12(shift_4_dout_i[12]), .A11(shift_4_dout_i[11]), .A10(shift_4_dout_i[10]), 
            .A9(shift_4_dout_i[9]), .A8(shift_4_dout_i[8]), .A7(shift_4_dout_i[7]), 
            .A6(shift_4_dout_i[6]), .A5(shift_4_dout_i[5]), .A4(shift_4_dout_i[4]), 
            .A3(shift_4_dout_i[3]), .A2(shift_4_dout_i[2]), .A1(shift_4_dout_i[1]), 
            .A0(shift_4_dout_i[0]), .B17(n119), .B16(n119), .B15(n119), 
            .B14(n119), .B13(n119), .B12(n119), .B11(n119), .B10(n119), 
            .B9(n119), .B8(n119), .B7(n119), .B6(n119), .B5(n119), 
            .B4(n119), .B3(n119), .B2(n119), .B1(n119), .B0(n119), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n17215), .ROA16(n17214), 
            .ROA15(n17213), .ROA14(n17212), .ROA13(n17211), .ROA12(n17210), 
            .ROA11(n17209), .ROA10(n17208), .ROA9(n17207), .ROA8(n17206), 
            .ROA7(n17205), .ROA6(n17204), .ROA5(n17203), .ROA4(n17202), 
            .ROA3(n17201), .ROA2(n17200), .ROA1(n17199), .ROA0(n17198), 
            .ROB17(n17233), .ROB16(n17232), .ROB15(n17231), .ROB14(n17230), 
            .ROB13(n17229), .ROB12(n17228), .ROB11(n17227), .ROB10(n17226), 
            .ROB9(n17225), .ROB8(n17224), .ROB7(n17223), .ROB6(n17222), 
            .ROB5(n17221), .ROB4(n17220), .ROB3(n17219), .ROB2(n17218), 
            .ROB1(n17217), .ROB0(n17216), .P35(n17270), .P34(n17269), 
            .P33(n17268), .P32(n17267), .P31(n17266), .P30(n17265), 
            .P29(n17264), .P28(n17263), .P27(n17262), .P26(n17261), 
            .P25(n17260), .P24(n17259), .P23(n17258), .P22(n17257), 
            .P21(n17256), .P20(n17255), .P19(n17254), .P18(n17253), 
            .P17(n17252), .P16(n17251), .P15(n17250), .P14(n17249), 
            .P13(n17248), .P12(n17247), .P11(n17246), .P10(n17245), 
            .P9(n17244), .P8(n17243), .P7(n17242), .P6(n17241), .P5(n17240), 
            .P4(n17239), .P3(n17238), .P2(n17237), .P1(n17236), .P0(n17235), 
            .SIGNEDP(n17234));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_56.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_56.REG_INPUTA_CE = "CE0";
    defparam lat_mult_56.REG_INPUTA_RST = "RST0";
    defparam lat_mult_56.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_56.REG_INPUTB_CE = "CE0";
    defparam lat_mult_56.REG_INPUTB_RST = "RST0";
    defparam lat_mult_56.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_56.REG_INPUTC_CE = "CE0";
    defparam lat_mult_56.REG_INPUTC_RST = "RST0";
    defparam lat_mult_56.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_56.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_56.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_56.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_56.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_56.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_56.CLK0_DIV = "ENABLED";
    defparam lat_mult_56.CLK1_DIV = "ENABLED";
    defparam lat_mult_56.CLK2_DIV = "ENABLED";
    defparam lat_mult_56.CLK3_DIV = "ENABLED";
    defparam lat_mult_56.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_56.GSR = "DISABLED";
    defparam lat_mult_56.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_56.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_56.MULT_BYPASS = "DISABLED";
    defparam lat_mult_56.RESETMODE = "SYNC";
    LUT4 i20_3_lut_4_lut (.A(op_i_23__N_1154[18]), .B(n34841), .C(n30179), 
         .D(\delay_i_23__N_1202[18] ), .Z(\dout_i_23__N_5777[18] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_200 (.A(op_i_23__N_1154[2]), .B(n34841), .C(n30179), 
         .D(\delay_i_23__N_1202[2] ), .Z(\dout_i_23__N_5777[2] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_200.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_201 (.A(op_i_23__N_1154[1]), .B(n34841), .C(n30179), 
         .D(\delay_i_23__N_1202[1] ), .Z(\dout_i_23__N_5777[1] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_201.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_202 (.A(op_i_23__N_1154[0]), .B(n34841), .C(n30179), 
         .D(\delay_i_23__N_1202[0] ), .Z(\dout_i_23__N_5777[0] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_202.init = 16'h8f80;
    LUT4 i1_2_lut_rep_248_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[12]), 
         .Z(n34610)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_248_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_247_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[13]), 
         .Z(n34609)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_247_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_214_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[22]), 
         .Z(n34576)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_214_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_213_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[23]), 
         .Z(n34575)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_213_3_lut.init = 16'h6060;
    LUT4 i12552_2_lut_rep_328_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[0]), 
         .Z(n34690)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12552_2_lut_rep_328_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_250_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[10]), 
         .Z(n34612)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_250_3_lut.init = 16'h6060;
    LUT4 i227_2_lut_rep_387_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(valid), 
         .Z(clk_c_enable_1396)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i227_2_lut_rep_387_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_rep_259_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[11]), 
         .Z(n34621)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_259_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_303_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[7]), 
         .Z(n34665)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_303_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_231_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[17]), 
         .Z(n34593)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_231_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_216_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[22]), 
         .Z(n34578)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_216_3_lut.init = 16'h6060;
    LUT4 i20_3_lut_4_lut_adj_203 (.A(op_r_23__N_1106[0]), .B(n34841), .C(n30179), 
         .D(\delay_r_23__N_1178[0] ), .Z(\dout_r_23__N_5681[0] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_203.init = 16'h8f80;
    LUT4 i1_2_lut_rep_262_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[8]), 
         .Z(n34624)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_262_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_217_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[21]), 
         .Z(n34579)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_217_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_225_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[17]), 
         .Z(n34587)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_225_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_226_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[16]), 
         .Z(n34588)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_226_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_304_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[6]), 
         .Z(n34666)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_304_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_232_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[16]), 
         .Z(n34594)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_232_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_260_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[10]), 
         .Z(n34622)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_260_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_215_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[23]), 
         .Z(n34577)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_215_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_261_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[9]), 
         .Z(n34623)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_261_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_249_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[11]), 
         .Z(n34611)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_249_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_327_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[1]), 
         .Z(n34689)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_327_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_271_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[9]), 
         .Z(n34633)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_271_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_218_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[20]), 
         .Z(n34580)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_218_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_272_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[8]), 
         .Z(n34634)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_272_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_219_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[21]), 
         .Z(n34581)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_219_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_273_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[7]), 
         .Z(n34635)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_273_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_220_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[20]), 
         .Z(n34582)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_220_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_274_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[6]), 
         .Z(n34636)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_274_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_221_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[19]), 
         .Z(n34583)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_221_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_283_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[5]), 
         .Z(n34645)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_283_3_lut.init = 16'h6060;
    LUT4 i12957_2_lut_rep_222_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[18]), 
         .Z(n34584)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12957_2_lut_rep_222_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_284_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[4]), 
         .Z(n34646)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_284_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_223_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[19]), 
         .Z(n34585)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_223_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_293_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[3]), 
         .Z(n34655)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_293_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_224_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[18]), 
         .Z(n34586)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_224_3_lut.init = 16'h6060;
    LUT4 i12941_2_lut_rep_294_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[2]), 
         .Z(n34656)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12941_2_lut_rep_294_3_lut.init = 16'h6060;
    LUT4 i12940_2_lut_rep_305_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[1]), 
         .Z(n34667)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12940_2_lut_rep_305_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_233_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[15]), 
         .Z(n34595)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_233_3_lut.init = 16'h6060;
    LUT4 i12553_2_lut_rep_306_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[0]), 
         .Z(n34668)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12553_2_lut_rep_306_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_234_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[14]), 
         .Z(n34596)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_234_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_311_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[5]), 
         .Z(n34673)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_311_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_239_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[15]), 
         .Z(n34601)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_239_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_312_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[4]), 
         .Z(n34674)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_312_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_240_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[14]), 
         .Z(n34602)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_240_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_317_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[3]), 
         .Z(n34679)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_317_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_241_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[13]), 
         .Z(n34603)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_241_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_242_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_i_23__N_1154[12]), 
         .Z(n34604)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_242_3_lut.init = 16'h6060;
    LUT4 i1_2_lut_rep_318_3_lut (.A(\rom4_state[0] ), .B(n34799), .C(op_r_23__N_1106[2]), 
         .Z(n34680)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i1_2_lut_rep_318_3_lut.init = 16'h6060;
    
endmodule
//
// Verilog Description of module shift_2
//

module shift_2 (shift_2_dout_r, clk_c, clk_c_enable_1396, \dout_i_23__N_5777[0] , 
            \dout_r_23__N_5681[0] , valid, clk_c_enable_2299, VCC_net, 
            \dout_i_23__N_5777[1] , \dout_i_23__N_5777[2] , \dout_i_23__N_5777[3] , 
            \dout_i_23__N_5777[4] , \dout_i_23__N_5777[5] , \dout_i_23__N_5777[6] , 
            \dout_i_23__N_5777[7] , \dout_i_23__N_5777[8] , \dout_i_23__N_5777[9] , 
            \dout_i_23__N_5777[10] , \dout_i_23__N_5777[11] , \dout_i_23__N_5777[12] , 
            \dout_i_23__N_5777[13] , \dout_i_23__N_5777[14] , \dout_i_23__N_5777[15] , 
            \dout_i_23__N_5777[16] , \dout_i_23__N_5777[17] , \dout_i_23__N_5777[18] , 
            \dout_i_23__N_5777[19] , \dout_i_23__N_5777[20] , \dout_i_23__N_5777[21] , 
            \dout_i_23__N_5777[22] , \dout_i_23__N_5777[23] , \dout_r_23__N_5681[1] , 
            \dout_r_23__N_5681[2] , \dout_r_23__N_5681[3] , \dout_r_23__N_5681[4] , 
            \dout_r_23__N_5681[5] , \dout_r_23__N_5681[6] , \dout_r_23__N_5681[7] , 
            \dout_r_23__N_5681[8] , \dout_r_23__N_5681[9] , \dout_r_23__N_5681[10] , 
            \dout_r_23__N_5681[11] , \dout_r_23__N_5681[12] , \dout_r_23__N_5681[13] , 
            \dout_r_23__N_5681[14] , \dout_r_23__N_5681[15] , \dout_r_23__N_5681[16] , 
            \dout_r_23__N_5681[17] , \dout_r_23__N_5681[18] , \dout_r_23__N_5681[19] , 
            \dout_r_23__N_5681[20] , \dout_r_23__N_5681[21] , \dout_r_23__N_5681[22] , 
            \dout_r_23__N_5681[23] , n34841, shift_2_dout_i) /* synthesis syn_module_defined=1 */ ;
    output [23:0]shift_2_dout_r;
    input clk_c;
    input clk_c_enable_1396;
    input \dout_i_23__N_5777[0] ;
    input \dout_r_23__N_5681[0] ;
    output valid;
    input clk_c_enable_2299;
    input VCC_net;
    input \dout_i_23__N_5777[1] ;
    input \dout_i_23__N_5777[2] ;
    input \dout_i_23__N_5777[3] ;
    input \dout_i_23__N_5777[4] ;
    input \dout_i_23__N_5777[5] ;
    input \dout_i_23__N_5777[6] ;
    input \dout_i_23__N_5777[7] ;
    input \dout_i_23__N_5777[8] ;
    input \dout_i_23__N_5777[9] ;
    input \dout_i_23__N_5777[10] ;
    input \dout_i_23__N_5777[11] ;
    input \dout_i_23__N_5777[12] ;
    input \dout_i_23__N_5777[13] ;
    input \dout_i_23__N_5777[14] ;
    input \dout_i_23__N_5777[15] ;
    input \dout_i_23__N_5777[16] ;
    input \dout_i_23__N_5777[17] ;
    input \dout_i_23__N_5777[18] ;
    input \dout_i_23__N_5777[19] ;
    input \dout_i_23__N_5777[20] ;
    input \dout_i_23__N_5777[21] ;
    input \dout_i_23__N_5777[22] ;
    input \dout_i_23__N_5777[23] ;
    input \dout_r_23__N_5681[1] ;
    input \dout_r_23__N_5681[2] ;
    input \dout_r_23__N_5681[3] ;
    input \dout_r_23__N_5681[4] ;
    input \dout_r_23__N_5681[5] ;
    input \dout_r_23__N_5681[6] ;
    input \dout_r_23__N_5681[7] ;
    input \dout_r_23__N_5681[8] ;
    input \dout_r_23__N_5681[9] ;
    input \dout_r_23__N_5681[10] ;
    input \dout_r_23__N_5681[11] ;
    input \dout_r_23__N_5681[12] ;
    input \dout_r_23__N_5681[13] ;
    input \dout_r_23__N_5681[14] ;
    input \dout_r_23__N_5681[15] ;
    input \dout_r_23__N_5681[16] ;
    input \dout_r_23__N_5681[17] ;
    input \dout_r_23__N_5681[18] ;
    input \dout_r_23__N_5681[19] ;
    input \dout_r_23__N_5681[20] ;
    input \dout_r_23__N_5681[21] ;
    input \dout_r_23__N_5681[22] ;
    input \dout_r_23__N_5681[23] ;
    input n34841;
    output [23:0]shift_2_dout_i;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire n29860, n29859;
    wire [47:0]dout_i_23__N_5777;
    wire [47:0]dout_r_23__N_5681;
    
    wire n29858, n29857, n29856, n29855, n29854, n29853, n29852, 
        n29851, n29850, n29849, n29848, n29847, n29861, n29862, 
        n29863, n29864, n29865, n29866, n29867, n29868, n29869, 
        n29870, n30016, n30017, n30018, n30019, n30020, n30021, 
        n30022, n30023, n30024, n30025, n30026, n30027, n30028, 
        n30029, n30030, n30031, n30032, n30033, n30034, n30035, 
        n30036, n30037, n30038, n30039;
    
    FD1S3AX shift_reg_r_i0_i34 (.D(n29860), .CK(clk_c), .Q(shift_2_dout_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i34.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i35 (.D(n29859), .CK(clk_c), .Q(shift_2_dout_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i35.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i0 (.D(\dout_i_23__N_5777[0] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i0.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i0 (.D(\dout_r_23__N_5681[0] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i0.GSR = "ENABLED";
    FD1P3AX valid_26 (.D(VCC_net), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam valid_26.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i36 (.D(n29858), .CK(clk_c), .Q(shift_2_dout_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i36.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i37 (.D(n29857), .CK(clk_c), .Q(shift_2_dout_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i37.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i38 (.D(n29856), .CK(clk_c), .Q(shift_2_dout_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i38.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i39 (.D(n29855), .CK(clk_c), .Q(shift_2_dout_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i39.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i40 (.D(n29854), .CK(clk_c), .Q(shift_2_dout_r[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i40.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i41 (.D(n29853), .CK(clk_c), .Q(shift_2_dout_r[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i41.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i42 (.D(n29852), .CK(clk_c), .Q(shift_2_dout_r[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i42.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i43 (.D(n29851), .CK(clk_c), .Q(shift_2_dout_r[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i43.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i44 (.D(n29850), .CK(clk_c), .Q(shift_2_dout_r[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i44.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i45 (.D(n29849), .CK(clk_c), .Q(shift_2_dout_r[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i45.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i46 (.D(n29848), .CK(clk_c), .Q(shift_2_dout_r[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i46.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i47 (.D(n29847), .CK(clk_c), .Q(shift_2_dout_r[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i47.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i1 (.D(\dout_i_23__N_5777[1] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i1.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i2 (.D(\dout_i_23__N_5777[2] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i2.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i3 (.D(\dout_i_23__N_5777[3] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i3.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i4 (.D(\dout_i_23__N_5777[4] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i4.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i5 (.D(\dout_i_23__N_5777[5] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i5.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i6 (.D(\dout_i_23__N_5777[6] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i6.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i7 (.D(\dout_i_23__N_5777[7] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i7.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i8 (.D(\dout_i_23__N_5777[8] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i8.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i9 (.D(\dout_i_23__N_5777[9] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i9.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i10 (.D(\dout_i_23__N_5777[10] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i10.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i11 (.D(\dout_i_23__N_5777[11] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i11.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i12 (.D(\dout_i_23__N_5777[12] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i12.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i13 (.D(\dout_i_23__N_5777[13] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i13.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i14 (.D(\dout_i_23__N_5777[14] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i14.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i15 (.D(\dout_i_23__N_5777[15] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i15.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i16 (.D(\dout_i_23__N_5777[16] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i16.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i17 (.D(\dout_i_23__N_5777[17] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i17.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i18 (.D(\dout_i_23__N_5777[18] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i18.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i19 (.D(\dout_i_23__N_5777[19] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i19.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i20 (.D(\dout_i_23__N_5777[20] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i20.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i21 (.D(\dout_i_23__N_5777[21] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i21.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i22 (.D(\dout_i_23__N_5777[22] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i22.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i23 (.D(\dout_i_23__N_5777[23] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_i_23__N_5777[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i23.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i1 (.D(\dout_r_23__N_5681[1] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i1.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i2 (.D(\dout_r_23__N_5681[2] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i2.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i3 (.D(\dout_r_23__N_5681[3] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i3.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i4 (.D(\dout_r_23__N_5681[4] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i4.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i5 (.D(\dout_r_23__N_5681[5] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i5.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i6 (.D(\dout_r_23__N_5681[6] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i6.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i7 (.D(\dout_r_23__N_5681[7] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i7.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i8 (.D(\dout_r_23__N_5681[8] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i8.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i9 (.D(\dout_r_23__N_5681[9] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i9.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i10 (.D(\dout_r_23__N_5681[10] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i10.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i11 (.D(\dout_r_23__N_5681[11] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i11.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i12 (.D(\dout_r_23__N_5681[12] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i12.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i13 (.D(\dout_r_23__N_5681[13] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i13.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i14 (.D(\dout_r_23__N_5681[14] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i14.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i15 (.D(\dout_r_23__N_5681[15] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i15.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i16 (.D(\dout_r_23__N_5681[16] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i16.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i17 (.D(\dout_r_23__N_5681[17] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i17.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i18 (.D(\dout_r_23__N_5681[18] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i18.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i19 (.D(\dout_r_23__N_5681[19] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i19.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i20 (.D(\dout_r_23__N_5681[20] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i20.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i21 (.D(\dout_r_23__N_5681[21] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i21.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i22 (.D(\dout_r_23__N_5681[22] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i22.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i23 (.D(\dout_r_23__N_5681[23] ), .SP(clk_c_enable_1396), 
            .CK(clk_c), .Q(dout_r_23__N_5681[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i23.GSR = "ENABLED";
    LUT4 i12151_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[33]), 
         .D(shift_2_dout_r[9]), .Z(n29861)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12151_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12152_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[32]), 
         .D(shift_2_dout_r[8]), .Z(n29862)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12152_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12153_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[31]), 
         .D(shift_2_dout_r[7]), .Z(n29863)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12153_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12154_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[30]), 
         .D(shift_2_dout_r[6]), .Z(n29864)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12154_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12155_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[29]), 
         .D(shift_2_dout_r[5]), .Z(n29865)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12155_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12156_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[28]), 
         .D(shift_2_dout_r[4]), .Z(n29866)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12156_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12157_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[27]), 
         .D(shift_2_dout_r[3]), .Z(n29867)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12157_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12158_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[26]), 
         .D(shift_2_dout_r[2]), .Z(n29868)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12158_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12159_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[25]), 
         .D(shift_2_dout_r[1]), .Z(n29869)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12159_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12160_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[24]), 
         .D(shift_2_dout_r[0]), .Z(n29870)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12160_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12306_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[47]), 
         .D(shift_2_dout_i[23]), .Z(n30016)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12306_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12307_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[46]), 
         .D(shift_2_dout_i[22]), .Z(n30017)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12307_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12308_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[45]), 
         .D(shift_2_dout_i[21]), .Z(n30018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12308_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12309_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[44]), 
         .D(shift_2_dout_i[20]), .Z(n30019)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12309_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12310_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[43]), 
         .D(shift_2_dout_i[19]), .Z(n30020)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12310_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12311_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[42]), 
         .D(shift_2_dout_i[18]), .Z(n30021)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12311_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12312_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[41]), 
         .D(shift_2_dout_i[17]), .Z(n30022)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12312_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12313_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[40]), 
         .D(shift_2_dout_i[16]), .Z(n30023)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12313_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12314_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[39]), 
         .D(shift_2_dout_i[15]), .Z(n30024)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12314_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12315_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[38]), 
         .D(shift_2_dout_i[14]), .Z(n30025)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12315_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12316_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[37]), 
         .D(shift_2_dout_i[13]), .Z(n30026)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12316_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12317_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[36]), 
         .D(shift_2_dout_i[12]), .Z(n30027)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12317_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12318_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[35]), 
         .D(shift_2_dout_i[11]), .Z(n30028)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12318_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12319_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[34]), 
         .D(shift_2_dout_i[10]), .Z(n30029)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12319_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12320_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[33]), 
         .D(shift_2_dout_i[9]), .Z(n30030)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12320_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12321_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[32]), 
         .D(shift_2_dout_i[8]), .Z(n30031)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12321_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12322_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[31]), 
         .D(shift_2_dout_i[7]), .Z(n30032)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12322_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12323_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[30]), 
         .D(shift_2_dout_i[6]), .Z(n30033)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12323_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12324_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[29]), 
         .D(shift_2_dout_i[5]), .Z(n30034)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12324_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12325_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[28]), 
         .D(shift_2_dout_i[4]), .Z(n30035)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12325_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12326_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[27]), 
         .D(shift_2_dout_i[3]), .Z(n30036)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12326_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12327_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[26]), 
         .D(shift_2_dout_i[2]), .Z(n30037)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12327_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12328_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[25]), 
         .D(shift_2_dout_i[1]), .Z(n30038)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12328_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12329_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_i_23__N_5777[24]), 
         .D(shift_2_dout_i[0]), .Z(n30039)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12329_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12137_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[47]), 
         .D(shift_2_dout_r[23]), .Z(n29847)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12137_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12138_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[46]), 
         .D(shift_2_dout_r[22]), .Z(n29848)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12138_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12139_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[45]), 
         .D(shift_2_dout_r[21]), .Z(n29849)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12139_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12140_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[44]), 
         .D(shift_2_dout_r[20]), .Z(n29850)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12140_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12141_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[43]), 
         .D(shift_2_dout_r[19]), .Z(n29851)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12141_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12142_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[42]), 
         .D(shift_2_dout_r[18]), .Z(n29852)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12142_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12143_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[41]), 
         .D(shift_2_dout_r[17]), .Z(n29853)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12143_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12144_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[40]), 
         .D(shift_2_dout_r[16]), .Z(n29854)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12144_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12145_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[39]), 
         .D(shift_2_dout_r[15]), .Z(n29855)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12145_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12146_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[38]), 
         .D(shift_2_dout_r[14]), .Z(n29856)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12146_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12147_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[37]), 
         .D(shift_2_dout_r[13]), .Z(n29857)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12147_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12148_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[36]), 
         .D(shift_2_dout_r[12]), .Z(n29858)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12148_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12149_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[35]), 
         .D(shift_2_dout_r[11]), .Z(n29859)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12149_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12150_3_lut_4_lut (.A(valid), .B(n34841), .C(dout_r_23__N_5681[34]), 
         .D(shift_2_dout_r[10]), .Z(n29860)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(41[14] 46[8])
    defparam i12150_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX shift_reg_i_i0_i24 (.D(n30039), .CK(clk_c), .Q(shift_2_dout_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i24.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i25 (.D(n30038), .CK(clk_c), .Q(shift_2_dout_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i25.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i26 (.D(n30037), .CK(clk_c), .Q(shift_2_dout_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i26.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i27 (.D(n30036), .CK(clk_c), .Q(shift_2_dout_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i27.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i28 (.D(n30035), .CK(clk_c), .Q(shift_2_dout_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i28.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i29 (.D(n30034), .CK(clk_c), .Q(shift_2_dout_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i29.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i30 (.D(n30033), .CK(clk_c), .Q(shift_2_dout_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i30.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i31 (.D(n30032), .CK(clk_c), .Q(shift_2_dout_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i31.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i32 (.D(n30031), .CK(clk_c), .Q(shift_2_dout_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i32.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i33 (.D(n30030), .CK(clk_c), .Q(shift_2_dout_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i33.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i34 (.D(n30029), .CK(clk_c), .Q(shift_2_dout_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i34.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i35 (.D(n30028), .CK(clk_c), .Q(shift_2_dout_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i35.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i36 (.D(n30027), .CK(clk_c), .Q(shift_2_dout_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i36.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i37 (.D(n30026), .CK(clk_c), .Q(shift_2_dout_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i37.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i38 (.D(n30025), .CK(clk_c), .Q(shift_2_dout_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i38.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i39 (.D(n30024), .CK(clk_c), .Q(shift_2_dout_i[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i39.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i40 (.D(n30023), .CK(clk_c), .Q(shift_2_dout_i[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i40.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i41 (.D(n30022), .CK(clk_c), .Q(shift_2_dout_i[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i41.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i42 (.D(n30021), .CK(clk_c), .Q(shift_2_dout_i[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i42.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i43 (.D(n30020), .CK(clk_c), .Q(shift_2_dout_i[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i43.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i44 (.D(n30019), .CK(clk_c), .Q(shift_2_dout_i[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i44.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i45 (.D(n30018), .CK(clk_c), .Q(shift_2_dout_i[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i45.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i46 (.D(n30017), .CK(clk_c), .Q(shift_2_dout_i[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i46.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i47 (.D(n30016), .CK(clk_c), .Q(shift_2_dout_i[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_i_i0_i47.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i24 (.D(n29870), .CK(clk_c), .Q(shift_2_dout_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i24.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i25 (.D(n29869), .CK(clk_c), .Q(shift_2_dout_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i25.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i26 (.D(n29868), .CK(clk_c), .Q(shift_2_dout_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i26.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i27 (.D(n29867), .CK(clk_c), .Q(shift_2_dout_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i27.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i28 (.D(n29866), .CK(clk_c), .Q(shift_2_dout_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i28.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i29 (.D(n29865), .CK(clk_c), .Q(shift_2_dout_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i29.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i30 (.D(n29864), .CK(clk_c), .Q(shift_2_dout_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i30.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i31 (.D(n29863), .CK(clk_c), .Q(shift_2_dout_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i31.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i32 (.D(n29862), .CK(clk_c), .Q(shift_2_dout_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i32.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i33 (.D(n29861), .CK(clk_c), .Q(shift_2_dout_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=198, LSE_RLINE=205 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_2.v(36[5] 46[8])
    defparam shift_reg_r_i0_i33.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module shift_4
//

module shift_4 (clk_c, clk_c_enable_1373, \dout_r_23__N_5203[0] , \dout_i_23__N_5395[0] , 
            valid, clk_c_enable_2305, VCC_net, \dout_r_23__N_5203[1] , 
            \dout_r_23__N_5203[2] , \dout_r_23__N_5203[3] , \dout_r_23__N_5203[4] , 
            \dout_r_23__N_5203[5] , \dout_r_23__N_5203[6] , \dout_r_23__N_5203[7] , 
            \dout_r_23__N_5203[8] , \dout_r_23__N_5203[9] , \dout_r_23__N_5203[10] , 
            \dout_r_23__N_5203[11] , \dout_r_23__N_5203[12] , \dout_r_23__N_5203[13] , 
            \dout_r_23__N_5203[14] , \dout_r_23__N_5203[15] , \dout_r_23__N_5203[16] , 
            \dout_r_23__N_5203[17] , \dout_r_23__N_5203[18] , \dout_r_23__N_5203[19] , 
            \dout_r_23__N_5203[20] , \dout_r_23__N_5203[21] , \dout_r_23__N_5203[22] , 
            \dout_r_23__N_5203[23] , \dout_i_23__N_5395[1] , \dout_i_23__N_5395[2] , 
            \dout_i_23__N_5395[3] , \dout_i_23__N_5395[4] , \dout_i_23__N_5395[5] , 
            \dout_i_23__N_5395[6] , \dout_i_23__N_5395[7] , \dout_i_23__N_5395[8] , 
            \dout_i_23__N_5395[9] , \dout_i_23__N_5395[10] , \dout_i_23__N_5395[11] , 
            \dout_i_23__N_5395[12] , \dout_i_23__N_5395[13] , \dout_i_23__N_5395[14] , 
            \dout_i_23__N_5395[15] , \dout_i_23__N_5395[16] , \dout_i_23__N_5395[17] , 
            \dout_i_23__N_5395[18] , \dout_i_23__N_5395[19] , \dout_i_23__N_5395[20] , 
            \dout_i_23__N_5395[21] , \dout_i_23__N_5395[22] , \dout_i_23__N_5395[23] , 
            n34842, shift_4_dout_r, shift_4_dout_i) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input clk_c_enable_1373;
    input \dout_r_23__N_5203[0] ;
    input \dout_i_23__N_5395[0] ;
    output valid;
    input clk_c_enable_2305;
    input VCC_net;
    input \dout_r_23__N_5203[1] ;
    input \dout_r_23__N_5203[2] ;
    input \dout_r_23__N_5203[3] ;
    input \dout_r_23__N_5203[4] ;
    input \dout_r_23__N_5203[5] ;
    input \dout_r_23__N_5203[6] ;
    input \dout_r_23__N_5203[7] ;
    input \dout_r_23__N_5203[8] ;
    input \dout_r_23__N_5203[9] ;
    input \dout_r_23__N_5203[10] ;
    input \dout_r_23__N_5203[11] ;
    input \dout_r_23__N_5203[12] ;
    input \dout_r_23__N_5203[13] ;
    input \dout_r_23__N_5203[14] ;
    input \dout_r_23__N_5203[15] ;
    input \dout_r_23__N_5203[16] ;
    input \dout_r_23__N_5203[17] ;
    input \dout_r_23__N_5203[18] ;
    input \dout_r_23__N_5203[19] ;
    input \dout_r_23__N_5203[20] ;
    input \dout_r_23__N_5203[21] ;
    input \dout_r_23__N_5203[22] ;
    input \dout_r_23__N_5203[23] ;
    input \dout_i_23__N_5395[1] ;
    input \dout_i_23__N_5395[2] ;
    input \dout_i_23__N_5395[3] ;
    input \dout_i_23__N_5395[4] ;
    input \dout_i_23__N_5395[5] ;
    input \dout_i_23__N_5395[6] ;
    input \dout_i_23__N_5395[7] ;
    input \dout_i_23__N_5395[8] ;
    input \dout_i_23__N_5395[9] ;
    input \dout_i_23__N_5395[10] ;
    input \dout_i_23__N_5395[11] ;
    input \dout_i_23__N_5395[12] ;
    input \dout_i_23__N_5395[13] ;
    input \dout_i_23__N_5395[14] ;
    input \dout_i_23__N_5395[15] ;
    input \dout_i_23__N_5395[16] ;
    input \dout_i_23__N_5395[17] ;
    input \dout_i_23__N_5395[18] ;
    input \dout_i_23__N_5395[19] ;
    input \dout_i_23__N_5395[20] ;
    input \dout_i_23__N_5395[21] ;
    input \dout_i_23__N_5395[22] ;
    input \dout_i_23__N_5395[23] ;
    input n34842;
    output [23:0]shift_4_dout_r;
    output [23:0]shift_4_dout_i;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    wire [95:0]dout_i_23__N_5395;
    wire [95:0]dout_r_23__N_5203;
    
    wire n30043, n30044, n30045, n30046, n30047, n30048, n30049, 
        n30050, n30051, n30052, n30053, n30054, n30055, n30056, 
        n30057, n30058, n30059, n30060, n30061, n30062, n30063, 
        n30064, n30065, n30066, n30067, n30068, n30069, n30070, 
        n30071, n30072, n30073, n30074, n30075, n30076, n30077, 
        n30078, n30079, n30080, n30081, n30082, n30083, n30084, 
        n30085, n30086, n30087, n30088, n30089, n30090;
    
    FD1P3AX shift_reg_i__i1 (.D(dout_i_23__N_5395[24]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i1.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i1 (.D(\dout_r_23__N_5203[0] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[24]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i1.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i1 (.D(dout_r_23__N_5203[24]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i1.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i1 (.D(\dout_i_23__N_5395[0] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[24]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i1.GSR = "ENABLED";
    FD1P3AX valid_26 (.D(VCC_net), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam valid_26.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i2 (.D(dout_i_23__N_5395[25]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i3 (.D(dout_i_23__N_5395[26]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i4 (.D(dout_i_23__N_5395[27]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i5 (.D(dout_i_23__N_5395[28]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i6 (.D(dout_i_23__N_5395[29]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i7 (.D(dout_i_23__N_5395[30]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i8 (.D(dout_i_23__N_5395[31]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i9 (.D(dout_i_23__N_5395[32]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i10 (.D(dout_i_23__N_5395[33]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i11 (.D(dout_i_23__N_5395[34]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i12 (.D(dout_i_23__N_5395[35]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i13 (.D(dout_i_23__N_5395[36]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i14 (.D(dout_i_23__N_5395[37]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i15 (.D(dout_i_23__N_5395[38]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i16 (.D(dout_i_23__N_5395[39]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i17 (.D(dout_i_23__N_5395[40]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i18 (.D(dout_i_23__N_5395[41]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i19 (.D(dout_i_23__N_5395[42]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i20 (.D(dout_i_23__N_5395[43]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i21 (.D(dout_i_23__N_5395[44]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i22 (.D(dout_i_23__N_5395[45]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i23 (.D(dout_i_23__N_5395[46]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i24 (.D(dout_i_23__N_5395[47]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i24.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i25 (.D(dout_i_23__N_5395[48]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i25.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i26 (.D(dout_i_23__N_5395[49]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i26.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i27 (.D(dout_i_23__N_5395[50]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i27.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i28 (.D(dout_i_23__N_5395[51]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i28.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i29 (.D(dout_i_23__N_5395[52]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i29.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i30 (.D(dout_i_23__N_5395[53]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[77])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i30.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i31 (.D(dout_i_23__N_5395[54]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[78])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i31.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i32 (.D(dout_i_23__N_5395[55]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[79])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i32.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i33 (.D(dout_i_23__N_5395[56]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i33.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i34 (.D(dout_i_23__N_5395[57]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i34.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i35 (.D(dout_i_23__N_5395[58]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i35.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i36 (.D(dout_i_23__N_5395[59]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i36.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i37 (.D(dout_i_23__N_5395[60]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i37.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i38 (.D(dout_i_23__N_5395[61]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[85])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i38.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i39 (.D(dout_i_23__N_5395[62]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[86])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i39.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i40 (.D(dout_i_23__N_5395[63]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[87])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i40.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i41 (.D(dout_i_23__N_5395[64]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i41.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i42 (.D(dout_i_23__N_5395[65]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i42.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i43 (.D(dout_i_23__N_5395[66]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i43.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i44 (.D(dout_i_23__N_5395[67]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i44.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i45 (.D(dout_i_23__N_5395[68]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i45.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i46 (.D(dout_i_23__N_5395[69]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[93])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i46.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i47 (.D(dout_i_23__N_5395[70]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[94])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i47.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i48 (.D(dout_i_23__N_5395[71]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[95])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i48.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i2 (.D(\dout_r_23__N_5203[1] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i3 (.D(\dout_r_23__N_5203[2] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[26]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i4 (.D(\dout_r_23__N_5203[3] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i5 (.D(\dout_r_23__N_5203[4] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[28]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i6 (.D(\dout_r_23__N_5203[5] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i7 (.D(\dout_r_23__N_5203[6] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[30]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i8 (.D(\dout_r_23__N_5203[7] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i9 (.D(\dout_r_23__N_5203[8] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[32]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i10 (.D(\dout_r_23__N_5203[9] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[33]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i11 (.D(\dout_r_23__N_5203[10] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[34]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i12 (.D(\dout_r_23__N_5203[11] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[35]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i13 (.D(\dout_r_23__N_5203[12] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[36]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i14 (.D(\dout_r_23__N_5203[13] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[37]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i15 (.D(\dout_r_23__N_5203[14] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[38]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i16 (.D(\dout_r_23__N_5203[15] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[39]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i17 (.D(\dout_r_23__N_5203[16] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[40]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i18 (.D(\dout_r_23__N_5203[17] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[41]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i19 (.D(\dout_r_23__N_5203[18] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[42]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i20 (.D(\dout_r_23__N_5203[19] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[43]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i21 (.D(\dout_r_23__N_5203[20] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[44]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i22 (.D(\dout_r_23__N_5203[21] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[45]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i23 (.D(\dout_r_23__N_5203[22] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[46]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res3__i24 (.D(\dout_r_23__N_5203[23] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[47]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r_res3__i24.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i2 (.D(dout_r_23__N_5203[25]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i3 (.D(dout_r_23__N_5203[26]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i4 (.D(dout_r_23__N_5203[27]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i5 (.D(dout_r_23__N_5203[28]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i6 (.D(dout_r_23__N_5203[29]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i7 (.D(dout_r_23__N_5203[30]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i8 (.D(dout_r_23__N_5203[31]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i9 (.D(dout_r_23__N_5203[32]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i10 (.D(dout_r_23__N_5203[33]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i11 (.D(dout_r_23__N_5203[34]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i12 (.D(dout_r_23__N_5203[35]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i13 (.D(dout_r_23__N_5203[36]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i14 (.D(dout_r_23__N_5203[37]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i15 (.D(dout_r_23__N_5203[38]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i16 (.D(dout_r_23__N_5203[39]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i17 (.D(dout_r_23__N_5203[40]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i18 (.D(dout_r_23__N_5203[41]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i19 (.D(dout_r_23__N_5203[42]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i20 (.D(dout_r_23__N_5203[43]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i21 (.D(dout_r_23__N_5203[44]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i22 (.D(dout_r_23__N_5203[45]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i23 (.D(dout_r_23__N_5203[46]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i24 (.D(dout_r_23__N_5203[47]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i24.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i25 (.D(dout_r_23__N_5203[48]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i25.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i26 (.D(dout_r_23__N_5203[49]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i26.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i27 (.D(dout_r_23__N_5203[50]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i27.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i28 (.D(dout_r_23__N_5203[51]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i28.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i29 (.D(dout_r_23__N_5203[52]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i29.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i30 (.D(dout_r_23__N_5203[53]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[77])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i30.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i31 (.D(dout_r_23__N_5203[54]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[78])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i31.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i32 (.D(dout_r_23__N_5203[55]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[79])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i32.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i33 (.D(dout_r_23__N_5203[56]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i33.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i34 (.D(dout_r_23__N_5203[57]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i34.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i35 (.D(dout_r_23__N_5203[58]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i35.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i36 (.D(dout_r_23__N_5203[59]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i36.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i37 (.D(dout_r_23__N_5203[60]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i37.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i38 (.D(dout_r_23__N_5203[61]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[85])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i38.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i39 (.D(dout_r_23__N_5203[62]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[86])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i39.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i40 (.D(dout_r_23__N_5203[63]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[87])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i40.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i41 (.D(dout_r_23__N_5203[64]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i41.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i42 (.D(dout_r_23__N_5203[65]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i42.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i43 (.D(dout_r_23__N_5203[66]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i43.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i44 (.D(dout_r_23__N_5203[67]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i44.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i45 (.D(dout_r_23__N_5203[68]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i45.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i46 (.D(dout_r_23__N_5203[69]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[93])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i46.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i47 (.D(dout_r_23__N_5203[70]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[94])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i47.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i48 (.D(dout_r_23__N_5203[71]), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_r_23__N_5203[95])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i48.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i2 (.D(\dout_i_23__N_5395[1] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i3 (.D(\dout_i_23__N_5395[2] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[26]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i4 (.D(\dout_i_23__N_5395[3] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i5 (.D(\dout_i_23__N_5395[4] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[28]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i6 (.D(\dout_i_23__N_5395[5] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i7 (.D(\dout_i_23__N_5395[6] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[30]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i8 (.D(\dout_i_23__N_5395[7] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i9 (.D(\dout_i_23__N_5395[8] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[32]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i10 (.D(\dout_i_23__N_5395[9] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[33]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i11 (.D(\dout_i_23__N_5395[10] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[34]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i12 (.D(\dout_i_23__N_5395[11] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[35]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i13 (.D(\dout_i_23__N_5395[12] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[36]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i14 (.D(\dout_i_23__N_5395[13] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[37]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i15 (.D(\dout_i_23__N_5395[14] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[38]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i16 (.D(\dout_i_23__N_5395[15] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[39]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i17 (.D(\dout_i_23__N_5395[16] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[40]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i18 (.D(\dout_i_23__N_5395[17] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[41]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i19 (.D(\dout_i_23__N_5395[18] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[42]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i20 (.D(\dout_i_23__N_5395[19] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[43]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i21 (.D(\dout_i_23__N_5395[20] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[44]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i22 (.D(\dout_i_23__N_5395[21] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[45]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i23 (.D(\dout_i_23__N_5395[22] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[46]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res2__i24 (.D(\dout_i_23__N_5395[23] ), .SP(clk_c_enable_1373), 
            .CK(clk_c), .Q(dout_i_23__N_5395[47]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i_res2__i24.GSR = "ENABLED";
    LUT4 i12333_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[95]), 
         .D(shift_4_dout_r[23]), .Z(n30043)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12333_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12334_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[94]), 
         .D(shift_4_dout_r[22]), .Z(n30044)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12334_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12335_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[93]), 
         .D(shift_4_dout_r[21]), .Z(n30045)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12335_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12336_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[92]), 
         .D(shift_4_dout_r[20]), .Z(n30046)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12336_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12337_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[91]), 
         .D(shift_4_dout_r[19]), .Z(n30047)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12337_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12338_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[90]), 
         .D(shift_4_dout_r[18]), .Z(n30048)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12338_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12339_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[89]), 
         .D(shift_4_dout_r[17]), .Z(n30049)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12339_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12340_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[88]), 
         .D(shift_4_dout_r[16]), .Z(n30050)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12340_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12341_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[87]), 
         .D(shift_4_dout_r[15]), .Z(n30051)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12341_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12342_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[86]), 
         .D(shift_4_dout_r[14]), .Z(n30052)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12342_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12343_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[85]), 
         .D(shift_4_dout_r[13]), .Z(n30053)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12343_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12344_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[84]), 
         .D(shift_4_dout_r[12]), .Z(n30054)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12344_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12345_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[83]), 
         .D(shift_4_dout_r[11]), .Z(n30055)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12345_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12346_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[82]), 
         .D(shift_4_dout_r[10]), .Z(n30056)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12346_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12347_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[81]), 
         .D(shift_4_dout_r[9]), .Z(n30057)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12347_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12348_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[80]), 
         .D(shift_4_dout_r[8]), .Z(n30058)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12348_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12349_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[79]), 
         .D(shift_4_dout_r[7]), .Z(n30059)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12349_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12350_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[78]), 
         .D(shift_4_dout_r[6]), .Z(n30060)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12350_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12351_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[77]), 
         .D(shift_4_dout_r[5]), .Z(n30061)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12351_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12352_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[76]), 
         .D(shift_4_dout_r[4]), .Z(n30062)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12352_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12353_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[75]), 
         .D(shift_4_dout_r[3]), .Z(n30063)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12353_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12354_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[74]), 
         .D(shift_4_dout_r[2]), .Z(n30064)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12354_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12355_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[73]), 
         .D(shift_4_dout_r[1]), .Z(n30065)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12355_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12356_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_r_23__N_5203[72]), 
         .D(shift_4_dout_r[0]), .Z(n30066)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12356_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12357_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[95]), 
         .D(shift_4_dout_i[23]), .Z(n30067)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12357_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12358_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[94]), 
         .D(shift_4_dout_i[22]), .Z(n30068)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12358_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12359_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[93]), 
         .D(shift_4_dout_i[21]), .Z(n30069)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12359_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12360_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[92]), 
         .D(shift_4_dout_i[20]), .Z(n30070)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12360_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12361_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[91]), 
         .D(shift_4_dout_i[19]), .Z(n30071)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12361_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12362_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[90]), 
         .D(shift_4_dout_i[18]), .Z(n30072)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12362_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12363_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[89]), 
         .D(shift_4_dout_i[17]), .Z(n30073)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12363_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12364_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[88]), 
         .D(shift_4_dout_i[16]), .Z(n30074)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12364_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12365_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[87]), 
         .D(shift_4_dout_i[15]), .Z(n30075)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12365_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12366_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[86]), 
         .D(shift_4_dout_i[14]), .Z(n30076)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12366_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12367_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[85]), 
         .D(shift_4_dout_i[13]), .Z(n30077)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12367_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12368_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[84]), 
         .D(shift_4_dout_i[12]), .Z(n30078)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12368_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12369_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[83]), 
         .D(shift_4_dout_i[11]), .Z(n30079)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12369_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12370_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[82]), 
         .D(shift_4_dout_i[10]), .Z(n30080)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12370_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12371_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[81]), 
         .D(shift_4_dout_i[9]), .Z(n30081)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12371_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12372_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[80]), 
         .D(shift_4_dout_i[8]), .Z(n30082)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12372_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12373_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[79]), 
         .D(shift_4_dout_i[7]), .Z(n30083)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12373_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12374_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[78]), 
         .D(shift_4_dout_i[6]), .Z(n30084)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12374_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12375_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[77]), 
         .D(shift_4_dout_i[5]), .Z(n30085)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12375_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12376_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[76]), 
         .D(shift_4_dout_i[4]), .Z(n30086)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12376_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12377_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[75]), 
         .D(shift_4_dout_i[3]), .Z(n30087)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12377_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12378_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[74]), 
         .D(shift_4_dout_i[2]), .Z(n30088)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12378_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12379_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[73]), 
         .D(shift_4_dout_i[1]), .Z(n30089)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12379_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12380_3_lut_4_lut (.A(valid), .B(n34842), .C(dout_i_23__N_5395[72]), 
         .D(shift_4_dout_i[0]), .Z(n30090)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(41[14] 46[8])
    defparam i12380_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX shift_reg_i__i49 (.D(n30090), .CK(clk_c), .Q(shift_4_dout_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i49.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i50 (.D(n30089), .CK(clk_c), .Q(shift_4_dout_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i50.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i51 (.D(n30088), .CK(clk_c), .Q(shift_4_dout_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i51.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i52 (.D(n30087), .CK(clk_c), .Q(shift_4_dout_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i52.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i53 (.D(n30086), .CK(clk_c), .Q(shift_4_dout_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i53.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i54 (.D(n30085), .CK(clk_c), .Q(shift_4_dout_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i54.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i55 (.D(n30084), .CK(clk_c), .Q(shift_4_dout_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i55.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i56 (.D(n30083), .CK(clk_c), .Q(shift_4_dout_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i56.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i57 (.D(n30082), .CK(clk_c), .Q(shift_4_dout_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i57.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i58 (.D(n30081), .CK(clk_c), .Q(shift_4_dout_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i58.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i59 (.D(n30080), .CK(clk_c), .Q(shift_4_dout_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i59.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i60 (.D(n30079), .CK(clk_c), .Q(shift_4_dout_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i60.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i61 (.D(n30078), .CK(clk_c), .Q(shift_4_dout_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i61.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i62 (.D(n30077), .CK(clk_c), .Q(shift_4_dout_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i62.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i63 (.D(n30076), .CK(clk_c), .Q(shift_4_dout_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i63.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i64 (.D(n30075), .CK(clk_c), .Q(shift_4_dout_i[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i64.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i65 (.D(n30074), .CK(clk_c), .Q(shift_4_dout_i[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i65.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i66 (.D(n30073), .CK(clk_c), .Q(shift_4_dout_i[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i66.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i67 (.D(n30072), .CK(clk_c), .Q(shift_4_dout_i[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i67.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i68 (.D(n30071), .CK(clk_c), .Q(shift_4_dout_i[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i68.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i69 (.D(n30070), .CK(clk_c), .Q(shift_4_dout_i[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i69.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i70 (.D(n30069), .CK(clk_c), .Q(shift_4_dout_i[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i70.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i71 (.D(n30068), .CK(clk_c), .Q(shift_4_dout_i[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i71.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i72 (.D(n30067), .CK(clk_c), .Q(shift_4_dout_i[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_i__i72.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i49 (.D(n30066), .CK(clk_c), .Q(shift_4_dout_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i49.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i50 (.D(n30065), .CK(clk_c), .Q(shift_4_dout_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i50.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i51 (.D(n30064), .CK(clk_c), .Q(shift_4_dout_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i51.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i52 (.D(n30063), .CK(clk_c), .Q(shift_4_dout_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i52.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i53 (.D(n30062), .CK(clk_c), .Q(shift_4_dout_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i53.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i54 (.D(n30061), .CK(clk_c), .Q(shift_4_dout_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i54.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i55 (.D(n30060), .CK(clk_c), .Q(shift_4_dout_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i55.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i56 (.D(n30059), .CK(clk_c), .Q(shift_4_dout_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i56.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i57 (.D(n30058), .CK(clk_c), .Q(shift_4_dout_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i57.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i58 (.D(n30057), .CK(clk_c), .Q(shift_4_dout_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i58.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i59 (.D(n30056), .CK(clk_c), .Q(shift_4_dout_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i59.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i60 (.D(n30055), .CK(clk_c), .Q(shift_4_dout_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i60.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i61 (.D(n30054), .CK(clk_c), .Q(shift_4_dout_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i61.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i62 (.D(n30053), .CK(clk_c), .Q(shift_4_dout_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i62.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i63 (.D(n30052), .CK(clk_c), .Q(shift_4_dout_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i63.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i64 (.D(n30051), .CK(clk_c), .Q(shift_4_dout_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i64.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i65 (.D(n30050), .CK(clk_c), .Q(shift_4_dout_r[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i65.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i66 (.D(n30049), .CK(clk_c), .Q(shift_4_dout_r[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i66.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i67 (.D(n30048), .CK(clk_c), .Q(shift_4_dout_r[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i67.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i68 (.D(n30047), .CK(clk_c), .Q(shift_4_dout_r[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i68.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i69 (.D(n30046), .CK(clk_c), .Q(shift_4_dout_r[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i69.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i70 (.D(n30045), .CK(clk_c), .Q(shift_4_dout_r[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i70.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i71 (.D(n30044), .CK(clk_c), .Q(shift_4_dout_r[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i71.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i72 (.D(n30043), .CK(clk_c), .Q(shift_4_dout_r[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=164, LSE_RLINE=171 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_4.v(36[5] 46[8])
    defparam shift_reg_r__i72.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module ROM_8
//

module ROM_8 (n29816, n29815, n34532, \rom8_state[0] , s_count, clk_c, 
            clk_c_enable_2285, clk_c_enable_2310, n34726, n34788, \rom8_w_i[12] , 
            n29782, n5, n29824, n29823, n29822, n34842, n30191, 
            GND_net, VCC_net, n34762, n34761, n34760, \rom8_w_i[1] , 
            n34785, n34734, \rom8_w_i[4] , \rom8_w_i[3] , n34787, 
            \rom8_w_i[0] , \rom8_w_i[6] , n34742, \rom8_w_i[2] , n6, 
            n34778, \rom8_w_r[0] , \rom8_w_r[7] , n34752, n34753, 
            \rom8_w_r[4] , \rom8_w_r[3] , \rom8_w_r[6] , n34779, \rom8_w_r[1] , 
            n34754, \rom8_w_r[8] , \rom8_w_r[5] , \rom8_w_r[10] , n34794, 
            n34755, n34756, clk_c_enable_2305, n30040) /* synthesis syn_module_defined=1 */ ;
    output n29816;
    output n29815;
    output n34532;
    output \rom8_state[0] ;
    output [3:0]s_count;
    input clk_c;
    output clk_c_enable_2285;
    input clk_c_enable_2310;
    output n34726;
    output n34788;
    output \rom8_w_i[12] ;
    output n29782;
    output n5;
    output n29824;
    output n29823;
    output n29822;
    output n34842;
    output n30191;
    input GND_net;
    input VCC_net;
    output n34762;
    output n34761;
    output n34760;
    output \rom8_w_i[1] ;
    output n34785;
    output n34734;
    output \rom8_w_i[4] ;
    output \rom8_w_i[3] ;
    output n34787;
    output \rom8_w_i[0] ;
    output \rom8_w_i[6] ;
    output n34742;
    output \rom8_w_i[2] ;
    output n6;
    output n34778;
    output \rom8_w_r[0] ;
    output \rom8_w_r[7] ;
    output n34752;
    output n34753;
    output \rom8_w_r[4] ;
    output \rom8_w_r[3] ;
    output \rom8_w_r[6] ;
    output n34779;
    output \rom8_w_r[1] ;
    output n34754;
    output \rom8_w_r[8] ;
    output \rom8_w_r[5] ;
    output \rom8_w_r[10] ;
    output n34794;
    output n34755;
    output n34756;
    output clk_c_enable_2305;
    input n30040;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire n34773;
    wire [5:0]n51;
    wire [5:0]n29;
    wire [3:0]n21;
    
    wire n32401;
    wire [5:0]count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(11[11:16])
    
    wire n32400, n32399;
    
    LUT4 i12107_3_lut (.A(n29816), .B(n29815), .C(n34532), .Z(\rom8_state[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(14[1] 73[4])
    defparam i12107_3_lut.init = 16'hcaca;
    FD1P3AX s_count_691__i0 (.D(n34773), .SP(clk_c_enable_2285), .CK(clk_c), 
            .Q(s_count[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam s_count_691__i0.GSR = "ENABLED";
    FD1P3AX count_692__i0 (.D(n29[0]), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(n51[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692__i0.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(s_count[0]), .B(n34726), .C(s_count[1]), .D(n34788), 
         .Z(\rom8_w_i[12] )) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i2_4_lut.init = 16'h3733;
    LUT4 i1_2_lut (.A(s_count[0]), .B(s_count[1]), .Z(n29782)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(60[5:10])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_adj_198 (.A(s_count[3]), .B(s_count[1]), .Z(n5)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_198.init = 16'h2222;
    LUT4 i2352_2_lut_rep_446 (.A(n29824), .B(n29823), .C(n29822), .D(\rom8_state[0] ), 
         .Z(n34842)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(14[1] 73[4])
    defparam i2352_2_lut_rep_446.init = 16'h35ca;
    LUT4 i13999_2_lut (.A(s_count[1]), .B(s_count[0]), .Z(n21[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam i13999_2_lut.init = 16'h6666;
    LUT4 s_count_3__bdd_4_lut (.A(s_count[3]), .B(s_count[2]), .C(s_count[1]), 
         .D(s_count[0]), .Z(n30191)) /* synthesis lut_function=((B (C+!(D))+!B !(C (D)))+!A) */ ;
    defparam s_count_3__bdd_4_lut.init = 16'hd7ff;
    CCU2C count_692_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32401), .S0(n29[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692_add_4_7.INIT0 = 16'haaa0;
    defparam count_692_add_4_7.INIT1 = 16'h0000;
    defparam count_692_add_4_7.INJECT1_0 = "NO";
    defparam count_692_add_4_7.INJECT1_1 = "NO";
    CCU2C count_692_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32400), .COUT(n32401), .S0(n29[3]), .S1(n29[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692_add_4_5.INIT0 = 16'haaa0;
    defparam count_692_add_4_5.INIT1 = 16'haaa0;
    defparam count_692_add_4_5.INJECT1_0 = "NO";
    defparam count_692_add_4_5.INJECT1_1 = "NO";
    CCU2C count_692_add_4_3 (.A0(n51[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n51[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32399), .COUT(n32400), .S0(n29[1]), .S1(n29[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692_add_4_3.INIT0 = 16'haaa0;
    defparam count_692_add_4_3.INIT1 = 16'haaa0;
    defparam count_692_add_4_3.INJECT1_0 = "NO";
    defparam count_692_add_4_3.INJECT1_1 = "NO";
    CCU2C count_692_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n51[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32399), .S1(n29[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692_add_4_1.INIT0 = 16'h0000;
    defparam count_692_add_4_1.INIT1 = 16'h555f;
    defparam count_692_add_4_1.INJECT1_0 = "NO";
    defparam count_692_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_400_4_lut_2_lut_4_lut (.A(s_count[3]), .B(s_count[0]), 
         .C(s_count[1]), .Z(n34762)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i1_3_lut_rep_400_4_lut_2_lut_4_lut.init = 16'hdfdf;
    LUT4 i12539_2_lut_rep_364_3_lut_4_lut (.A(n34761), .B(n34760), .C(n30191), 
         .D(n34762), .Z(n34726)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i12539_2_lut_rep_364_3_lut_4_lut.init = 16'h2000;
    LUT4 i12540_1_lut_2_lut_3_lut_4_lut (.A(n34761), .B(n34760), .C(n30191), 
         .D(n34762), .Z(\rom8_w_i[1] )) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i12540_1_lut_2_lut_3_lut_4_lut.init = 16'hdfff;
    LUT4 i16395_3_lut_3_lut (.A(clk_c_enable_2285), .B(s_count[3]), .C(n29816), 
         .Z(n29816)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i16395_3_lut_3_lut.init = 16'h2020;
    LUT4 i16399_3_lut_3_lut (.A(clk_c_enable_2285), .B(s_count[3]), .C(n29815), 
         .Z(n29815)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam i16399_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i16379_3_lut_3_lut (.A(s_count[3]), .B(clk_c_enable_2285), .C(n29824), 
         .Z(n29824)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(27[10] 34[8])
    defparam i16379_3_lut_3_lut.init = 16'h8080;
    LUT4 i16383_4_lut_2_lut_3_lut (.A(s_count[3]), .B(clk_c_enable_2285), 
         .C(n29823), .Z(n29823)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(27[10] 34[8])
    defparam i16383_4_lut_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i12483_2_lut_rep_372_3_lut_4_lut (.A(n34788), .B(n34785), .C(n34762), 
         .D(n34761), .Z(n34734)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i12483_2_lut_rep_372_3_lut_4_lut.init = 16'h7000;
    LUT4 i16330_2_lut_3_lut_4_lut (.A(n34788), .B(n34785), .C(n30191), 
         .D(n34761), .Z(\rom8_w_i[4] )) /* synthesis lut_function=(A (B+!(C (D)))+!A !(C (D))) */ ;
    defparam i16330_2_lut_3_lut_4_lut.init = 16'h8fff;
    LUT4 i12484_1_lut_2_lut_3_lut_4_lut (.A(n34788), .B(n34785), .C(n34762), 
         .D(n34761), .Z(\rom8_w_i[3] )) /* synthesis lut_function=(A (B+!(C (D)))+!A !(C (D))) */ ;
    defparam i12484_1_lut_2_lut_3_lut_4_lut.init = 16'h8fff;
    LUT4 i16327_2_lut_4_lut (.A(n29782), .B(n34787), .C(n34788), .D(n30191), 
         .Z(\rom8_w_i[0] )) /* synthesis lut_function=(!(A (D)+!A !((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(60[5:10])
    defparam i16327_2_lut_4_lut.init = 16'h51ff;
    LUT4 i12480_1_lut_3_lut_4_lut_2_lut_4_lut (.A(s_count[3]), .B(s_count[0]), 
         .C(s_count[1]), .Z(\rom8_w_i[6] )) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i12480_1_lut_3_lut_4_lut_2_lut_4_lut.init = 16'h2020;
    LUT4 i12477_2_lut_rep_380_3_lut_4_lut_4_lut (.A(s_count[2]), .B(s_count[3]), 
         .C(s_count[1]), .D(s_count[0]), .Z(n34742)) /* synthesis lut_function=(!(A (B (C (D)))+!A !((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(56[5:10])
    defparam i12477_2_lut_rep_380_3_lut_4_lut_4_lut.init = 16'h7bff;
    LUT4 i12478_1_lut_2_lut_3_lut_4_lut_4_lut (.A(s_count[2]), .B(s_count[3]), 
         .C(s_count[1]), .D(s_count[0]), .Z(\rom8_w_i[2] )) /* synthesis lut_function=(A (B (C (D)))+!A !((C+!(D))+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(56[5:10])
    defparam i12478_1_lut_2_lut_3_lut_4_lut_4_lut.init = 16'h8400;
    LUT4 i2_1_lut_rep_411 (.A(s_count[0]), .Z(n34773)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut_rep_411.init = 16'h5555;
    LUT4 i2_2_lut_2_lut (.A(s_count[0]), .B(s_count[2]), .Z(n6)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i2_2_lut_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_rep_412 (.A(count[4]), .B(count[5]), .C(count[3]), .Z(clk_c_enable_2285)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_412.init = 16'hfefe;
    LUT4 i16367_3_lut_2_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .D(s_count[3]), .Z(n34532)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i16367_3_lut_2_lut_4_lut.init = 16'h00fe;
    LUT4 i16359_3_lut_2_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .D(s_count[3]), .Z(n29822)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i16359_3_lut_2_lut_4_lut.init = 16'hfe00;
    LUT4 i10884_3_lut_rep_416 (.A(s_count[1]), .B(s_count[2]), .C(s_count[0]), 
         .Z(n34778)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C))) */ ;
    defparam i10884_3_lut_rep_416.init = 16'h9a9a;
    LUT4 i12502_2_lut_4_lut (.A(s_count[1]), .B(s_count[2]), .C(s_count[0]), 
         .D(s_count[3]), .Z(\rom8_w_r[0] )) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B+!(C (D)))) */ ;
    defparam i12502_2_lut_4_lut.init = 16'h9a00;
    LUT4 i12450_2_lut_4_lut_4_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[3]), 
         .D(s_count[0]), .Z(\rom8_w_r[7] )) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B ((D)+!C)+!B !(C (D))))) */ ;
    defparam i12450_2_lut_4_lut_4_lut.init = 16'h3040;
    LUT4 i10878_3_lut_rep_390_3_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), 
         .Z(n34752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C)+!B !(C))) */ ;
    defparam i10878_3_lut_rep_390_3_lut.init = 16'hcbcb;
    LUT4 i2377_3_lut_rep_391_3_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), 
         .Z(n34753)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;
    defparam i2377_3_lut_rep_391_3_lut.init = 16'h5b5b;
    LUT4 i12507_2_lut_4_lut_4_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[3]), 
         .D(s_count[0]), .Z(\rom8_w_r[4] )) /* synthesis lut_function=(A (C (D))+!A !(((D)+!C)+!B)) */ ;
    defparam i12507_2_lut_4_lut_4_lut.init = 16'ha040;
    LUT4 i12459_4_lut_4_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), 
         .D(s_count[3]), .Z(\rom8_w_r[3] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+!(C (D))))) */ ;
    defparam i12459_4_lut_4_lut.init = 16'h3800;
    LUT4 i12476_4_lut_4_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), 
         .D(s_count[3]), .Z(\rom8_w_r[6] )) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(C (D)))) */ ;
    defparam i12476_4_lut_4_lut.init = 16'h5800;
    LUT4 i10882_4_lut_3_lut_rep_417 (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), 
         .Z(n34779)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;
    defparam i10882_4_lut_3_lut_rep_417.init = 16'he8e8;
    LUT4 i12501_2_lut_4_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), 
         .D(s_count[3]), .Z(\rom8_w_r[1] )) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (C (D)))) */ ;
    defparam i12501_2_lut_4_lut.init = 16'he800;
    LUT4 i13337_3_lut_rep_392_4_lut (.A(s_count[0]), .B(s_count[1]), .C(s_count[2]), 
         .D(s_count[3]), .Z(n34754)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C (D))))) */ ;
    defparam i13337_3_lut_rep_392_4_lut.init = 16'h1e00;
    LUT4 i13338_1_lut_3_lut_4_lut (.A(s_count[0]), .B(s_count[1]), .C(s_count[2]), 
         .D(s_count[3]), .Z(\rom8_w_r[8] )) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam i13338_1_lut_3_lut_4_lut.init = 16'he1ff;
    LUT4 i1_2_lut_3_lut_4_lut (.A(s_count[0]), .B(s_count[1]), .C(s_count[2]), 
         .D(s_count[3]), .Z(\rom8_w_r[5] )) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_199 (.A(s_count[0]), .B(s_count[1]), .C(s_count[2]), 
         .D(s_count[3]), .Z(\rom8_w_r[10] )) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_199.init = 16'he000;
    LUT4 i14002_2_lut_rep_423 (.A(s_count[1]), .B(s_count[0]), .Z(n34785)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam i14002_2_lut_rep_423.init = 16'h8888;
    LUT4 i14006_2_lut_3_lut (.A(s_count[1]), .B(s_count[0]), .C(s_count[2]), 
         .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam i14006_2_lut_3_lut.init = 16'h7878;
    LUT4 s_count_3__I_0_65_i6_2_lut_rep_425 (.A(s_count[2]), .B(s_count[3]), 
         .Z(n34787)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(44[5:10])
    defparam s_count_3__I_0_65_i6_2_lut_rep_425.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_399_3_lut_4_lut (.A(s_count[2]), .B(s_count[3]), .C(s_count[0]), 
         .D(s_count[1]), .Z(n34761)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(44[5:10])
    defparam i1_2_lut_rep_399_3_lut_4_lut.init = 16'hffbf;
    LUT4 i12547_2_lut_rep_426 (.A(s_count[2]), .B(s_count[3]), .Z(n34788)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12547_2_lut_rep_426.init = 16'h8888;
    LUT4 i13306_2_lut_rep_398_3_lut_4_lut (.A(s_count[2]), .B(s_count[3]), 
         .C(s_count[0]), .D(s_count[1]), .Z(n34760)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13306_2_lut_rep_398_3_lut_4_lut.init = 16'h8000;
    LUT4 i12115_3_lut_rep_432 (.A(n29824), .B(n29823), .C(n29822), .Z(n34794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(14[1] 73[4])
    defparam i12115_3_lut_rep_432.init = 16'hcaca;
    LUT4 equal_370_i3_2_lut_rep_393_4_lut (.A(n29824), .B(n29823), .C(n29822), 
         .D(\rom8_state[0] ), .Z(n34755)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(14[1] 73[4])
    defparam equal_370_i3_2_lut_rep_393_4_lut.init = 16'hcaff;
    LUT4 i166_2_lut_rep_394_4_lut (.A(n29824), .B(n29823), .C(n29822), 
         .D(\rom8_state[0] ), .Z(n34756)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(14[1] 73[4])
    defparam i166_2_lut_rep_394_4_lut.init = 16'h00ca;
    LUT4 i2352_2_lut_rep_403_4_lut (.A(n29824), .B(n29823), .C(n29822), 
         .D(\rom8_state[0] ), .Z(clk_c_enable_2305)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(14[1] 73[4])
    defparam i2352_2_lut_rep_403_4_lut.init = 16'h35ca;
    FD1S3AX s_count_691__i3 (.D(n30040), .CK(clk_c), .Q(s_count[3]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam s_count_691__i3.GSR = "ENABLED";
    FD1P3AX s_count_691__i1 (.D(n21[1]), .SP(clk_c_enable_2285), .CK(clk_c), 
            .Q(s_count[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam s_count_691__i1.GSR = "ENABLED";
    FD1P3AX s_count_691__i2 (.D(n21[2]), .SP(clk_c_enable_2285), .CK(clk_c), 
            .Q(s_count[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(33[24:35])
    defparam s_count_691__i2.GSR = "ENABLED";
    FD1P3AX count_692__i1 (.D(n29[1]), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(n51[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692__i1.GSR = "ENABLED";
    FD1P3AX count_692__i2 (.D(n29[2]), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(n51[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692__i2.GSR = "ENABLED";
    FD1P3AX count_692__i3 (.D(n29[3]), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692__i3.GSR = "ENABLED";
    FD1P3AX count_692__i4 (.D(n29[4]), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692__i4.GSR = "ENABLED";
    FD1P3AX count_692__i5 (.D(n29[5]), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_8.v(17[22:31])
    defparam count_692__i5.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module radix2_U3
//

module radix2_U3 (op_r_23__N_1106, \count[5] , \count[4] , \op_r_23__N_1082[8] , 
            \radix_no1_op_r[0] , \op_r_23__N_1082[9] , \radix_no1_op_r[1] , 
            GND_net, \op_r_23__N_1268[0] , \op_r_23__N_1268[1] , \op_r_23__N_1268[2] , 
            \op_r_23__N_1268[3] , \op_r_23__N_1268[4] , \op_r_23__N_1268[5] , 
            \op_r_23__N_1268[6] , \op_r_23__N_1268[7] , \op_r_23__N_1268[8] , 
            \op_r_23__N_1268[9] , \op_r_23__N_1268[10] , \op_r_23__N_1268[11] , 
            \op_r_23__N_1268[12] , \op_r_23__N_1268[13] , \op_r_23__N_1268[14] , 
            \op_r_23__N_1268[15] , \op_r_23__N_1268[16] , \op_r_23__N_1268[17] , 
            VCC_net, \op_r_23__N_1082[10] , \radix_no1_op_r[2] , \op_r_23__N_1082[11] , 
            \radix_no1_op_r[3] , \op_r_23__N_1082[12] , \radix_no1_op_r[4] , 
            \op_i_23__N_1310[0] , \op_i_23__N_1310[1] , \op_i_23__N_1310[2] , 
            \op_i_23__N_1310[3] , \op_i_23__N_1310[4] , \op_i_23__N_1310[5] , 
            n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, 
            n79, n78, n77, n76, n75, n74, n73, n72, n71, n70, 
            n69, n68, n67, n66, n65, \rom16_w_i[8] , n9983, n9984, 
            n9985, n9986, n9987, n9988, \rom16_w_i[0] , \rom16_w_i[1] , 
            \rom16_w_i[2] , \rom16_w_i[3] , \rom16_w_i[4] , \rom16_w_i[5] , 
            \rom16_w_i[6] , \rom16_w_i[7] , \op_r_23__N_1082[13] , \radix_no1_op_r[5] , 
            \op_r_23__N_1226[0] , \op_r_23__N_1226[1] , \op_r_23__N_1226[2] , 
            \op_r_23__N_1226[3] , \op_r_23__N_1226[4] , \op_r_23__N_1226[5] , 
            \op_r_23__N_1226[6] , \op_r_23__N_1226[7] , \op_r_23__N_1226[8] , 
            \op_r_23__N_1226[9] , \op_r_23__N_1226[10] , \op_r_23__N_1226[11] , 
            \op_r_23__N_1226[12] , \op_r_23__N_1226[13] , \op_r_23__N_1226[14] , 
            \op_r_23__N_1226[15] , \op_r_23__N_1226[16] , \op_r_23__N_1226[17] , 
            \op_r_23__N_1226[18] , \op_r_23__N_1226[19] , \op_r_23__N_1226[20] , 
            \op_r_23__N_1226[21] , \op_r_23__N_1226[22] , \op_r_23__N_1226[23] , 
            \op_r_23__N_1226[24] , \op_r_23__N_1226[25] , \op_r_23__N_1226[26] , 
            \op_r_23__N_1226[27] , \op_r_23__N_1226[28] , \op_r_23__N_1226[29] , 
            \op_r_23__N_1226[30] , \op_r_23__N_1226[31] , \op_r_23__N_1082[14] , 
            \radix_no1_op_r[6] , \op_r_23__N_1268[18] , \op_r_23__N_1268[19] , 
            \op_r_23__N_1268[20] , \op_r_23__N_1268[21] , \op_r_23__N_1268[22] , 
            \op_r_23__N_1268[23] , \op_r_23__N_1268[24] , \op_r_23__N_1268[25] , 
            \op_r_23__N_1268[26] , \op_r_23__N_1268[27] , \op_r_23__N_1268[28] , 
            \op_r_23__N_1268[29] , \op_r_23__N_1268[30] , \op_r_23__N_1268[31] , 
            \rom16_w_r[9] , n12332, n12333, n12334, n12335, n12336, 
            n12337, n12338, \rom16_w_r[0] , \rom16_w_r[1] , \rom16_w_r[2] , 
            \rom16_w_r[3] , \rom16_w_r[4] , \rom16_w_r[5] , \rom16_w_r[6] , 
            \rom16_w_r[7] , \rom16_w_r[8] , n12314, n12315, n12316, 
            n12317, n12318, n12319, n12320, n12321, n12322, n12323, 
            n12324, n12325, n12326, n12327, n12328, n12329, n12330, 
            n12331, \op_r_23__N_1082[15] , \radix_no1_op_r[7] , op_i_23__N_1154, 
            \op_i_23__N_1130[8] , \radix_no1_op_i[0] , \op_i_23__N_1130[9] , 
            \radix_no1_op_i[1] , \op_i_23__N_1130[10] , \radix_no1_op_i[2] , 
            \op_i_23__N_1130[11] , \radix_no1_op_i[3] , \op_i_23__N_1130[12] , 
            \radix_no1_op_i[4] , \op_i_23__N_1130[13] , \radix_no1_op_i[5] , 
            \op_i_23__N_1130[14] , \radix_no1_op_i[6] , \op_i_23__N_1130[15] , 
            \radix_no1_op_i[7] , n8593, n8592, n8591, n8590, n8589, 
            n8588, n8587, n8586, n8585, n8584, n8583, n8582, n8581, 
            n8580, n8579, n8578, n8577, n8576, n8575, n8574, n8573, 
            n8572, n8571, n8570, n8569, n8568, n319, n9989, n9990, 
            n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, 
            n9999, n10000, n10001, n10002, n10003, n10004, n10005, 
            n10006, \shift_16_dout_i[8] , \shift_16_dout_i[9] , \shift_16_dout_i[10] , 
            \shift_16_dout_i[11] , \shift_16_dout_i[12] , \shift_16_dout_i[13] , 
            \shift_16_dout_i[14] , \shift_16_dout_i[15] , \shift_16_dout_i[16] , 
            \shift_16_dout_i[17] , n12344, n12345, n12346, n12347, 
            n12348, n12349, n12350, n12351, n12352, n12353, n12368, 
            \shift_16_dout_i[18] , \shift_16_dout_i[19] , \shift_16_dout_i[20] , 
            \shift_16_dout_i[21] , \shift_16_dout_i[22] , \shift_16_dout_i[23] , 
            clk_c_enable_2310, n34755, \shift_8_dout_r[22] , n7539, 
            n34756, \op_r_23__N_1082[30] , n31574, \shift_8_dout_r[23] , 
            n7538, \op_r_23__N_1082[31] , n31572, \shift_8_dout_i[22] , 
            n7486, \op_i_23__N_1130[30] , n31378, \shift_8_dout_i[23] , 
            n7485, \op_i_23__N_1130[31] , n31376, \shift_8_dout_r[20] , 
            n7541, \op_r_23__N_1082[28] , n31578, \shift_8_dout_r[21] , 
            n7540, \op_r_23__N_1082[29] , n31576, \shift_8_dout_i[20] , 
            n7488, \op_i_23__N_1130[28] , n31382, \shift_8_dout_i[21] , 
            n7487, \op_i_23__N_1130[29] , n31380, \shift_8_dout_r[18] , 
            n7543, \op_r_23__N_1082[26] , n31582, \shift_8_dout_r[19] , 
            n7542, \op_r_23__N_1082[27] , n31580, \shift_8_dout_i[18] , 
            n7490, \op_i_23__N_1130[26] , n31386, \shift_8_dout_i[19] , 
            n7489, \op_i_23__N_1130[27] , n31384, \shift_8_dout_r[16] , 
            n7545, \op_r_23__N_1082[24] , n31586, \shift_8_dout_r[17] , 
            n7544, \op_r_23__N_1082[25] , n31584, \shift_8_dout_i[16] , 
            n7492, \op_i_23__N_1130[24] , n31390, \shift_8_dout_i[17] , 
            n7491, \op_i_23__N_1130[25] , n31388, \shift_8_dout_r[14] , 
            n7547, \op_r_23__N_1082[22] , n31590, \shift_8_dout_r[15] , 
            n7546, \op_r_23__N_1082[23] , n31588, \shift_8_dout_i[14] , 
            n7494, \op_i_23__N_1130[22] , n31394, \shift_8_dout_i[15] , 
            n7493, \op_i_23__N_1130[23] , n31392, \shift_8_dout_r[12] , 
            n7549, \op_r_23__N_1082[20] , n31594, \shift_8_dout_r[13] , 
            n7548, \op_r_23__N_1082[21] , n31592, \shift_8_dout_i[12] , 
            n7496, \op_i_23__N_1130[20] , n31398, \shift_8_dout_i[13] , 
            n7495, \op_i_23__N_1130[21] , n31396, \shift_8_dout_r[10] , 
            n7551, \op_r_23__N_1082[18] , n31598, \shift_8_dout_r[11] , 
            n7550, \op_r_23__N_1082[19] , n31596, \shift_8_dout_i[10] , 
            n7498, \op_i_23__N_1130[18] , n31402, \shift_8_dout_i[11] , 
            n7497, \op_i_23__N_1130[19] , n31400, \shift_8_dout_r[8] , 
            n7553, \op_r_23__N_1082[16] , n31602, \shift_8_dout_r[9] , 
            n7552, \op_r_23__N_1082[17] , n31600, \shift_8_dout_i[8] , 
            n7500, \op_i_23__N_1130[16] , n31406, \shift_8_dout_i[9] , 
            n7499, \op_i_23__N_1130[17] , n31404, \din_r_reg[8] , \delay_r_23__N_1178[8] , 
            \dout_r_23__N_2506[8] , \din_r_reg[9] , \delay_r_23__N_1178[9] , 
            \dout_r_23__N_2506[9] , \din_r_reg[10] , \delay_r_23__N_1178[10] , 
            \dout_r_23__N_2506[10] , \din_r_reg[11] , \delay_r_23__N_1178[11] , 
            \dout_r_23__N_2506[11] , \din_r_reg[12] , \delay_r_23__N_1178[12] , 
            \dout_r_23__N_2506[12] , \din_r_reg[13] , \delay_r_23__N_1178[13] , 
            \dout_r_23__N_2506[13] , \din_r_reg[14] , \delay_r_23__N_1178[14] , 
            \dout_r_23__N_2506[14] , \din_r_reg[15] , \delay_r_23__N_1178[15] , 
            \dout_r_23__N_2506[15] , \din_r_reg[16] , \delay_r_23__N_1178[16] , 
            \dout_r_23__N_2506[16] , \din_r_reg[17] , \delay_r_23__N_1178[17] , 
            \dout_r_23__N_2506[17] , \din_r_reg[18] , \delay_r_23__N_1178[18] , 
            \dout_r_23__N_2506[18] , \din_r_reg[23] , \delay_r_23__N_1178[19] , 
            \dout_r_23__N_2506[19] , \delay_r_23__N_1178[20] , \dout_r_23__N_2506[20] , 
            \delay_r_23__N_1178[21] , \dout_r_23__N_2506[21] , \delay_r_23__N_1178[22] , 
            \dout_r_23__N_2506[22] , \delay_r_23__N_1178[23] , \dout_r_23__N_2506[23] , 
            \din_i_reg[8] , \delay_i_23__N_1202[8] , \dout_i_23__N_3274[8] , 
            \din_i_reg[9] , \delay_i_23__N_1202[9] , \dout_i_23__N_3274[9] , 
            \din_i_reg[10] , \delay_i_23__N_1202[10] , \dout_i_23__N_3274[10] , 
            \din_i_reg[11] , \delay_i_23__N_1202[11] , \dout_i_23__N_3274[11] , 
            \din_i_reg[12] , \delay_i_23__N_1202[12] , \dout_i_23__N_3274[12] , 
            \din_i_reg[13] , \delay_i_23__N_1202[13] , \dout_i_23__N_3274[13] , 
            \din_i_reg[14] , \delay_i_23__N_1202[14] , \dout_i_23__N_3274[14] , 
            \din_i_reg[15] , \delay_i_23__N_1202[15] , \dout_i_23__N_3274[15] , 
            \din_i_reg[16] , \delay_i_23__N_1202[16] , \dout_i_23__N_3274[16] , 
            \din_i_reg[17] , \delay_i_23__N_1202[17] , \dout_i_23__N_3274[17] , 
            \din_i_reg[18] , \delay_i_23__N_1202[18] , \dout_i_23__N_3274[18] , 
            \din_i_reg[23] , \delay_i_23__N_1202[19] , \dout_i_23__N_3274[19] , 
            \delay_i_23__N_1202[20] , \dout_i_23__N_3274[20] , \delay_i_23__N_1202[21] , 
            \dout_i_23__N_3274[21] , \delay_i_23__N_1202[22] , \dout_i_23__N_3274[22] , 
            \delay_i_23__N_1202[23] , \dout_i_23__N_3274[23] , n34659, 
            n34652, n34651, n34650, n34649, n34642, n34641, n34640, 
            n34639, n34630, n34629, n34628, n34627, n34618, n34617, 
            n34616, n34615, n34660, n34661, n34662, n34669, n34670, 
            n34671, n34672, n34675, n34676, n34677, n34678, n34683, 
            n34684, n34685, n34686, valid, clk_c_enable_1419) /* synthesis syn_module_defined=1 */ ;
    input [23:0]op_r_23__N_1106;
    input \count[5] ;
    input \count[4] ;
    input \op_r_23__N_1082[8] ;
    output \radix_no1_op_r[0] ;
    input \op_r_23__N_1082[9] ;
    output \radix_no1_op_r[1] ;
    input GND_net;
    output \op_r_23__N_1268[0] ;
    output \op_r_23__N_1268[1] ;
    output \op_r_23__N_1268[2] ;
    output \op_r_23__N_1268[3] ;
    output \op_r_23__N_1268[4] ;
    output \op_r_23__N_1268[5] ;
    output \op_r_23__N_1268[6] ;
    output \op_r_23__N_1268[7] ;
    output \op_r_23__N_1268[8] ;
    output \op_r_23__N_1268[9] ;
    output \op_r_23__N_1268[10] ;
    output \op_r_23__N_1268[11] ;
    output \op_r_23__N_1268[12] ;
    output \op_r_23__N_1268[13] ;
    output \op_r_23__N_1268[14] ;
    output \op_r_23__N_1268[15] ;
    output \op_r_23__N_1268[16] ;
    output \op_r_23__N_1268[17] ;
    input VCC_net;
    input \op_r_23__N_1082[10] ;
    output \radix_no1_op_r[2] ;
    input \op_r_23__N_1082[11] ;
    output \radix_no1_op_r[3] ;
    input \op_r_23__N_1082[12] ;
    output \radix_no1_op_r[4] ;
    output \op_i_23__N_1310[0] ;
    output \op_i_23__N_1310[1] ;
    output \op_i_23__N_1310[2] ;
    output \op_i_23__N_1310[3] ;
    output \op_i_23__N_1310[4] ;
    output \op_i_23__N_1310[5] ;
    output n89;
    output n88;
    output n87;
    output n86;
    output n85;
    output n84;
    output n83;
    output n82;
    output n81;
    output n80;
    output n79;
    output n78;
    output n77;
    output n76;
    output n75;
    output n74;
    output n73;
    output n72;
    output n71;
    output n70;
    output n69;
    output n68;
    output n67;
    output n66;
    output n65;
    input \rom16_w_i[8] ;
    input n9983;
    input n9984;
    input n9985;
    input n9986;
    input n9987;
    input n9988;
    input \rom16_w_i[0] ;
    input \rom16_w_i[1] ;
    input \rom16_w_i[2] ;
    input \rom16_w_i[3] ;
    input \rom16_w_i[4] ;
    input \rom16_w_i[5] ;
    input \rom16_w_i[6] ;
    input \rom16_w_i[7] ;
    input \op_r_23__N_1082[13] ;
    output \radix_no1_op_r[5] ;
    output \op_r_23__N_1226[0] ;
    output \op_r_23__N_1226[1] ;
    output \op_r_23__N_1226[2] ;
    output \op_r_23__N_1226[3] ;
    output \op_r_23__N_1226[4] ;
    output \op_r_23__N_1226[5] ;
    output \op_r_23__N_1226[6] ;
    output \op_r_23__N_1226[7] ;
    output \op_r_23__N_1226[8] ;
    output \op_r_23__N_1226[9] ;
    output \op_r_23__N_1226[10] ;
    output \op_r_23__N_1226[11] ;
    output \op_r_23__N_1226[12] ;
    output \op_r_23__N_1226[13] ;
    output \op_r_23__N_1226[14] ;
    output \op_r_23__N_1226[15] ;
    output \op_r_23__N_1226[16] ;
    output \op_r_23__N_1226[17] ;
    output \op_r_23__N_1226[18] ;
    output \op_r_23__N_1226[19] ;
    output \op_r_23__N_1226[20] ;
    output \op_r_23__N_1226[21] ;
    output \op_r_23__N_1226[22] ;
    output \op_r_23__N_1226[23] ;
    output \op_r_23__N_1226[24] ;
    output \op_r_23__N_1226[25] ;
    output \op_r_23__N_1226[26] ;
    output \op_r_23__N_1226[27] ;
    output \op_r_23__N_1226[28] ;
    output \op_r_23__N_1226[29] ;
    output \op_r_23__N_1226[30] ;
    output \op_r_23__N_1226[31] ;
    input \op_r_23__N_1082[14] ;
    output \radix_no1_op_r[6] ;
    output \op_r_23__N_1268[18] ;
    output \op_r_23__N_1268[19] ;
    output \op_r_23__N_1268[20] ;
    output \op_r_23__N_1268[21] ;
    output \op_r_23__N_1268[22] ;
    output \op_r_23__N_1268[23] ;
    output \op_r_23__N_1268[24] ;
    output \op_r_23__N_1268[25] ;
    output \op_r_23__N_1268[26] ;
    output \op_r_23__N_1268[27] ;
    output \op_r_23__N_1268[28] ;
    output \op_r_23__N_1268[29] ;
    output \op_r_23__N_1268[30] ;
    output \op_r_23__N_1268[31] ;
    input \rom16_w_r[9] ;
    input n12332;
    input n12333;
    input n12334;
    input n12335;
    input n12336;
    input n12337;
    input n12338;
    input \rom16_w_r[0] ;
    input \rom16_w_r[1] ;
    input \rom16_w_r[2] ;
    input \rom16_w_r[3] ;
    input \rom16_w_r[4] ;
    input \rom16_w_r[5] ;
    input \rom16_w_r[6] ;
    input \rom16_w_r[7] ;
    input \rom16_w_r[8] ;
    input n12314;
    input n12315;
    input n12316;
    input n12317;
    input n12318;
    input n12319;
    input n12320;
    input n12321;
    input n12322;
    input n12323;
    input n12324;
    input n12325;
    input n12326;
    input n12327;
    input n12328;
    input n12329;
    input n12330;
    input n12331;
    input \op_r_23__N_1082[15] ;
    output \radix_no1_op_r[7] ;
    input [23:0]op_i_23__N_1154;
    input \op_i_23__N_1130[8] ;
    output \radix_no1_op_i[0] ;
    input \op_i_23__N_1130[9] ;
    output \radix_no1_op_i[1] ;
    input \op_i_23__N_1130[10] ;
    output \radix_no1_op_i[2] ;
    input \op_i_23__N_1130[11] ;
    output \radix_no1_op_i[3] ;
    input \op_i_23__N_1130[12] ;
    output \radix_no1_op_i[4] ;
    input \op_i_23__N_1130[13] ;
    output \radix_no1_op_i[5] ;
    input \op_i_23__N_1130[14] ;
    output \radix_no1_op_i[6] ;
    input \op_i_23__N_1130[15] ;
    output \radix_no1_op_i[7] ;
    output n8593;
    output n8592;
    output n8591;
    output n8590;
    output n8589;
    output n8588;
    output n8587;
    output n8586;
    output n8585;
    output n8584;
    output n8583;
    output n8582;
    output n8581;
    output n8580;
    output n8579;
    output n8578;
    output n8577;
    output n8576;
    output n8575;
    output n8574;
    output n8573;
    output n8572;
    output n8571;
    output n8570;
    output n8569;
    output n8568;
    input n319;
    input n9989;
    input n9990;
    input n9991;
    input n9992;
    input n9993;
    input n9994;
    input n9995;
    input n9996;
    input n9997;
    input n9998;
    input n9999;
    input n10000;
    input n10001;
    input n10002;
    input n10003;
    input n10004;
    input n10005;
    input n10006;
    input \shift_16_dout_i[8] ;
    input \shift_16_dout_i[9] ;
    input \shift_16_dout_i[10] ;
    input \shift_16_dout_i[11] ;
    input \shift_16_dout_i[12] ;
    input \shift_16_dout_i[13] ;
    input \shift_16_dout_i[14] ;
    input \shift_16_dout_i[15] ;
    input \shift_16_dout_i[16] ;
    input \shift_16_dout_i[17] ;
    input n12344;
    input n12345;
    input n12346;
    input n12347;
    input n12348;
    input n12349;
    input n12350;
    input n12351;
    input n12352;
    input n12353;
    input n12368;
    input \shift_16_dout_i[18] ;
    input \shift_16_dout_i[19] ;
    input \shift_16_dout_i[20] ;
    input \shift_16_dout_i[21] ;
    input \shift_16_dout_i[22] ;
    input \shift_16_dout_i[23] ;
    output clk_c_enable_2310;
    input n34755;
    input \shift_8_dout_r[22] ;
    output n7539;
    input n34756;
    input \op_r_23__N_1082[30] ;
    output n31574;
    input \shift_8_dout_r[23] ;
    output n7538;
    input \op_r_23__N_1082[31] ;
    output n31572;
    input \shift_8_dout_i[22] ;
    output n7486;
    input \op_i_23__N_1130[30] ;
    output n31378;
    input \shift_8_dout_i[23] ;
    output n7485;
    input \op_i_23__N_1130[31] ;
    output n31376;
    input \shift_8_dout_r[20] ;
    output n7541;
    input \op_r_23__N_1082[28] ;
    output n31578;
    input \shift_8_dout_r[21] ;
    output n7540;
    input \op_r_23__N_1082[29] ;
    output n31576;
    input \shift_8_dout_i[20] ;
    output n7488;
    input \op_i_23__N_1130[28] ;
    output n31382;
    input \shift_8_dout_i[21] ;
    output n7487;
    input \op_i_23__N_1130[29] ;
    output n31380;
    input \shift_8_dout_r[18] ;
    output n7543;
    input \op_r_23__N_1082[26] ;
    output n31582;
    input \shift_8_dout_r[19] ;
    output n7542;
    input \op_r_23__N_1082[27] ;
    output n31580;
    input \shift_8_dout_i[18] ;
    output n7490;
    input \op_i_23__N_1130[26] ;
    output n31386;
    input \shift_8_dout_i[19] ;
    output n7489;
    input \op_i_23__N_1130[27] ;
    output n31384;
    input \shift_8_dout_r[16] ;
    output n7545;
    input \op_r_23__N_1082[24] ;
    output n31586;
    input \shift_8_dout_r[17] ;
    output n7544;
    input \op_r_23__N_1082[25] ;
    output n31584;
    input \shift_8_dout_i[16] ;
    output n7492;
    input \op_i_23__N_1130[24] ;
    output n31390;
    input \shift_8_dout_i[17] ;
    output n7491;
    input \op_i_23__N_1130[25] ;
    output n31388;
    input \shift_8_dout_r[14] ;
    output n7547;
    input \op_r_23__N_1082[22] ;
    output n31590;
    input \shift_8_dout_r[15] ;
    output n7546;
    input \op_r_23__N_1082[23] ;
    output n31588;
    input \shift_8_dout_i[14] ;
    output n7494;
    input \op_i_23__N_1130[22] ;
    output n31394;
    input \shift_8_dout_i[15] ;
    output n7493;
    input \op_i_23__N_1130[23] ;
    output n31392;
    input \shift_8_dout_r[12] ;
    output n7549;
    input \op_r_23__N_1082[20] ;
    output n31594;
    input \shift_8_dout_r[13] ;
    output n7548;
    input \op_r_23__N_1082[21] ;
    output n31592;
    input \shift_8_dout_i[12] ;
    output n7496;
    input \op_i_23__N_1130[20] ;
    output n31398;
    input \shift_8_dout_i[13] ;
    output n7495;
    input \op_i_23__N_1130[21] ;
    output n31396;
    input \shift_8_dout_r[10] ;
    output n7551;
    input \op_r_23__N_1082[18] ;
    output n31598;
    input \shift_8_dout_r[11] ;
    output n7550;
    input \op_r_23__N_1082[19] ;
    output n31596;
    input \shift_8_dout_i[10] ;
    output n7498;
    input \op_i_23__N_1130[18] ;
    output n31402;
    input \shift_8_dout_i[11] ;
    output n7497;
    input \op_i_23__N_1130[19] ;
    output n31400;
    input \shift_8_dout_r[8] ;
    output n7553;
    input \op_r_23__N_1082[16] ;
    output n31602;
    input \shift_8_dout_r[9] ;
    output n7552;
    input \op_r_23__N_1082[17] ;
    output n31600;
    input \shift_8_dout_i[8] ;
    output n7500;
    input \op_i_23__N_1130[16] ;
    output n31406;
    input \shift_8_dout_i[9] ;
    output n7499;
    input \op_i_23__N_1130[17] ;
    output n31404;
    input \din_r_reg[8] ;
    input \delay_r_23__N_1178[8] ;
    output \dout_r_23__N_2506[8] ;
    input \din_r_reg[9] ;
    input \delay_r_23__N_1178[9] ;
    output \dout_r_23__N_2506[9] ;
    input \din_r_reg[10] ;
    input \delay_r_23__N_1178[10] ;
    output \dout_r_23__N_2506[10] ;
    input \din_r_reg[11] ;
    input \delay_r_23__N_1178[11] ;
    output \dout_r_23__N_2506[11] ;
    input \din_r_reg[12] ;
    input \delay_r_23__N_1178[12] ;
    output \dout_r_23__N_2506[12] ;
    input \din_r_reg[13] ;
    input \delay_r_23__N_1178[13] ;
    output \dout_r_23__N_2506[13] ;
    input \din_r_reg[14] ;
    input \delay_r_23__N_1178[14] ;
    output \dout_r_23__N_2506[14] ;
    input \din_r_reg[15] ;
    input \delay_r_23__N_1178[15] ;
    output \dout_r_23__N_2506[15] ;
    input \din_r_reg[16] ;
    input \delay_r_23__N_1178[16] ;
    output \dout_r_23__N_2506[16] ;
    input \din_r_reg[17] ;
    input \delay_r_23__N_1178[17] ;
    output \dout_r_23__N_2506[17] ;
    input \din_r_reg[18] ;
    input \delay_r_23__N_1178[18] ;
    output \dout_r_23__N_2506[18] ;
    input \din_r_reg[23] ;
    input \delay_r_23__N_1178[19] ;
    output \dout_r_23__N_2506[19] ;
    input \delay_r_23__N_1178[20] ;
    output \dout_r_23__N_2506[20] ;
    input \delay_r_23__N_1178[21] ;
    output \dout_r_23__N_2506[21] ;
    input \delay_r_23__N_1178[22] ;
    output \dout_r_23__N_2506[22] ;
    input \delay_r_23__N_1178[23] ;
    output \dout_r_23__N_2506[23] ;
    input \din_i_reg[8] ;
    input \delay_i_23__N_1202[8] ;
    output \dout_i_23__N_3274[8] ;
    input \din_i_reg[9] ;
    input \delay_i_23__N_1202[9] ;
    output \dout_i_23__N_3274[9] ;
    input \din_i_reg[10] ;
    input \delay_i_23__N_1202[10] ;
    output \dout_i_23__N_3274[10] ;
    input \din_i_reg[11] ;
    input \delay_i_23__N_1202[11] ;
    output \dout_i_23__N_3274[11] ;
    input \din_i_reg[12] ;
    input \delay_i_23__N_1202[12] ;
    output \dout_i_23__N_3274[12] ;
    input \din_i_reg[13] ;
    input \delay_i_23__N_1202[13] ;
    output \dout_i_23__N_3274[13] ;
    input \din_i_reg[14] ;
    input \delay_i_23__N_1202[14] ;
    output \dout_i_23__N_3274[14] ;
    input \din_i_reg[15] ;
    input \delay_i_23__N_1202[15] ;
    output \dout_i_23__N_3274[15] ;
    input \din_i_reg[16] ;
    input \delay_i_23__N_1202[16] ;
    output \dout_i_23__N_3274[16] ;
    input \din_i_reg[17] ;
    input \delay_i_23__N_1202[17] ;
    output \dout_i_23__N_3274[17] ;
    input \din_i_reg[18] ;
    input \delay_i_23__N_1202[18] ;
    output \dout_i_23__N_3274[18] ;
    input \din_i_reg[23] ;
    input \delay_i_23__N_1202[19] ;
    output \dout_i_23__N_3274[19] ;
    input \delay_i_23__N_1202[20] ;
    output \dout_i_23__N_3274[20] ;
    input \delay_i_23__N_1202[21] ;
    output \dout_i_23__N_3274[21] ;
    input \delay_i_23__N_1202[22] ;
    output \dout_i_23__N_3274[22] ;
    input \delay_i_23__N_1202[23] ;
    output \dout_i_23__N_3274[23] ;
    output n34659;
    output n34652;
    output n34651;
    output n34650;
    output n34649;
    output n34642;
    output n34641;
    output n34640;
    output n34639;
    output n34630;
    output n34629;
    output n34628;
    output n34627;
    output n34618;
    output n34617;
    output n34616;
    output n34615;
    output n34660;
    output n34661;
    output n34662;
    output n34669;
    output n34670;
    output n34671;
    output n34672;
    output n34675;
    output n34676;
    output n34677;
    output n34678;
    output n34683;
    output n34684;
    output n34685;
    output n34686;
    input valid;
    output clk_c_enable_1419;
    
    
    wire n18090, n18091, n18092, n18093, n18094, n18095, n18096, 
        n18097, n18098, n18099, n18100, n18101, n18102, n18103, 
        n18104, n18105, n18106, n18107, n18108, n18109, n18110, 
        n18111, n18112, n18113, n18114, n18115, n18116, n18117, 
        n18118, n18119, n18120, n18121, n18122, n18123, n18124, 
        n18125, n18126, n18127, n18128, n18129, n18130, n18131, 
        n18132, n18133, n18134, n18135, n18136, n18137, n18138, 
        n18139, n18140, n18141, n18142, n18143, n18144, n18145, 
        n18146, n18147, n18148, n18149, n18150, n18151, n18152, 
        n18153, n18154, n18155, n18156, n18157, n18158, n18159, 
        n18160, n18161, n18162, n18163, n18164, n18165, n18166, 
        n18167, n18168, n18169, n18170, n18171, n18172, n18173, 
        n18174, n18175, n18176, n18177, n18178, n18179, n18180, 
        n18181, n18182, n18183, n18184, n18185, n18186, n18187, 
        n18188, n18189, n18190, n18191, n18192, n18193, n18194, 
        n18195, n18196, n18197, n18198, n18199, n18200, n18201, 
        n18202, n18203, n18204, n18205, n18206, n18207, n18208, 
        n18209, n18210, n18211, n18212, n18213, n18214, n18215, 
        n18216, n18217, n18218, n18219, n18220, n18221, n18222, 
        n18223, n18224, n18225, n18226, n18227, n18228, n18229, 
        n18230, n18231, n18232, n18233, n18234, n18235, n18382, 
        n18383, n18384, n18385, n18386, n18387, n18388, n18389, 
        n18390, n18391, n18392, n18393, n18394, n18395, n18396, 
        n18397, n18398, n18399, n18400, n18401, n18402, n18403, 
        n18404, n18405, n18406, n18407, n18408, n18409, n18410, 
        n18411, n18412, n18413, n18414, n18415, n18416, n18417, 
        n18418, n18565, n18566, n18567, n18568, n18569, n18570, 
        n18571, n18572, n18573, n18574, n18575, n18576, n18577, 
        n18578, n18579, n18580, n18581, n18582, n18583, n18584, 
        n18585, n18586, n18587, n18588, n18589, n18590, n18591, 
        n18592, n18593, n18594, n18595, n18596, n18597, n18598, 
        n18599, n18600, n18601, n18602, n18603, n18604, n18605, 
        n18606, n18607, n18608, n18609, n18610, n18611, n18612, 
        n18613, n18614, n18615, n18616, n18617, n18618, n18619, 
        n18620, n18621, n18622, n18623, n18624, n18625, n18626, 
        n18627, n18628, n18629, n18630, n18631, n18632, n18633, 
        n18634, n18635, n18636, n18637, n18638, n18639, n18640, 
        n18641, n18642, n18643, n18644, n18645, n18646, n18647, 
        n18648, n18649, n18650, n18651, n18652, n18653, n18654, 
        n18655, n18656, n18657, n18658, n18659, n18660, n18661, 
        n18662, n18663, n18664, n18665, n18666, n18667, n18668, 
        n18669, n18670, n18671, n18672, n18673, n18674, n18675, 
        n18676, n18677, n18678, n18679, n18680, n18681, n18682, 
        n18683, n18684, n18685, n18686, n18687, n18688, n18689, 
        n18690, n18691, n18692, n18693, n18694, n18695, n18696, 
        n18697, n18698, n18699, n18700, n18701, n18702, n18703, 
        n18704, n18705, n18706, n18707, n18708, n18709, n18710, 
        n15122, n15123, n15124, n15125, n15126, n15127, n15128, 
        n15129, n15130, n15131, n15132, n15133, n15134, n15135, 
        n15136, n15137, n15138, n15139, n15140, n15141, n15142, 
        n15143, n15144, n15145, n15146, n15147, n15148, n15149, 
        n15150, n15151, n15152, n15153, n15154, n15155, n15156, 
        n15157, n15158, n15159, n15160, n15161, n15162, n15163, 
        n15164, n15165, n15166, n15167, n15168, n15169, n15170, 
        n15171, n15172, n15173, n15174, n15175, n15176, n15177, 
        n15178, n15179, n15180, n15181, n15182, n15183, n15184, 
        n15185, n15186, n15187, n15188, n15189, n15190, n15191, 
        n15192, n15193, n15194, n15195, n15196, n15197, n15198, 
        n15199, n15200, n15201, n15202, n15203, n15204, n15205, 
        n15206, n15207, n15208, n15209, n15210, n15211, n15212, 
        n15213, n15214, n15215, n15216, n15217, n15218, n15219, 
        n15220, n15221, n15222, n15223, n15224, n15225, n15226, 
        n15227, n15228, n15229, n15230, n15231, n15232, n15233, 
        n15234, n15235, n15236, n15237, n15238, n15239, n15240, 
        n15241, n15242, n15243, n15244, n15245, n15246, n15247, 
        n15248, n15249, n15250, n15251, n15252, n15253, n15254, 
        n15255, n15256, n15257, n15258, n15259, n15260, n15261, 
        n15262, n15263, n15264, n15265, n15266, n15267, n15268, 
        n15269, n15270, n15271, n15272, n15273, n15274, n15275, 
        n15276, n15277, n15278, n15279, n15280, n15281, n15282, 
        n15283, n15284, n15285, n15286, n15287, n15288, n15289, 
        n15290, n15291, n15292, n15293, n15294, n15295, n15296, 
        n15297, n15298, n15299, n15300, n15301, n15302, n15303, 
        n15304, n14976, n14977, n14978, n14979, n14980, n14981, 
        n14982, n14983, n14984, n14985, n14986, n14987, n14988, 
        n14989, n14990, n14991, n14992, n14993, n14994, n14995, 
        n14996, n14997, n14998, n14999, n15000, n15001, n15002, 
        n15003, n15004, n15005, n15006, n15007, n15008, n15009, 
        n15010, n15011, n15012, n15013, n15014, n15015, n15016, 
        n15017, n15018, n15019, n15020, n15021, n15022, n15023, 
        n15024, n15025, n15026, n15027, n15028, n15029, n15030, 
        n15031, n15032, n15033, n15034, n15035, n15036, n15037, 
        n15038, n15039, n15040, n15041, n15042, n15043, n15044, 
        n15045, n15046, n15047, n15048, n15049, n15050, n15051, 
        n15052, n15053, n15054, n15055, n15056, n15057, n15058, 
        n15059, n15060, n15061, n15062, n15063, n15064, n15065, 
        n15066, n15067, n15068, n15069, n15070, n15071, n15072, 
        n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
        n15080, n15081, n15082, n15083, n15084, n15085, n15086, 
        n15087, n15088, n15089, n15090, n15091, n15092, n15093, 
        n15094, n15095, n15096, n15097, n15098, n15099, n15100, 
        n15101, n15102, n15103, n15104, n15105, n15106, n15107, 
        n15108, n15109, n15110, n15111, n15112, n15113, n15114, 
        n15115, n15116, n15117, n15118, n15119, n15120, n15121, 
        n18236, n18237, n18238, n18239, n18240, n18241, n18242, 
        n18243, n18244, n18245, n18246, n18247, n18248, n18249, 
        n18250, n18251, n18252, n18253, n18254, n18255, n18256, 
        n18257, n18258, n18259, n18260, n18261, n18262, n18263, 
        n18264, n18265, n18266, n18267, n18268, n18269, n18270, 
        n18271, n18272, n18273, n18274, n18275, n18276, n18277, 
        n18278, n18279, n18280, n18281, n18282, n18283, n18284, 
        n18285, n18286, n18287, n18288, n18289, n18290, n18291, 
        n18292, n18293, n18294, n18295, n18296, n18297, n18298, 
        n18299, n18300, n18301, n18302, n18303, n18304, n18305, 
        n18306, n18307, n18308, n18309, n18310, n18311, n18312, 
        n18313, n18314, n18315, n18316, n18317, n18318, n18319, 
        n18320, n18321, n18322, n18323, n18324, n18325, n18326, 
        n18327, n18328, n18329, n18330, n18331, n18332, n18333, 
        n18334, n18335, n18336, n18337, n18338, n18339, n18340, 
        n18341, n18342, n18343, n18344, n18345, n18346, n18347, 
        n18348, n18349, n18350, n18351, n18352, n18353, n18354, 
        n18355, n18356, n18357, n18358, n18359, n18360, n18361, 
        n18362, n18363, n18364, n18365, n18366, n18367, n18368, 
        n18369, n18370, n18371, n18372, n18373, n18374, n18375, 
        n18376, n18377, n18378, n18379, n18380, n18381, n13324, 
        n13325, n13326, n13327, n13328, n13329, n13330, n13331, 
        n13332, n13333, n13334, n13335, n13336, n13337, n13338, 
        n13339, n13340, n13341, n13342, n13343, n13344, n13345, 
        n13346, n13347, n13348, n13349, n13350, n13351, n13352, 
        n13353, n13354, n13355, n13356, n13357, n13358, n13359, 
        n13360, n13361, n13362, n13363, n13364, n13365, n13366, 
        n13367, n13368, n13369, n13370, n13371, n13372, n13373, 
        n13374, n13375, n13376, n13377, n13378, n13379, n13380, 
        n13381, n13382, n13383, n13384, n13385, n13386, n13387, 
        n13388, n13389, n13390, n13391, n13392, n13393, n13394, 
        n13395, n13396, n13397, n13398, n13399, n13400, n13401, 
        n13402, n13403, n13404, n13405, n13406, n13407, n13408, 
        n13409, n13410, n13411, n13412, n13413, n13414, n13415, 
        n13416, n13417, n13418, n13419, n13420, n13421, n13422, 
        n13423, n13424, n13425, n13426, n13427, n13428, n13429, 
        n13430, n13431, n13432, n13433, n13434, n13435, n13436, 
        n13437, n13438, n13439, n13440, n13441, n13442, n13443, 
        n13444, n13445, n13446, n13447, n13448, n13449, n13450, 
        n13451, n13452, n13453, n13454, n13455, n13456, n13457, 
        n13458, n13459, n13460, n13461, n13462, n13463, n13464, 
        n13465, n13466, n13467, n13468, n13469, n13470, n13471, 
        n13472, n13473, n13474, n13475, n13476, n13477, n13478, 
        n13479, n13480, n13481, n13482, n13483, n13484, n13485, 
        n13486, n13487, n13488, n13489, n13490, n13491, n13492, 
        n13493, n13494, n13495, n13496, n13497, n13498, n13499, 
        n13500, n13501, n13502, n13503, n13504, n13505, n13506, 
        n13178, n13179, n13180, n13181, n13182, n13183, n13184, 
        n13185, n13186, n13187, n13188, n13189, n13190, n13191, 
        n13192, n13193, n13194, n13195, n13196, n13197, n13198, 
        n13199, n13200, n13201, n13202, n13203, n13204, n13205, 
        n13206, n13207, n13208, n13209, n13210, n13211, n13212, 
        n13213, n13214, n13215, n13216, n13217, n13218, n13219, 
        n13220, n13221, n13222, n13223, n13224, n13225, n13226, 
        n13227, n13228, n13229, n13230, n13231, n13232, n13233, 
        n13234, n13235, n13236, n13237, n13238, n13239, n13240, 
        n13241, n13242, n13243, n13244, n13245, n13246, n13247, 
        n13248, n13249, n13250, n13251, n13252, n13253, n13254, 
        n13255, n13256, n13257, n13258, n13259, n13260, n13261, 
        n13262, n13263, n13264, n13265, n13266, n13267, n13268, 
        n13269, n13270, n13271, n13272, n13273, n13274, n13275, 
        n13276, n13277, n13278, n13279, n13280, n13281, n13282, 
        n13283, n13284, n13285, n13286, n13287, n13288, n13289, 
        n13290, n13291, n13292, n13293, n13294, n13295, n13296, 
        n13297, n13298, n13299, n13300, n13301, n13302, n13303, 
        n13304, n13305, n13306, n13307, n13308, n13309, n13310, 
        n13311, n13312, n13313, n13314, n13315, n13316, n13317, 
        n13318, n13319, n13320, n13321, n13322, n13323;
    
    LUT4 i12536_4_lut_4_lut (.A(op_r_23__N_1106[0]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[8] ), .Z(\radix_no1_op_r[0] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12536_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12825_4_lut_4_lut (.A(op_r_23__N_1106[1]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[9] ), .Z(\radix_no1_op_r[1] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12825_4_lut_4_lut.init = 16'h2c20;
    ALU54B lat_alu_73 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18126), .SIGNEDIB(n18199), .SIGNEDCIN(GND_net), 
           .A35(n18125), .A34(n18124), .A33(n18123), .A32(n18122), .A31(n18121), 
           .A30(n18120), .A29(n18119), .A28(n18118), .A27(n18117), .A26(n18116), 
           .A25(n18115), .A24(n18114), .A23(n18113), .A22(n18112), .A21(n18111), 
           .A20(n18110), .A19(n18109), .A18(n18108), .A17(n18107), .A16(n18106), 
           .A15(n18105), .A14(n18104), .A13(n18103), .A12(n18102), .A11(n18101), 
           .A10(n18100), .A9(n18099), .A8(n18098), .A7(n18097), .A6(n18096), 
           .A5(n18095), .A4(n18094), .A3(n18093), .A2(n18092), .A1(n18091), 
           .A0(n18090), .B35(n18198), .B34(n18197), .B33(n18196), .B32(n18195), 
           .B31(n18194), .B30(n18193), .B29(n18192), .B28(n18191), .B27(n18190), 
           .B26(n18189), .B25(n18188), .B24(n18187), .B23(n18186), .B22(n18185), 
           .B21(n18184), .B20(n18183), .B19(n18182), .B18(n18181), .B17(n18180), 
           .B16(n18179), .B15(n18178), .B14(n18177), .B13(n18176), .B12(n18175), 
           .B11(n18174), .B10(n18173), .B9(n18172), .B8(n18171), .B7(n18170), 
           .B6(n18169), .B5(n18168), .B4(n18167), .B3(n18166), .B2(n18165), 
           .B1(n18164), .B0(n18163), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18162), .MA34(n18161), .MA33(n18160), .MA32(n18159), 
           .MA31(n18158), .MA30(n18157), .MA29(n18156), .MA28(n18155), 
           .MA27(n18154), .MA26(n18153), .MA25(n18152), .MA24(n18151), 
           .MA23(n18150), .MA22(n18149), .MA21(n18148), .MA20(n18147), 
           .MA19(n18146), .MA18(n18145), .MA17(n18144), .MA16(n18143), 
           .MA15(n18142), .MA14(n18141), .MA13(n18140), .MA12(n18139), 
           .MA11(n18138), .MA10(n18137), .MA9(n18136), .MA8(n18135), 
           .MA7(n18134), .MA6(n18133), .MA5(n18132), .MA4(n18131), .MA3(n18130), 
           .MA2(n18129), .MA1(n18128), .MA0(n18127), .MB35(n18235), 
           .MB34(n18234), .MB33(n18233), .MB32(n18232), .MB31(n18231), 
           .MB30(n18230), .MB29(n18229), .MB28(n18228), .MB27(n18227), 
           .MB26(n18226), .MB25(n18225), .MB24(n18224), .MB23(n18223), 
           .MB22(n18222), .MB21(n18221), .MB20(n18220), .MB19(n18219), 
           .MB18(n18218), .MB17(n18217), .MB16(n18216), .MB15(n18215), 
           .MB14(n18214), .MB13(n18213), .MB12(n18212), .MB11(n18211), 
           .MB10(n18210), .MB9(n18209), .MB8(n18208), .MB7(n18207), 
           .MB6(n18206), .MB5(n18205), .MB4(n18204), .MB3(n18203), .MB2(n18202), 
           .MB1(n18201), .MB0(n18200), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n18417), 
           .R52(n18416), .R51(n18415), .R50(n18414), .R49(n18413), .R48(n18412), 
           .R47(n18411), .R46(n18410), .R45(n18409), .R44(n18408), .R43(n18407), 
           .R42(n18406), .R41(n18405), .R40(n18404), .R39(n18403), .R38(n18402), 
           .R37(n18401), .R36(n18400), .R35(n18399), .R34(n18398), .R33(n18397), 
           .R32(n18396), .R31(n18395), .R30(n18394), .R29(n18393), .R28(n18392), 
           .R27(n18391), .R26(n18390), .R25(n18389), .R24(n18388), .R23(n18387), 
           .R22(n18386), .R21(n18385), .R20(n18384), .R19(n18383), .R18(n18382), 
           .R17(\op_r_23__N_1268[17] ), .R16(\op_r_23__N_1268[16] ), .R15(\op_r_23__N_1268[15] ), 
           .R14(\op_r_23__N_1268[14] ), .R13(\op_r_23__N_1268[13] ), .R12(\op_r_23__N_1268[12] ), 
           .R11(\op_r_23__N_1268[11] ), .R10(\op_r_23__N_1268[10] ), .R9(\op_r_23__N_1268[9] ), 
           .R8(\op_r_23__N_1268[8] ), .R7(\op_r_23__N_1268[7] ), .R6(\op_r_23__N_1268[6] ), 
           .R5(\op_r_23__N_1268[5] ), .R4(\op_r_23__N_1268[4] ), .R3(\op_r_23__N_1268[3] ), 
           .R2(\op_r_23__N_1268[2] ), .R1(\op_r_23__N_1268[1] ), .R0(\op_r_23__N_1268[0] ), 
           .SIGNEDR(n18418));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_73.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_73.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_73.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_73.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_73.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_73.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_73.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_73.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_73.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_73.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_73.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_73.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_73.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_73.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_73.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_73.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_73.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_73.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_73.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_73.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_73.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_73.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_73.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_73.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_73.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_73.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_73.REG_FLAG_CLK = "NONE";
    defparam lat_alu_73.REG_FLAG_CE = "CE0";
    defparam lat_alu_73.REG_FLAG_RST = "RST0";
    defparam lat_alu_73.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_73.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_73.MASK01 = "0x00000000000000";
    defparam lat_alu_73.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_73.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_73.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_73.CLK0_DIV = "ENABLED";
    defparam lat_alu_73.CLK1_DIV = "ENABLED";
    defparam lat_alu_73.CLK2_DIV = "ENABLED";
    defparam lat_alu_73.CLK3_DIV = "ENABLED";
    defparam lat_alu_73.MCPAT = "0x00000000000000";
    defparam lat_alu_73.MASKPAT = "0x00000000000000";
    defparam lat_alu_73.RNDPAT = "0x00000000000000";
    defparam lat_alu_73.GSR = "DISABLED";
    defparam lat_alu_73.RESETMODE = "SYNC";
    defparam lat_alu_73.MULT9_MODE = "DISABLED";
    defparam lat_alu_73.LEGACY = "DISABLED";
    LUT4 i12826_4_lut_4_lut (.A(op_r_23__N_1106[2]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[10] ), .Z(\radix_no1_op_r[2] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12826_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12827_4_lut_4_lut (.A(op_r_23__N_1106[3]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[11] ), .Z(\radix_no1_op_r[3] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12827_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12828_4_lut_4_lut (.A(op_r_23__N_1106[4]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[12] ), .Z(\radix_no1_op_r[4] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12828_4_lut_4_lut.init = 16'h2c20;
    ALU54B lat_alu_78 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18601), .SIGNEDIB(n18674), .SIGNEDCIN(GND_net), 
           .A35(n18600), .A34(n18599), .A33(n18598), .A32(n18597), .A31(n18596), 
           .A30(n18595), .A29(n18594), .A28(n18593), .A27(n18592), .A26(n18591), 
           .A25(n18590), .A24(n18589), .A23(n18588), .A22(n18587), .A21(n18586), 
           .A20(n18585), .A19(n18584), .A18(n18583), .A17(n18582), .A16(n18581), 
           .A15(n18580), .A14(n18579), .A13(n18578), .A12(n18577), .A11(n18576), 
           .A10(n18575), .A9(n18574), .A8(n18573), .A7(n18572), .A6(n18571), 
           .A5(n18570), .A4(n18569), .A3(n18568), .A2(n18567), .A1(n18566), 
           .A0(n18565), .B35(n18673), .B34(n18672), .B33(n18671), .B32(n18670), 
           .B31(n18669), .B30(n18668), .B29(n18667), .B28(n18666), .B27(n18665), 
           .B26(n18664), .B25(n18663), .B24(n18662), .B23(n18661), .B22(n18660), 
           .B21(n18659), .B20(n18658), .B19(n18657), .B18(n18656), .B17(n18655), 
           .B16(n18654), .B15(n18653), .B14(n18652), .B13(n18651), .B12(n18650), 
           .B11(n18649), .B10(n18648), .B9(n18647), .B8(n18646), .B7(n18645), 
           .B6(n18644), .B5(n18643), .B4(n18642), .B3(n18641), .B2(n18640), 
           .B1(n18639), .B0(n18638), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18637), .MA34(n18636), .MA33(n18635), .MA32(n18634), 
           .MA31(n18633), .MA30(n18632), .MA29(n18631), .MA28(n18630), 
           .MA27(n18629), .MA26(n18628), .MA25(n18627), .MA24(n18626), 
           .MA23(n18625), .MA22(n18624), .MA21(n18623), .MA20(n18622), 
           .MA19(n18621), .MA18(n18620), .MA17(n18619), .MA16(n18618), 
           .MA15(n18617), .MA14(n18616), .MA13(n18615), .MA12(n18614), 
           .MA11(n18613), .MA10(n18612), .MA9(n18611), .MA8(n18610), 
           .MA7(n18609), .MA6(n18608), .MA5(n18607), .MA4(n18606), .MA3(n18605), 
           .MA2(n18604), .MA1(n18603), .MA0(n18602), .MB35(n18710), 
           .MB34(n18709), .MB33(n18708), .MB32(n18707), .MB31(n18706), 
           .MB30(n18705), .MB29(n18704), .MB28(n18703), .MB27(n18702), 
           .MB26(n18701), .MB25(n18700), .MB24(n18699), .MB23(n18698), 
           .MB22(n18697), .MB21(n18696), .MB20(n18695), .MB19(n18694), 
           .MB18(n18693), .MB17(n18692), .MB16(n18691), .MB15(n18690), 
           .MB14(n18689), .MB13(n18688), .MB12(n18687), .MB11(n18686), 
           .MB10(n18685), .MB9(n18684), .MB8(n18683), .MB7(n18682), 
           .MB6(n18681), .MB5(n18680), .MB4(n18679), .MB3(n18678), .MB2(n18677), 
           .MB1(n18676), .MB0(n18675), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R30(n65), .R29(n66), 
           .R28(n67), .R27(n68), .R26(n69), .R25(n70), .R24(n71), 
           .R23(n72), .R22(n73), .R21(n74), .R20(n75), .R19(n76), 
           .R18(n77), .R17(n78), .R16(n79), .R15(n80), .R14(n81), 
           .R13(n82), .R12(n83), .R11(n84), .R10(n85), .R9(n86), .R8(n87), 
           .R7(n88), .R6(n89), .R5(\op_i_23__N_1310[5] ), .R4(\op_i_23__N_1310[4] ), 
           .R3(\op_i_23__N_1310[3] ), .R2(\op_i_23__N_1310[2] ), .R1(\op_i_23__N_1310[1] ), 
           .R0(\op_i_23__N_1310[0] ));
    defparam lat_alu_78.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_78.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_78.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_78.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_78.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_78.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_78.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_78.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_78.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_78.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_78.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_78.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_78.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_78.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_78.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_78.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_78.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_78.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_78.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_78.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_78.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_78.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_78.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_78.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_78.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_78.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_78.REG_FLAG_CLK = "NONE";
    defparam lat_alu_78.REG_FLAG_CE = "CE0";
    defparam lat_alu_78.REG_FLAG_RST = "RST0";
    defparam lat_alu_78.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_78.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_78.MASK01 = "0x00000000000000";
    defparam lat_alu_78.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_78.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_78.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_78.CLK0_DIV = "ENABLED";
    defparam lat_alu_78.CLK1_DIV = "ENABLED";
    defparam lat_alu_78.CLK2_DIV = "ENABLED";
    defparam lat_alu_78.CLK3_DIV = "ENABLED";
    defparam lat_alu_78.MCPAT = "0x00000000000000";
    defparam lat_alu_78.MASKPAT = "0x00000000000000";
    defparam lat_alu_78.RNDPAT = "0x00000000000000";
    defparam lat_alu_78.GSR = "DISABLED";
    defparam lat_alu_78.RESETMODE = "SYNC";
    defparam lat_alu_78.MULT9_MODE = "DISABLED";
    defparam lat_alu_78.LEGACY = "DISABLED";
    MULT18X18D lat_mult_77 (.A17(\rom16_w_i[8] ), .A16(\rom16_w_i[8] ), 
            .A15(\rom16_w_i[8] ), .A14(\rom16_w_i[8] ), .A13(\rom16_w_i[8] ), 
            .A12(\rom16_w_i[8] ), .A11(\rom16_w_i[8] ), .A10(\rom16_w_i[8] ), 
            .A9(\rom16_w_i[8] ), .A8(\rom16_w_i[8] ), .A7(\rom16_w_i[8] ), 
            .A6(\rom16_w_i[8] ), .A5(\rom16_w_i[8] ), .A4(\rom16_w_i[8] ), 
            .A3(\rom16_w_i[8] ), .A2(\rom16_w_i[8] ), .A1(\rom16_w_i[8] ), 
            .A0(\rom16_w_i[8] ), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(GND_net), .B7(GND_net), 
            .B6(GND_net), .B5(n9988), .B4(n9987), .B3(n9986), .B2(n9985), 
            .B1(n9984), .B0(n9983), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18655), 
            .ROA16(n18654), .ROA15(n18653), .ROA14(n18652), .ROA13(n18651), 
            .ROA12(n18650), .ROA11(n18649), .ROA10(n18648), .ROA9(n18647), 
            .ROA8(n18646), .ROA7(n18645), .ROA6(n18644), .ROA5(n18643), 
            .ROA4(n18642), .ROA3(n18641), .ROA2(n18640), .ROA1(n18639), 
            .ROA0(n18638), .ROB17(n18673), .ROB16(n18672), .ROB15(n18671), 
            .ROB14(n18670), .ROB13(n18669), .ROB12(n18668), .ROB11(n18667), 
            .ROB10(n18666), .ROB9(n18665), .ROB8(n18664), .ROB7(n18663), 
            .ROB6(n18662), .ROB5(n18661), .ROB4(n18660), .ROB3(n18659), 
            .ROB2(n18658), .ROB1(n18657), .ROB0(n18656), .P35(n18710), 
            .P34(n18709), .P33(n18708), .P32(n18707), .P31(n18706), 
            .P30(n18705), .P29(n18704), .P28(n18703), .P27(n18702), 
            .P26(n18701), .P25(n18700), .P24(n18699), .P23(n18698), 
            .P22(n18697), .P21(n18696), .P20(n18695), .P19(n18694), 
            .P18(n18693), .P17(n18692), .P16(n18691), .P15(n18690), 
            .P14(n18689), .P13(n18688), .P12(n18687), .P11(n18686), 
            .P10(n18685), .P9(n18684), .P8(n18683), .P7(n18682), .P6(n18681), 
            .P5(n18680), .P4(n18679), .P3(n18678), .P2(n18677), .P1(n18676), 
            .P0(n18675), .SIGNEDP(n18674));
    defparam lat_mult_77.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_77.REG_INPUTA_CE = "CE0";
    defparam lat_mult_77.REG_INPUTA_RST = "RST0";
    defparam lat_mult_77.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_77.REG_INPUTB_CE = "CE0";
    defparam lat_mult_77.REG_INPUTB_RST = "RST0";
    defparam lat_mult_77.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_77.REG_INPUTC_CE = "CE0";
    defparam lat_mult_77.REG_INPUTC_RST = "RST0";
    defparam lat_mult_77.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_77.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_77.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_77.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_77.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_77.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_77.CLK0_DIV = "ENABLED";
    defparam lat_mult_77.CLK1_DIV = "ENABLED";
    defparam lat_mult_77.CLK2_DIV = "ENABLED";
    defparam lat_mult_77.CLK3_DIV = "ENABLED";
    defparam lat_mult_77.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_77.GSR = "DISABLED";
    defparam lat_mult_77.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_77.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_77.MULT_BYPASS = "DISABLED";
    defparam lat_mult_77.RESETMODE = "SYNC";
    MULT18X18D mult_967_mult_2 (.A17(\rom16_w_i[8] ), .A16(\rom16_w_i[8] ), 
            .A15(\rom16_w_i[8] ), .A14(\rom16_w_i[8] ), .A13(\rom16_w_i[8] ), 
            .A12(\rom16_w_i[8] ), .A11(\rom16_w_i[8] ), .A10(\rom16_w_i[8] ), 
            .A9(\rom16_w_i[8] ), .A8(\rom16_w_i[8] ), .A7(\rom16_w_i[7] ), 
            .A6(\rom16_w_i[6] ), .A5(\rom16_w_i[5] ), .A4(\rom16_w_i[4] ), 
            .A3(\rom16_w_i[3] ), .A2(\rom16_w_i[2] ), .A1(\rom16_w_i[1] ), 
            .A0(\rom16_w_i[0] ), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(GND_net), .B7(GND_net), 
            .B6(GND_net), .B5(n9988), .B4(n9987), .B3(n9986), .B2(n9985), 
            .B1(n9984), .B0(n9983), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18582), 
            .ROA16(n18581), .ROA15(n18580), .ROA14(n18579), .ROA13(n18578), 
            .ROA12(n18577), .ROA11(n18576), .ROA10(n18575), .ROA9(n18574), 
            .ROA8(n18573), .ROA7(n18572), .ROA6(n18571), .ROA5(n18570), 
            .ROA4(n18569), .ROA3(n18568), .ROA2(n18567), .ROA1(n18566), 
            .ROA0(n18565), .ROB17(n18600), .ROB16(n18599), .ROB15(n18598), 
            .ROB14(n18597), .ROB13(n18596), .ROB12(n18595), .ROB11(n18594), 
            .ROB10(n18593), .ROB9(n18592), .ROB8(n18591), .ROB7(n18590), 
            .ROB6(n18589), .ROB5(n18588), .ROB4(n18587), .ROB3(n18586), 
            .ROB2(n18585), .ROB1(n18584), .ROB0(n18583), .P35(n18637), 
            .P34(n18636), .P33(n18635), .P32(n18634), .P31(n18633), 
            .P30(n18632), .P29(n18631), .P28(n18630), .P27(n18629), 
            .P26(n18628), .P25(n18627), .P24(n18626), .P23(n18625), 
            .P22(n18624), .P21(n18623), .P20(n18622), .P19(n18621), 
            .P18(n18620), .P17(n18619), .P16(n18618), .P15(n18617), 
            .P14(n18616), .P13(n18615), .P12(n18614), .P11(n18613), 
            .P10(n18612), .P9(n18611), .P8(n18610), .P7(n18609), .P6(n18608), 
            .P5(n18607), .P4(n18606), .P3(n18605), .P2(n18604), .P1(n18603), 
            .P0(n18602), .SIGNEDP(n18601));
    defparam mult_967_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_967_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_967_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_967_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_967_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_967_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_967_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_967_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_967_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_967_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_967_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_967_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_967_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_967_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_967_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_967_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_967_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_967_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_967_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_967_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_967_mult_2.GSR = "DISABLED";
    defparam mult_967_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_967_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_967_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_967_mult_2.RESETMODE = "SYNC";
    LUT4 i12829_4_lut_4_lut (.A(op_r_23__N_1106[5]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[13] ), .Z(\radix_no1_op_r[5] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12829_4_lut_4_lut.init = 16'h2c20;
    ALU54B lat_alu_29 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n15158), .SIGNEDIB(n15231), .SIGNEDCIN(n15304), .A35(n15157), 
           .A34(n15156), .A33(n15155), .A32(n15154), .A31(n15153), .A30(n15152), 
           .A29(n15151), .A28(n15150), .A27(n15149), .A26(n15148), .A25(n15147), 
           .A24(n15146), .A23(n15145), .A22(n15144), .A21(n15143), .A20(n15142), 
           .A19(n15141), .A18(n15140), .A17(n15139), .A16(n15138), .A15(n15137), 
           .A14(n15136), .A13(n15135), .A12(n15134), .A11(n15133), .A10(n15132), 
           .A9(n15131), .A8(n15130), .A7(n15129), .A6(n15128), .A5(n15127), 
           .A4(n15126), .A3(n15125), .A2(n15124), .A1(n15123), .A0(n15122), 
           .B35(n15230), .B34(n15229), .B33(n15228), .B32(n15227), .B31(n15226), 
           .B30(n15225), .B29(n15224), .B28(n15223), .B27(n15222), .B26(n15221), 
           .B25(n15220), .B24(n15219), .B23(n15218), .B22(n15217), .B21(n15216), 
           .B20(n15215), .B19(n15214), .B18(n15213), .B17(n15212), .B16(n15211), 
           .B15(n15210), .B14(n15209), .B13(n15208), .B12(n15207), .B11(n15206), 
           .B10(n15205), .B9(n15204), .B8(n15203), .B7(n15202), .B6(n15201), 
           .B5(n15200), .B4(n15199), .B3(n15198), .B2(n15197), .B1(n15196), 
           .B0(n15195), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n15194), .MA34(n15193), .MA33(n15192), .MA32(n15191), 
           .MA31(n15190), .MA30(n15189), .MA29(n15188), .MA28(n15187), 
           .MA27(n15186), .MA26(n15185), .MA25(n15184), .MA24(n15183), 
           .MA23(n15182), .MA22(n15181), .MA21(n15180), .MA20(n15179), 
           .MA19(n15178), .MA18(n15177), .MA17(n15176), .MA16(n15175), 
           .MA15(n15174), .MA14(n15173), .MA13(n15172), .MA12(n15171), 
           .MA11(n15170), .MA10(n15169), .MA9(n15168), .MA8(n15167), 
           .MA7(n15166), .MA6(n15165), .MA5(n15164), .MA4(n15163), .MA3(n15162), 
           .MA2(n15161), .MA1(n15160), .MA0(n15159), .MB35(n15267), 
           .MB34(n15266), .MB33(n15265), .MB32(n15264), .MB31(n15263), 
           .MB30(n15262), .MB29(n15261), .MB28(n15260), .MB27(n15259), 
           .MB26(n15258), .MB25(n15257), .MB24(n15256), .MB23(n15255), 
           .MB22(n15254), .MB21(n15253), .MB20(n15252), .MB19(n15251), 
           .MB18(n15250), .MB17(n15249), .MB16(n15248), .MB15(n15247), 
           .MB14(n15246), .MB13(n15245), .MB12(n15244), .MB11(n15243), 
           .MB10(n15242), .MB9(n15241), .MB8(n15240), .MB7(n15239), 
           .MB6(n15238), .MB5(n15237), .MB4(n15236), .MB3(n15235), .MB2(n15234), 
           .MB1(n15233), .MB0(n15232), .CIN53(n15303), .CIN52(n15302), 
           .CIN51(n15301), .CIN50(n15300), .CIN49(n15299), .CIN48(n15298), 
           .CIN47(n15297), .CIN46(n15296), .CIN45(n15295), .CIN44(n15294), 
           .CIN43(n15293), .CIN42(n15292), .CIN41(n15291), .CIN40(n15290), 
           .CIN39(n15289), .CIN38(n15288), .CIN37(n15287), .CIN36(n15286), 
           .CIN35(n15285), .CIN34(n15284), .CIN33(n15283), .CIN32(n15282), 
           .CIN31(n15281), .CIN30(n15280), .CIN29(n15279), .CIN28(n15278), 
           .CIN27(n15277), .CIN26(n15276), .CIN25(n15275), .CIN24(n15274), 
           .CIN23(n15273), .CIN22(n15272), .CIN21(n15271), .CIN20(n15270), 
           .CIN19(n15269), .CIN18(n15268), .CIN17(\op_r_23__N_1226[17] ), 
           .CIN16(\op_r_23__N_1226[16] ), .CIN15(\op_r_23__N_1226[15] ), 
           .CIN14(\op_r_23__N_1226[14] ), .CIN13(\op_r_23__N_1226[13] ), 
           .CIN12(\op_r_23__N_1226[12] ), .CIN11(\op_r_23__N_1226[11] ), 
           .CIN10(\op_r_23__N_1226[10] ), .CIN9(\op_r_23__N_1226[9] ), .CIN8(\op_r_23__N_1226[8] ), 
           .CIN7(\op_r_23__N_1226[7] ), .CIN6(\op_r_23__N_1226[6] ), .CIN5(\op_r_23__N_1226[5] ), 
           .CIN4(\op_r_23__N_1226[4] ), .CIN3(\op_r_23__N_1226[3] ), .CIN2(\op_r_23__N_1226[2] ), 
           .CIN1(\op_r_23__N_1226[1] ), .CIN0(\op_r_23__N_1226[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1226[31] ), 
           .R12(\op_r_23__N_1226[30] ), .R11(\op_r_23__N_1226[29] ), .R10(\op_r_23__N_1226[28] ), 
           .R9(\op_r_23__N_1226[27] ), .R8(\op_r_23__N_1226[26] ), .R7(\op_r_23__N_1226[25] ), 
           .R6(\op_r_23__N_1226[24] ), .R5(\op_r_23__N_1226[23] ), .R4(\op_r_23__N_1226[22] ), 
           .R3(\op_r_23__N_1226[21] ), .R2(\op_r_23__N_1226[20] ), .R1(\op_r_23__N_1226[19] ), 
           .R0(\op_r_23__N_1226[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_29.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_29.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_29.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_29.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_29.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_29.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_29.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_29.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_29.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_29.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_29.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_29.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_29.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_29.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_29.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_29.REG_FLAG_CLK = "NONE";
    defparam lat_alu_29.REG_FLAG_CE = "CE0";
    defparam lat_alu_29.REG_FLAG_RST = "RST0";
    defparam lat_alu_29.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_29.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_29.MASK01 = "0x00000000000000";
    defparam lat_alu_29.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_29.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_29.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_29.CLK0_DIV = "ENABLED";
    defparam lat_alu_29.CLK1_DIV = "ENABLED";
    defparam lat_alu_29.CLK2_DIV = "ENABLED";
    defparam lat_alu_29.CLK3_DIV = "ENABLED";
    defparam lat_alu_29.MCPAT = "0x00000000000000";
    defparam lat_alu_29.MASKPAT = "0x00000000000000";
    defparam lat_alu_29.RNDPAT = "0x00000000000000";
    defparam lat_alu_29.GSR = "DISABLED";
    defparam lat_alu_29.RESETMODE = "SYNC";
    defparam lat_alu_29.MULT9_MODE = "DISABLED";
    defparam lat_alu_29.LEGACY = "DISABLED";
    ALU54B lat_alu_28 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n15012), .SIGNEDIB(n15085), .SIGNEDCIN(GND_net), 
           .A35(n15011), .A34(n15010), .A33(n15009), .A32(n15008), .A31(n15007), 
           .A30(n15006), .A29(n15005), .A28(n15004), .A27(n15003), .A26(n15002), 
           .A25(n15001), .A24(n15000), .A23(n14999), .A22(n14998), .A21(n14997), 
           .A20(n14996), .A19(n14995), .A18(n14994), .A17(n14993), .A16(n14992), 
           .A15(n14991), .A14(n14990), .A13(n14989), .A12(n14988), .A11(n14987), 
           .A10(n14986), .A9(n14985), .A8(n14984), .A7(n14983), .A6(n14982), 
           .A5(n14981), .A4(n14980), .A3(n14979), .A2(n14978), .A1(n14977), 
           .A0(n14976), .B35(n15084), .B34(n15083), .B33(n15082), .B32(n15081), 
           .B31(n15080), .B30(n15079), .B29(n15078), .B28(n15077), .B27(n15076), 
           .B26(n15075), .B25(n15074), .B24(n15073), .B23(n15072), .B22(n15071), 
           .B21(n15070), .B20(n15069), .B19(n15068), .B18(n15067), .B17(n15066), 
           .B16(n15065), .B15(n15064), .B14(n15063), .B13(n15062), .B12(n15061), 
           .B11(n15060), .B10(n15059), .B9(n15058), .B8(n15057), .B7(n15056), 
           .B6(n15055), .B5(n15054), .B4(n15053), .B3(n15052), .B2(n15051), 
           .B1(n15050), .B0(n15049), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n15048), .MA34(n15047), .MA33(n15046), .MA32(n15045), 
           .MA31(n15044), .MA30(n15043), .MA29(n15042), .MA28(n15041), 
           .MA27(n15040), .MA26(n15039), .MA25(n15038), .MA24(n15037), 
           .MA23(n15036), .MA22(n15035), .MA21(n15034), .MA20(n15033), 
           .MA19(n15032), .MA18(n15031), .MA17(n15030), .MA16(n15029), 
           .MA15(n15028), .MA14(n15027), .MA13(n15026), .MA12(n15025), 
           .MA11(n15024), .MA10(n15023), .MA9(n15022), .MA8(n15021), 
           .MA7(n15020), .MA6(n15019), .MA5(n15018), .MA4(n15017), .MA3(n15016), 
           .MA2(n15015), .MA1(n15014), .MA0(n15013), .MB35(n15121), 
           .MB34(n15120), .MB33(n15119), .MB32(n15118), .MB31(n15117), 
           .MB30(n15116), .MB29(n15115), .MB28(n15114), .MB27(n15113), 
           .MB26(n15112), .MB25(n15111), .MB24(n15110), .MB23(n15109), 
           .MB22(n15108), .MB21(n15107), .MB20(n15106), .MB19(n15105), 
           .MB18(n15104), .MB17(n15103), .MB16(n15102), .MB15(n15101), 
           .MB14(n15100), .MB13(n15099), .MB12(n15098), .MB11(n15097), 
           .MB10(n15096), .MB9(n15095), .MB8(n15094), .MB7(n15093), 
           .MB6(n15092), .MB5(n15091), .MB4(n15090), .MB3(n15089), .MB2(n15088), 
           .MB1(n15087), .MB0(n15086), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n15303), 
           .R52(n15302), .R51(n15301), .R50(n15300), .R49(n15299), .R48(n15298), 
           .R47(n15297), .R46(n15296), .R45(n15295), .R44(n15294), .R43(n15293), 
           .R42(n15292), .R41(n15291), .R40(n15290), .R39(n15289), .R38(n15288), 
           .R37(n15287), .R36(n15286), .R35(n15285), .R34(n15284), .R33(n15283), 
           .R32(n15282), .R31(n15281), .R30(n15280), .R29(n15279), .R28(n15278), 
           .R27(n15277), .R26(n15276), .R25(n15275), .R24(n15274), .R23(n15273), 
           .R22(n15272), .R21(n15271), .R20(n15270), .R19(n15269), .R18(n15268), 
           .R17(\op_r_23__N_1226[17] ), .R16(\op_r_23__N_1226[16] ), .R15(\op_r_23__N_1226[15] ), 
           .R14(\op_r_23__N_1226[14] ), .R13(\op_r_23__N_1226[13] ), .R12(\op_r_23__N_1226[12] ), 
           .R11(\op_r_23__N_1226[11] ), .R10(\op_r_23__N_1226[10] ), .R9(\op_r_23__N_1226[9] ), 
           .R8(\op_r_23__N_1226[8] ), .R7(\op_r_23__N_1226[7] ), .R6(\op_r_23__N_1226[6] ), 
           .R5(\op_r_23__N_1226[5] ), .R4(\op_r_23__N_1226[4] ), .R3(\op_r_23__N_1226[3] ), 
           .R2(\op_r_23__N_1226[2] ), .R1(\op_r_23__N_1226[1] ), .R0(\op_r_23__N_1226[0] ), 
           .SIGNEDR(n15304));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_28.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_28.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_28.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_28.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_28.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_28.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_28.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_28.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_28.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_28.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_28.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_28.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_28.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_28.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_28.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_28.REG_FLAG_CLK = "NONE";
    defparam lat_alu_28.REG_FLAG_CE = "CE0";
    defparam lat_alu_28.REG_FLAG_RST = "RST0";
    defparam lat_alu_28.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_28.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_28.MASK01 = "0x00000000000000";
    defparam lat_alu_28.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_28.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_28.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_28.CLK0_DIV = "ENABLED";
    defparam lat_alu_28.CLK1_DIV = "ENABLED";
    defparam lat_alu_28.CLK2_DIV = "ENABLED";
    defparam lat_alu_28.CLK3_DIV = "ENABLED";
    defparam lat_alu_28.MCPAT = "0x00000000000000";
    defparam lat_alu_28.MASKPAT = "0x00000000000000";
    defparam lat_alu_28.RNDPAT = "0x00000000000000";
    defparam lat_alu_28.GSR = "DISABLED";
    defparam lat_alu_28.RESETMODE = "SYNC";
    defparam lat_alu_28.MULT9_MODE = "DISABLED";
    defparam lat_alu_28.LEGACY = "DISABLED";
    LUT4 i12830_4_lut_4_lut (.A(op_r_23__N_1106[6]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[14] ), .Z(\radix_no1_op_r[6] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12830_4_lut_4_lut.init = 16'h2c20;
    ALU54B lat_alu_74 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18272), .SIGNEDIB(n18345), .SIGNEDCIN(n18418), .A35(n18271), 
           .A34(n18270), .A33(n18269), .A32(n18268), .A31(n18267), .A30(n18266), 
           .A29(n18265), .A28(n18264), .A27(n18263), .A26(n18262), .A25(n18261), 
           .A24(n18260), .A23(n18259), .A22(n18258), .A21(n18257), .A20(n18256), 
           .A19(n18255), .A18(n18254), .A17(n18253), .A16(n18252), .A15(n18251), 
           .A14(n18250), .A13(n18249), .A12(n18248), .A11(n18247), .A10(n18246), 
           .A9(n18245), .A8(n18244), .A7(n18243), .A6(n18242), .A5(n18241), 
           .A4(n18240), .A3(n18239), .A2(n18238), .A1(n18237), .A0(n18236), 
           .B35(n18344), .B34(n18343), .B33(n18342), .B32(n18341), .B31(n18340), 
           .B30(n18339), .B29(n18338), .B28(n18337), .B27(n18336), .B26(n18335), 
           .B25(n18334), .B24(n18333), .B23(n18332), .B22(n18331), .B21(n18330), 
           .B20(n18329), .B19(n18328), .B18(n18327), .B17(n18326), .B16(n18325), 
           .B15(n18324), .B14(n18323), .B13(n18322), .B12(n18321), .B11(n18320), 
           .B10(n18319), .B9(n18318), .B8(n18317), .B7(n18316), .B6(n18315), 
           .B5(n18314), .B4(n18313), .B3(n18312), .B2(n18311), .B1(n18310), 
           .B0(n18309), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18308), .MA34(n18307), .MA33(n18306), .MA32(n18305), 
           .MA31(n18304), .MA30(n18303), .MA29(n18302), .MA28(n18301), 
           .MA27(n18300), .MA26(n18299), .MA25(n18298), .MA24(n18297), 
           .MA23(n18296), .MA22(n18295), .MA21(n18294), .MA20(n18293), 
           .MA19(n18292), .MA18(n18291), .MA17(n18290), .MA16(n18289), 
           .MA15(n18288), .MA14(n18287), .MA13(n18286), .MA12(n18285), 
           .MA11(n18284), .MA10(n18283), .MA9(n18282), .MA8(n18281), 
           .MA7(n18280), .MA6(n18279), .MA5(n18278), .MA4(n18277), .MA3(n18276), 
           .MA2(n18275), .MA1(n18274), .MA0(n18273), .MB35(n18381), 
           .MB34(n18380), .MB33(n18379), .MB32(n18378), .MB31(n18377), 
           .MB30(n18376), .MB29(n18375), .MB28(n18374), .MB27(n18373), 
           .MB26(n18372), .MB25(n18371), .MB24(n18370), .MB23(n18369), 
           .MB22(n18368), .MB21(n18367), .MB20(n18366), .MB19(n18365), 
           .MB18(n18364), .MB17(n18363), .MB16(n18362), .MB15(n18361), 
           .MB14(n18360), .MB13(n18359), .MB12(n18358), .MB11(n18357), 
           .MB10(n18356), .MB9(n18355), .MB8(n18354), .MB7(n18353), 
           .MB6(n18352), .MB5(n18351), .MB4(n18350), .MB3(n18349), .MB2(n18348), 
           .MB1(n18347), .MB0(n18346), .CIN53(n18417), .CIN52(n18416), 
           .CIN51(n18415), .CIN50(n18414), .CIN49(n18413), .CIN48(n18412), 
           .CIN47(n18411), .CIN46(n18410), .CIN45(n18409), .CIN44(n18408), 
           .CIN43(n18407), .CIN42(n18406), .CIN41(n18405), .CIN40(n18404), 
           .CIN39(n18403), .CIN38(n18402), .CIN37(n18401), .CIN36(n18400), 
           .CIN35(n18399), .CIN34(n18398), .CIN33(n18397), .CIN32(n18396), 
           .CIN31(n18395), .CIN30(n18394), .CIN29(n18393), .CIN28(n18392), 
           .CIN27(n18391), .CIN26(n18390), .CIN25(n18389), .CIN24(n18388), 
           .CIN23(n18387), .CIN22(n18386), .CIN21(n18385), .CIN20(n18384), 
           .CIN19(n18383), .CIN18(n18382), .CIN17(\op_r_23__N_1268[17] ), 
           .CIN16(\op_r_23__N_1268[16] ), .CIN15(\op_r_23__N_1268[15] ), 
           .CIN14(\op_r_23__N_1268[14] ), .CIN13(\op_r_23__N_1268[13] ), 
           .CIN12(\op_r_23__N_1268[12] ), .CIN11(\op_r_23__N_1268[11] ), 
           .CIN10(\op_r_23__N_1268[10] ), .CIN9(\op_r_23__N_1268[9] ), .CIN8(\op_r_23__N_1268[8] ), 
           .CIN7(\op_r_23__N_1268[7] ), .CIN6(\op_r_23__N_1268[6] ), .CIN5(\op_r_23__N_1268[5] ), 
           .CIN4(\op_r_23__N_1268[4] ), .CIN3(\op_r_23__N_1268[3] ), .CIN2(\op_r_23__N_1268[2] ), 
           .CIN1(\op_r_23__N_1268[1] ), .CIN0(\op_r_23__N_1268[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1268[31] ), 
           .R12(\op_r_23__N_1268[30] ), .R11(\op_r_23__N_1268[29] ), .R10(\op_r_23__N_1268[28] ), 
           .R9(\op_r_23__N_1268[27] ), .R8(\op_r_23__N_1268[26] ), .R7(\op_r_23__N_1268[25] ), 
           .R6(\op_r_23__N_1268[24] ), .R5(\op_r_23__N_1268[23] ), .R4(\op_r_23__N_1268[22] ), 
           .R3(\op_r_23__N_1268[21] ), .R2(\op_r_23__N_1268[20] ), .R1(\op_r_23__N_1268[19] ), 
           .R0(\op_r_23__N_1268[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_74.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_74.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_74.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_74.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_74.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_74.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_74.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_74.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_74.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_74.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_74.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_74.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_74.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_74.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_74.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_74.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_74.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_74.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_74.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_74.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_74.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_74.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_74.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_74.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_74.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_74.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_74.REG_FLAG_CLK = "NONE";
    defparam lat_alu_74.REG_FLAG_CE = "CE0";
    defparam lat_alu_74.REG_FLAG_RST = "RST0";
    defparam lat_alu_74.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_74.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_74.MASK01 = "0x00000000000000";
    defparam lat_alu_74.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_74.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_74.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_74.CLK0_DIV = "ENABLED";
    defparam lat_alu_74.CLK1_DIV = "ENABLED";
    defparam lat_alu_74.CLK2_DIV = "ENABLED";
    defparam lat_alu_74.CLK3_DIV = "ENABLED";
    defparam lat_alu_74.MCPAT = "0x00000000000000";
    defparam lat_alu_74.MASKPAT = "0x00000000000000";
    defparam lat_alu_74.RNDPAT = "0x00000000000000";
    defparam lat_alu_74.GSR = "DISABLED";
    defparam lat_alu_74.RESETMODE = "SYNC";
    defparam lat_alu_74.MULT9_MODE = "DISABLED";
    defparam lat_alu_74.LEGACY = "DISABLED";
    MULT18X18D lat_mult_27 (.A17(\rom16_w_r[9] ), .A16(\rom16_w_r[9] ), 
            .A15(\rom16_w_r[9] ), .A14(\rom16_w_r[9] ), .A13(\rom16_w_r[9] ), 
            .A12(\rom16_w_r[9] ), .A11(\rom16_w_r[9] ), .A10(\rom16_w_r[9] ), 
            .A9(\rom16_w_r[9] ), .A8(\rom16_w_r[9] ), .A7(\rom16_w_r[9] ), 
            .A6(\rom16_w_r[9] ), .A5(\rom16_w_r[9] ), .A4(\rom16_w_r[9] ), 
            .A3(\rom16_w_r[9] ), .A2(\rom16_w_r[9] ), .A1(\rom16_w_r[9] ), 
            .A0(\rom16_w_r[9] ), .B17(n12338), .B16(n12338), .B15(n12338), 
            .B14(n12338), .B13(n12338), .B12(n12338), .B11(n12338), 
            .B10(n12338), .B9(n12338), .B8(n12338), .B7(n12338), .B6(n12338), 
            .B5(n12337), .B4(n12336), .B3(n12335), .B2(n12334), .B1(n12333), 
            .B0(n12332), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n15212), 
            .ROA16(n15211), .ROA15(n15210), .ROA14(n15209), .ROA13(n15208), 
            .ROA12(n15207), .ROA11(n15206), .ROA10(n15205), .ROA9(n15204), 
            .ROA8(n15203), .ROA7(n15202), .ROA6(n15201), .ROA5(n15200), 
            .ROA4(n15199), .ROA3(n15198), .ROA2(n15197), .ROA1(n15196), 
            .ROA0(n15195), .ROB17(n15230), .ROB16(n15229), .ROB15(n15228), 
            .ROB14(n15227), .ROB13(n15226), .ROB12(n15225), .ROB11(n15224), 
            .ROB10(n15223), .ROB9(n15222), .ROB8(n15221), .ROB7(n15220), 
            .ROB6(n15219), .ROB5(n15218), .ROB4(n15217), .ROB3(n15216), 
            .ROB2(n15215), .ROB1(n15214), .ROB0(n15213), .P35(n15267), 
            .P34(n15266), .P33(n15265), .P32(n15264), .P31(n15263), 
            .P30(n15262), .P29(n15261), .P28(n15260), .P27(n15259), 
            .P26(n15258), .P25(n15257), .P24(n15256), .P23(n15255), 
            .P22(n15254), .P21(n15253), .P20(n15252), .P19(n15251), 
            .P18(n15250), .P17(n15249), .P16(n15248), .P15(n15247), 
            .P14(n15246), .P13(n15245), .P12(n15244), .P11(n15243), 
            .P10(n15242), .P9(n15241), .P8(n15240), .P7(n15239), .P6(n15238), 
            .P5(n15237), .P4(n15236), .P3(n15235), .P2(n15234), .P1(n15233), 
            .P0(n15232), .SIGNEDP(n15231));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_27.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_27.REG_INPUTA_CE = "CE0";
    defparam lat_mult_27.REG_INPUTA_RST = "RST0";
    defparam lat_mult_27.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_27.REG_INPUTB_CE = "CE0";
    defparam lat_mult_27.REG_INPUTB_RST = "RST0";
    defparam lat_mult_27.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_27.REG_INPUTC_CE = "CE0";
    defparam lat_mult_27.REG_INPUTC_RST = "RST0";
    defparam lat_mult_27.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_27.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_27.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_27.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_27.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_27.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_27.CLK0_DIV = "ENABLED";
    defparam lat_mult_27.CLK1_DIV = "ENABLED";
    defparam lat_mult_27.CLK2_DIV = "ENABLED";
    defparam lat_mult_27.CLK3_DIV = "ENABLED";
    defparam lat_mult_27.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_27.GSR = "DISABLED";
    defparam lat_mult_27.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_27.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_27.MULT_BYPASS = "DISABLED";
    defparam lat_mult_27.RESETMODE = "SYNC";
    MULT18X18D lat_mult_26 (.A17(\rom16_w_r[9] ), .A16(\rom16_w_r[9] ), 
            .A15(\rom16_w_r[9] ), .A14(\rom16_w_r[9] ), .A13(\rom16_w_r[9] ), 
            .A12(\rom16_w_r[9] ), .A11(\rom16_w_r[9] ), .A10(\rom16_w_r[9] ), 
            .A9(\rom16_w_r[9] ), .A8(\rom16_w_r[8] ), .A7(\rom16_w_r[7] ), 
            .A6(\rom16_w_r[6] ), .A5(\rom16_w_r[5] ), .A4(\rom16_w_r[4] ), 
            .A3(\rom16_w_r[3] ), .A2(\rom16_w_r[2] ), .A1(\rom16_w_r[1] ), 
            .A0(\rom16_w_r[0] ), .B17(n12338), .B16(n12338), .B15(n12338), 
            .B14(n12338), .B13(n12338), .B12(n12338), .B11(n12338), 
            .B10(n12338), .B9(n12338), .B8(n12338), .B7(n12338), .B6(n12338), 
            .B5(n12337), .B4(n12336), .B3(n12335), .B2(n12334), .B1(n12333), 
            .B0(n12332), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n15139), 
            .ROA16(n15138), .ROA15(n15137), .ROA14(n15136), .ROA13(n15135), 
            .ROA12(n15134), .ROA11(n15133), .ROA10(n15132), .ROA9(n15131), 
            .ROA8(n15130), .ROA7(n15129), .ROA6(n15128), .ROA5(n15127), 
            .ROA4(n15126), .ROA3(n15125), .ROA2(n15124), .ROA1(n15123), 
            .ROA0(n15122), .ROB17(n15157), .ROB16(n15156), .ROB15(n15155), 
            .ROB14(n15154), .ROB13(n15153), .ROB12(n15152), .ROB11(n15151), 
            .ROB10(n15150), .ROB9(n15149), .ROB8(n15148), .ROB7(n15147), 
            .ROB6(n15146), .ROB5(n15145), .ROB4(n15144), .ROB3(n15143), 
            .ROB2(n15142), .ROB1(n15141), .ROB0(n15140), .P35(n15194), 
            .P34(n15193), .P33(n15192), .P32(n15191), .P31(n15190), 
            .P30(n15189), .P29(n15188), .P28(n15187), .P27(n15186), 
            .P26(n15185), .P25(n15184), .P24(n15183), .P23(n15182), 
            .P22(n15181), .P21(n15180), .P20(n15179), .P19(n15178), 
            .P18(n15177), .P17(n15176), .P16(n15175), .P15(n15174), 
            .P14(n15173), .P13(n15172), .P12(n15171), .P11(n15170), 
            .P10(n15169), .P9(n15168), .P8(n15167), .P7(n15166), .P6(n15165), 
            .P5(n15164), .P4(n15163), .P3(n15162), .P2(n15161), .P1(n15160), 
            .P0(n15159), .SIGNEDP(n15158));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_26.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_26.REG_INPUTA_CE = "CE0";
    defparam lat_mult_26.REG_INPUTA_RST = "RST0";
    defparam lat_mult_26.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_26.REG_INPUTB_CE = "CE0";
    defparam lat_mult_26.REG_INPUTB_RST = "RST0";
    defparam lat_mult_26.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_26.REG_INPUTC_CE = "CE0";
    defparam lat_mult_26.REG_INPUTC_RST = "RST0";
    defparam lat_mult_26.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_26.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_26.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_26.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_26.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_26.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_26.CLK0_DIV = "ENABLED";
    defparam lat_mult_26.CLK1_DIV = "ENABLED";
    defparam lat_mult_26.CLK2_DIV = "ENABLED";
    defparam lat_mult_26.CLK3_DIV = "ENABLED";
    defparam lat_mult_26.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_26.GSR = "DISABLED";
    defparam lat_mult_26.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_26.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_26.MULT_BYPASS = "DISABLED";
    defparam lat_mult_26.RESETMODE = "SYNC";
    MULT18X18D lat_mult_25 (.A17(\rom16_w_r[9] ), .A16(\rom16_w_r[9] ), 
            .A15(\rom16_w_r[9] ), .A14(\rom16_w_r[9] ), .A13(\rom16_w_r[9] ), 
            .A12(\rom16_w_r[9] ), .A11(\rom16_w_r[9] ), .A10(\rom16_w_r[9] ), 
            .A9(\rom16_w_r[9] ), .A8(\rom16_w_r[9] ), .A7(\rom16_w_r[9] ), 
            .A6(\rom16_w_r[9] ), .A5(\rom16_w_r[9] ), .A4(\rom16_w_r[9] ), 
            .A3(\rom16_w_r[9] ), .A2(\rom16_w_r[9] ), .A1(\rom16_w_r[9] ), 
            .A0(\rom16_w_r[9] ), .B17(n12331), .B16(n12330), .B15(n12329), 
            .B14(n12328), .B13(n12327), .B12(n12326), .B11(n12325), 
            .B10(n12324), .B9(n12323), .B8(n12322), .B7(n12321), .B6(n12320), 
            .B5(n12319), .B4(n12318), .B3(n12317), .B2(n12316), .B1(n12315), 
            .B0(n12314), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n15066), 
            .ROA16(n15065), .ROA15(n15064), .ROA14(n15063), .ROA13(n15062), 
            .ROA12(n15061), .ROA11(n15060), .ROA10(n15059), .ROA9(n15058), 
            .ROA8(n15057), .ROA7(n15056), .ROA6(n15055), .ROA5(n15054), 
            .ROA4(n15053), .ROA3(n15052), .ROA2(n15051), .ROA1(n15050), 
            .ROA0(n15049), .ROB17(n15084), .ROB16(n15083), .ROB15(n15082), 
            .ROB14(n15081), .ROB13(n15080), .ROB12(n15079), .ROB11(n15078), 
            .ROB10(n15077), .ROB9(n15076), .ROB8(n15075), .ROB7(n15074), 
            .ROB6(n15073), .ROB5(n15072), .ROB4(n15071), .ROB3(n15070), 
            .ROB2(n15069), .ROB1(n15068), .ROB0(n15067), .P35(n15121), 
            .P34(n15120), .P33(n15119), .P32(n15118), .P31(n15117), 
            .P30(n15116), .P29(n15115), .P28(n15114), .P27(n15113), 
            .P26(n15112), .P25(n15111), .P24(n15110), .P23(n15109), 
            .P22(n15108), .P21(n15107), .P20(n15106), .P19(n15105), 
            .P18(n15104), .P17(n15103), .P16(n15102), .P15(n15101), 
            .P14(n15100), .P13(n15099), .P12(n15098), .P11(n15097), 
            .P10(n15096), .P9(n15095), .P8(n15094), .P7(n15093), .P6(n15092), 
            .P5(n15091), .P4(n15090), .P3(n15089), .P2(n15088), .P1(n15087), 
            .P0(n15086), .SIGNEDP(n15085));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_25.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_25.REG_INPUTA_CE = "CE0";
    defparam lat_mult_25.REG_INPUTA_RST = "RST0";
    defparam lat_mult_25.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_25.REG_INPUTB_CE = "CE0";
    defparam lat_mult_25.REG_INPUTB_RST = "RST0";
    defparam lat_mult_25.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_25.REG_INPUTC_CE = "CE0";
    defparam lat_mult_25.REG_INPUTC_RST = "RST0";
    defparam lat_mult_25.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_25.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_25.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_25.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_25.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_25.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_25.CLK0_DIV = "ENABLED";
    defparam lat_mult_25.CLK1_DIV = "ENABLED";
    defparam lat_mult_25.CLK2_DIV = "ENABLED";
    defparam lat_mult_25.CLK3_DIV = "ENABLED";
    defparam lat_mult_25.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_25.GSR = "DISABLED";
    defparam lat_mult_25.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_25.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_25.MULT_BYPASS = "DISABLED";
    defparam lat_mult_25.RESETMODE = "SYNC";
    LUT4 i12831_4_lut_4_lut (.A(op_r_23__N_1106[7]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_r_23__N_1082[15] ), .Z(\radix_no1_op_r[7] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12831_4_lut_4_lut.init = 16'h2c20;
    MULT18X18D mult_10_mult_2 (.A17(\rom16_w_r[9] ), .A16(\rom16_w_r[9] ), 
            .A15(\rom16_w_r[9] ), .A14(\rom16_w_r[9] ), .A13(\rom16_w_r[9] ), 
            .A12(\rom16_w_r[9] ), .A11(\rom16_w_r[9] ), .A10(\rom16_w_r[9] ), 
            .A9(\rom16_w_r[9] ), .A8(\rom16_w_r[8] ), .A7(\rom16_w_r[7] ), 
            .A6(\rom16_w_r[6] ), .A5(\rom16_w_r[5] ), .A4(\rom16_w_r[4] ), 
            .A3(\rom16_w_r[3] ), .A2(\rom16_w_r[2] ), .A1(\rom16_w_r[1] ), 
            .A0(\rom16_w_r[0] ), .B17(n12331), .B16(n12330), .B15(n12329), 
            .B14(n12328), .B13(n12327), .B12(n12326), .B11(n12325), 
            .B10(n12324), .B9(n12323), .B8(n12322), .B7(n12321), .B6(n12320), 
            .B5(n12319), .B4(n12318), .B3(n12317), .B2(n12316), .B1(n12315), 
            .B0(n12314), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14993), 
            .ROA16(n14992), .ROA15(n14991), .ROA14(n14990), .ROA13(n14989), 
            .ROA12(n14988), .ROA11(n14987), .ROA10(n14986), .ROA9(n14985), 
            .ROA8(n14984), .ROA7(n14983), .ROA6(n14982), .ROA5(n14981), 
            .ROA4(n14980), .ROA3(n14979), .ROA2(n14978), .ROA1(n14977), 
            .ROA0(n14976), .ROB17(n15011), .ROB16(n15010), .ROB15(n15009), 
            .ROB14(n15008), .ROB13(n15007), .ROB12(n15006), .ROB11(n15005), 
            .ROB10(n15004), .ROB9(n15003), .ROB8(n15002), .ROB7(n15001), 
            .ROB6(n15000), .ROB5(n14999), .ROB4(n14998), .ROB3(n14997), 
            .ROB2(n14996), .ROB1(n14995), .ROB0(n14994), .P35(n15048), 
            .P34(n15047), .P33(n15046), .P32(n15045), .P31(n15044), 
            .P30(n15043), .P29(n15042), .P28(n15041), .P27(n15040), 
            .P26(n15039), .P25(n15038), .P24(n15037), .P23(n15036), 
            .P22(n15035), .P21(n15034), .P20(n15033), .P19(n15032), 
            .P18(n15031), .P17(n15030), .P16(n15029), .P15(n15028), 
            .P14(n15027), .P13(n15026), .P12(n15025), .P11(n15024), 
            .P10(n15023), .P9(n15022), .P8(n15021), .P7(n15020), .P6(n15019), 
            .P5(n15018), .P4(n15017), .P3(n15016), .P2(n15015), .P1(n15014), 
            .P0(n15013), .SIGNEDP(n15012));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam mult_10_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_10_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_10_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_10_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_10_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_10_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_10_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_10_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_10_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_10_mult_2.GSR = "DISABLED";
    defparam mult_10_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_10_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_10_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_10_mult_2.RESETMODE = "SYNC";
    LUT4 i12549_4_lut_4_lut (.A(op_i_23__N_1154[0]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[8] ), .Z(\radix_no1_op_i[0] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12549_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12848_4_lut_4_lut (.A(op_i_23__N_1154[1]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[9] ), .Z(\radix_no1_op_i[1] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12848_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12849_4_lut_4_lut (.A(op_i_23__N_1154[2]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[10] ), .Z(\radix_no1_op_i[2] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12849_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12850_4_lut_4_lut (.A(op_i_23__N_1154[3]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[11] ), .Z(\radix_no1_op_i[3] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12850_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12851_4_lut_4_lut (.A(op_i_23__N_1154[4]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[12] ), .Z(\radix_no1_op_i[4] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12851_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12852_4_lut_4_lut (.A(op_i_23__N_1154[5]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[13] ), .Z(\radix_no1_op_i[5] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12852_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12853_4_lut_4_lut (.A(op_i_23__N_1154[6]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[14] ), .Z(\radix_no1_op_i[6] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12853_4_lut_4_lut.init = 16'h2c20;
    LUT4 i12854_4_lut_4_lut (.A(op_i_23__N_1154[7]), .B(\count[5] ), .C(\count[4] ), 
         .D(\op_i_23__N_1130[15] ), .Z(\radix_no1_op_i[7] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12854_4_lut_4_lut.init = 16'h2c20;
    ALU54B lat_alu_4 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n13360), .SIGNEDIB(n13433), .SIGNEDCIN(n13506), .A35(n13359), 
           .A34(n13358), .A33(n13357), .A32(n13356), .A31(n13355), .A30(n13354), 
           .A29(n13353), .A28(n13352), .A27(n13351), .A26(n13350), .A25(n13349), 
           .A24(n13348), .A23(n13347), .A22(n13346), .A21(n13345), .A20(n13344), 
           .A19(n13343), .A18(n13342), .A17(n13341), .A16(n13340), .A15(n13339), 
           .A14(n13338), .A13(n13337), .A12(n13336), .A11(n13335), .A10(n13334), 
           .A9(n13333), .A8(n13332), .A7(n13331), .A6(n13330), .A5(n13329), 
           .A4(n13328), .A3(n13327), .A2(n13326), .A1(n13325), .A0(n13324), 
           .B35(n13432), .B34(n13431), .B33(n13430), .B32(n13429), .B31(n13428), 
           .B30(n13427), .B29(n13426), .B28(n13425), .B27(n13424), .B26(n13423), 
           .B25(n13422), .B24(n13421), .B23(n13420), .B22(n13419), .B21(n13418), 
           .B20(n13417), .B19(n13416), .B18(n13415), .B17(n13414), .B16(n13413), 
           .B15(n13412), .B14(n13411), .B13(n13410), .B12(n13409), .B11(n13408), 
           .B10(n13407), .B9(n13406), .B8(n13405), .B7(n13404), .B6(n13403), 
           .B5(n13402), .B4(n13401), .B3(n13400), .B2(n13399), .B1(n13398), 
           .B0(n13397), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n13396), .MA34(n13395), .MA33(n13394), .MA32(n13393), 
           .MA31(n13392), .MA30(n13391), .MA29(n13390), .MA28(n13389), 
           .MA27(n13388), .MA26(n13387), .MA25(n13386), .MA24(n13385), 
           .MA23(n13384), .MA22(n13383), .MA21(n13382), .MA20(n13381), 
           .MA19(n13380), .MA18(n13379), .MA17(n13378), .MA16(n13377), 
           .MA15(n13376), .MA14(n13375), .MA13(n13374), .MA12(n13373), 
           .MA11(n13372), .MA10(n13371), .MA9(n13370), .MA8(n13369), 
           .MA7(n13368), .MA6(n13367), .MA5(n13366), .MA4(n13365), .MA3(n13364), 
           .MA2(n13363), .MA1(n13362), .MA0(n13361), .MB35(n13469), 
           .MB34(n13468), .MB33(n13467), .MB32(n13466), .MB31(n13465), 
           .MB30(n13464), .MB29(n13463), .MB28(n13462), .MB27(n13461), 
           .MB26(n13460), .MB25(n13459), .MB24(n13458), .MB23(n13457), 
           .MB22(n13456), .MB21(n13455), .MB20(n13454), .MB19(n13453), 
           .MB18(n13452), .MB17(n13451), .MB16(n13450), .MB15(n13449), 
           .MB14(n13448), .MB13(n13447), .MB12(n13446), .MB11(n13445), 
           .MB10(n13444), .MB9(n13443), .MB8(n13442), .MB7(n13441), 
           .MB6(n13440), .MB5(n13439), .MB4(n13438), .MB3(n13437), .MB2(n13436), 
           .MB1(n13435), .MB0(n13434), .CIN53(n13505), .CIN52(n13504), 
           .CIN51(n13503), .CIN50(n13502), .CIN49(n13501), .CIN48(n13500), 
           .CIN47(n13499), .CIN46(n13498), .CIN45(n13497), .CIN44(n13496), 
           .CIN43(n13495), .CIN42(n13494), .CIN41(n13493), .CIN40(n13492), 
           .CIN39(n13491), .CIN38(n13490), .CIN37(n13489), .CIN36(n13488), 
           .CIN35(n13487), .CIN34(n13486), .CIN33(n13485), .CIN32(n13484), 
           .CIN31(n13483), .CIN30(n13482), .CIN29(n13481), .CIN28(n13480), 
           .CIN27(n13479), .CIN26(n13478), .CIN25(n13477), .CIN24(n13476), 
           .CIN23(n13475), .CIN22(n13474), .CIN21(n13473), .CIN20(n13472), 
           .CIN19(n13471), .CIN18(n13470), .CIN17(n8576), .CIN16(n8577), 
           .CIN15(n8578), .CIN14(n8579), .CIN13(n8580), .CIN12(n8581), 
           .CIN11(n8582), .CIN10(n8583), .CIN9(n8584), .CIN8(n8585), 
           .CIN7(n8586), .CIN6(n8587), .CIN5(n8588), .CIN4(n8589), .CIN3(n8590), 
           .CIN2(n8591), .CIN1(n8592), .CIN0(n8593), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R7(n8568), .R6(n8569), .R5(n8570), 
           .R4(n8571), .R3(n8572), .R2(n8573), .R1(n8574), .R0(n8575));
    defparam lat_alu_4.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_4.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_4.REG_FLAG_CLK = "NONE";
    defparam lat_alu_4.REG_FLAG_CE = "CE0";
    defparam lat_alu_4.REG_FLAG_RST = "RST0";
    defparam lat_alu_4.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASK01 = "0x00000000000000";
    defparam lat_alu_4.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_4.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_4.CLK0_DIV = "ENABLED";
    defparam lat_alu_4.CLK1_DIV = "ENABLED";
    defparam lat_alu_4.CLK2_DIV = "ENABLED";
    defparam lat_alu_4.CLK3_DIV = "ENABLED";
    defparam lat_alu_4.MCPAT = "0x00000000000000";
    defparam lat_alu_4.MASKPAT = "0x00000000000000";
    defparam lat_alu_4.RNDPAT = "0x00000000000000";
    defparam lat_alu_4.GSR = "DISABLED";
    defparam lat_alu_4.RESETMODE = "SYNC";
    defparam lat_alu_4.MULT9_MODE = "DISABLED";
    defparam lat_alu_4.LEGACY = "DISABLED";
    ALU54B lat_alu_3 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n13214), .SIGNEDIB(n13287), .SIGNEDCIN(GND_net), 
           .A35(n13213), .A34(n13212), .A33(n13211), .A32(n13210), .A31(n13209), 
           .A30(n13208), .A29(n13207), .A28(n13206), .A27(n13205), .A26(n13204), 
           .A25(n13203), .A24(n13202), .A23(n13201), .A22(n13200), .A21(n13199), 
           .A20(n13198), .A19(n13197), .A18(n13196), .A17(n13195), .A16(n13194), 
           .A15(n13193), .A14(n13192), .A13(n13191), .A12(n13190), .A11(n13189), 
           .A10(n13188), .A9(n13187), .A8(n13186), .A7(n13185), .A6(n13184), 
           .A5(n13183), .A4(n13182), .A3(n13181), .A2(n13180), .A1(n13179), 
           .A0(n13178), .B35(n13286), .B34(n13285), .B33(n13284), .B32(n13283), 
           .B31(n13282), .B30(n13281), .B29(n13280), .B28(n13279), .B27(n13278), 
           .B26(n13277), .B25(n13276), .B24(n13275), .B23(n13274), .B22(n13273), 
           .B21(n13272), .B20(n13271), .B19(n13270), .B18(n13269), .B17(n13268), 
           .B16(n13267), .B15(n13266), .B14(n13265), .B13(n13264), .B12(n13263), 
           .B11(n13262), .B10(n13261), .B9(n13260), .B8(n13259), .B7(n13258), 
           .B6(n13257), .B5(n13256), .B4(n13255), .B3(n13254), .B2(n13253), 
           .B1(n13252), .B0(n13251), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n13250), .MA34(n13249), .MA33(n13248), .MA32(n13247), 
           .MA31(n13246), .MA30(n13245), .MA29(n13244), .MA28(n13243), 
           .MA27(n13242), .MA26(n13241), .MA25(n13240), .MA24(n13239), 
           .MA23(n13238), .MA22(n13237), .MA21(n13236), .MA20(n13235), 
           .MA19(n13234), .MA18(n13233), .MA17(n13232), .MA16(n13231), 
           .MA15(n13230), .MA14(n13229), .MA13(n13228), .MA12(n13227), 
           .MA11(n13226), .MA10(n13225), .MA9(n13224), .MA8(n13223), 
           .MA7(n13222), .MA6(n13221), .MA5(n13220), .MA4(n13219), .MA3(n13218), 
           .MA2(n13217), .MA1(n13216), .MA0(n13215), .MB35(n13323), 
           .MB34(n13322), .MB33(n13321), .MB32(n13320), .MB31(n13319), 
           .MB30(n13318), .MB29(n13317), .MB28(n13316), .MB27(n13315), 
           .MB26(n13314), .MB25(n13313), .MB24(n13312), .MB23(n13311), 
           .MB22(n13310), .MB21(n13309), .MB20(n13308), .MB19(n13307), 
           .MB18(n13306), .MB17(n13305), .MB16(n13304), .MB15(n13303), 
           .MB14(n13302), .MB13(n13301), .MB12(n13300), .MB11(n13299), 
           .MB10(n13298), .MB9(n13297), .MB8(n13296), .MB7(n13295), 
           .MB6(n13294), .MB5(n13293), .MB4(n13292), .MB3(n13291), .MB2(n13290), 
           .MB1(n13289), .MB0(n13288), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n13505), 
           .R52(n13504), .R51(n13503), .R50(n13502), .R49(n13501), .R48(n13500), 
           .R47(n13499), .R46(n13498), .R45(n13497), .R44(n13496), .R43(n13495), 
           .R42(n13494), .R41(n13493), .R40(n13492), .R39(n13491), .R38(n13490), 
           .R37(n13489), .R36(n13488), .R35(n13487), .R34(n13486), .R33(n13485), 
           .R32(n13484), .R31(n13483), .R30(n13482), .R29(n13481), .R28(n13480), 
           .R27(n13479), .R26(n13478), .R25(n13477), .R24(n13476), .R23(n13475), 
           .R22(n13474), .R21(n13473), .R20(n13472), .R19(n13471), .R18(n13470), 
           .R17(n8576), .R16(n8577), .R15(n8578), .R14(n8579), .R13(n8580), 
           .R12(n8581), .R11(n8582), .R10(n8583), .R9(n8584), .R8(n8585), 
           .R7(n8586), .R6(n8587), .R5(n8588), .R4(n8589), .R3(n8590), 
           .R2(n8591), .R1(n8592), .R0(n8593), .SIGNEDR(n13506));
    defparam lat_alu_3.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_3.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_3.REG_FLAG_CLK = "NONE";
    defparam lat_alu_3.REG_FLAG_CE = "CE0";
    defparam lat_alu_3.REG_FLAG_RST = "RST0";
    defparam lat_alu_3.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASK01 = "0x00000000000000";
    defparam lat_alu_3.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_3.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_3.CLK0_DIV = "ENABLED";
    defparam lat_alu_3.CLK1_DIV = "ENABLED";
    defparam lat_alu_3.CLK2_DIV = "ENABLED";
    defparam lat_alu_3.CLK3_DIV = "ENABLED";
    defparam lat_alu_3.MCPAT = "0x00000000000000";
    defparam lat_alu_3.MASKPAT = "0x00000000000000";
    defparam lat_alu_3.RNDPAT = "0x00000000000000";
    defparam lat_alu_3.GSR = "DISABLED";
    defparam lat_alu_3.RESETMODE = "SYNC";
    defparam lat_alu_3.MULT9_MODE = "DISABLED";
    defparam lat_alu_3.LEGACY = "DISABLED";
    MULT18X18D lat_mult_2 (.A17(\rom16_w_i[8] ), .A16(\rom16_w_i[8] ), .A15(\rom16_w_i[8] ), 
            .A14(\rom16_w_i[8] ), .A13(\rom16_w_i[8] ), .A12(\rom16_w_i[8] ), 
            .A11(\rom16_w_i[8] ), .A10(\rom16_w_i[8] ), .A9(\rom16_w_i[8] ), 
            .A8(\rom16_w_i[8] ), .A7(\rom16_w_i[8] ), .A6(\rom16_w_i[8] ), 
            .A5(\rom16_w_i[8] ), .A4(\rom16_w_i[8] ), .A3(\rom16_w_i[8] ), 
            .A2(\rom16_w_i[8] ), .A1(\rom16_w_i[8] ), .A0(\rom16_w_i[8] ), 
            .B17(n319), .B16(n319), .B15(n319), .B14(n319), .B13(n319), 
            .B12(n319), .B11(n319), .B10(n319), .B9(n319), .B8(n319), 
            .B7(n319), .B6(n319), .B5(n319), .B4(n319), .B3(n319), 
            .B2(n319), .B1(n319), .B0(n319), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n13414), .ROA16(n13413), .ROA15(n13412), .ROA14(n13411), 
            .ROA13(n13410), .ROA12(n13409), .ROA11(n13408), .ROA10(n13407), 
            .ROA9(n13406), .ROA8(n13405), .ROA7(n13404), .ROA6(n13403), 
            .ROA5(n13402), .ROA4(n13401), .ROA3(n13400), .ROA2(n13399), 
            .ROA1(n13398), .ROA0(n13397), .ROB17(n13432), .ROB16(n13431), 
            .ROB15(n13430), .ROB14(n13429), .ROB13(n13428), .ROB12(n13427), 
            .ROB11(n13426), .ROB10(n13425), .ROB9(n13424), .ROB8(n13423), 
            .ROB7(n13422), .ROB6(n13421), .ROB5(n13420), .ROB4(n13419), 
            .ROB3(n13418), .ROB2(n13417), .ROB1(n13416), .ROB0(n13415), 
            .P35(n13469), .P34(n13468), .P33(n13467), .P32(n13466), 
            .P31(n13465), .P30(n13464), .P29(n13463), .P28(n13462), 
            .P27(n13461), .P26(n13460), .P25(n13459), .P24(n13458), 
            .P23(n13457), .P22(n13456), .P21(n13455), .P20(n13454), 
            .P19(n13453), .P18(n13452), .P17(n13451), .P16(n13450), 
            .P15(n13449), .P14(n13448), .P13(n13447), .P12(n13446), 
            .P11(n13445), .P10(n13444), .P9(n13443), .P8(n13442), .P7(n13441), 
            .P6(n13440), .P5(n13439), .P4(n13438), .P3(n13437), .P2(n13436), 
            .P1(n13435), .P0(n13434), .SIGNEDP(n13433));
    defparam lat_mult_2.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTA_CE = "CE0";
    defparam lat_mult_2.REG_INPUTA_RST = "RST0";
    defparam lat_mult_2.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTB_CE = "CE0";
    defparam lat_mult_2.REG_INPUTB_RST = "RST0";
    defparam lat_mult_2.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTC_CE = "CE0";
    defparam lat_mult_2.REG_INPUTC_RST = "RST0";
    defparam lat_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_2.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_2.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_2.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_2.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_2.CLK0_DIV = "ENABLED";
    defparam lat_mult_2.CLK1_DIV = "ENABLED";
    defparam lat_mult_2.CLK2_DIV = "ENABLED";
    defparam lat_mult_2.CLK3_DIV = "ENABLED";
    defparam lat_mult_2.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_2.GSR = "DISABLED";
    defparam lat_mult_2.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_2.MULT_BYPASS = "DISABLED";
    defparam lat_mult_2.RESETMODE = "SYNC";
    MULT18X18D lat_mult_1 (.A17(\rom16_w_i[8] ), .A16(\rom16_w_i[8] ), .A15(\rom16_w_i[8] ), 
            .A14(\rom16_w_i[8] ), .A13(\rom16_w_i[8] ), .A12(\rom16_w_i[8] ), 
            .A11(\rom16_w_i[8] ), .A10(\rom16_w_i[8] ), .A9(\rom16_w_i[8] ), 
            .A8(\rom16_w_i[8] ), .A7(\rom16_w_i[7] ), .A6(\rom16_w_i[6] ), 
            .A5(\rom16_w_i[5] ), .A4(\rom16_w_i[4] ), .A3(\rom16_w_i[3] ), 
            .A2(\rom16_w_i[2] ), .A1(\rom16_w_i[1] ), .A0(\rom16_w_i[0] ), 
            .B17(n319), .B16(n319), .B15(n319), .B14(n319), .B13(n319), 
            .B12(n319), .B11(n319), .B10(n319), .B9(n319), .B8(n319), 
            .B7(n319), .B6(n319), .B5(n319), .B4(n319), .B3(n319), 
            .B2(n319), .B1(n319), .B0(n319), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n13341), .ROA16(n13340), .ROA15(n13339), .ROA14(n13338), 
            .ROA13(n13337), .ROA12(n13336), .ROA11(n13335), .ROA10(n13334), 
            .ROA9(n13333), .ROA8(n13332), .ROA7(n13331), .ROA6(n13330), 
            .ROA5(n13329), .ROA4(n13328), .ROA3(n13327), .ROA2(n13326), 
            .ROA1(n13325), .ROA0(n13324), .ROB17(n13359), .ROB16(n13358), 
            .ROB15(n13357), .ROB14(n13356), .ROB13(n13355), .ROB12(n13354), 
            .ROB11(n13353), .ROB10(n13352), .ROB9(n13351), .ROB8(n13350), 
            .ROB7(n13349), .ROB6(n13348), .ROB5(n13347), .ROB4(n13346), 
            .ROB3(n13345), .ROB2(n13344), .ROB1(n13343), .ROB0(n13342), 
            .P35(n13396), .P34(n13395), .P33(n13394), .P32(n13393), 
            .P31(n13392), .P30(n13391), .P29(n13390), .P28(n13389), 
            .P27(n13388), .P26(n13387), .P25(n13386), .P24(n13385), 
            .P23(n13384), .P22(n13383), .P21(n13382), .P20(n13381), 
            .P19(n13380), .P18(n13379), .P17(n13378), .P16(n13377), 
            .P15(n13376), .P14(n13375), .P13(n13374), .P12(n13373), 
            .P11(n13372), .P10(n13371), .P9(n13370), .P8(n13369), .P7(n13368), 
            .P6(n13367), .P5(n13366), .P4(n13365), .P3(n13364), .P2(n13363), 
            .P1(n13362), .P0(n13361), .SIGNEDP(n13360));
    defparam lat_mult_1.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTA_CE = "CE0";
    defparam lat_mult_1.REG_INPUTA_RST = "RST0";
    defparam lat_mult_1.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTB_CE = "CE0";
    defparam lat_mult_1.REG_INPUTB_RST = "RST0";
    defparam lat_mult_1.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTC_CE = "CE0";
    defparam lat_mult_1.REG_INPUTC_RST = "RST0";
    defparam lat_mult_1.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_1.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_1.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_1.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_1.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_1.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_1.CLK0_DIV = "ENABLED";
    defparam lat_mult_1.CLK1_DIV = "ENABLED";
    defparam lat_mult_1.CLK2_DIV = "ENABLED";
    defparam lat_mult_1.CLK3_DIV = "ENABLED";
    defparam lat_mult_1.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_1.GSR = "DISABLED";
    defparam lat_mult_1.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_1.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_1.MULT_BYPASS = "DISABLED";
    defparam lat_mult_1.RESETMODE = "SYNC";
    MULT18X18D lat_mult_0 (.A17(\rom16_w_i[8] ), .A16(\rom16_w_i[8] ), .A15(\rom16_w_i[8] ), 
            .A14(\rom16_w_i[8] ), .A13(\rom16_w_i[8] ), .A12(\rom16_w_i[8] ), 
            .A11(\rom16_w_i[8] ), .A10(\rom16_w_i[8] ), .A9(\rom16_w_i[8] ), 
            .A8(\rom16_w_i[8] ), .A7(\rom16_w_i[8] ), .A6(\rom16_w_i[8] ), 
            .A5(\rom16_w_i[8] ), .A4(\rom16_w_i[8] ), .A3(\rom16_w_i[8] ), 
            .A2(\rom16_w_i[8] ), .A1(\rom16_w_i[8] ), .A0(\rom16_w_i[8] ), 
            .B17(n10006), .B16(n10005), .B15(n10004), .B14(n10003), 
            .B13(n10002), .B12(n10001), .B11(n10000), .B10(n9999), .B9(n9998), 
            .B8(n9997), .B7(n9996), .B6(n9995), .B5(n9994), .B4(n9993), 
            .B3(n9992), .B2(n9991), .B1(n9990), .B0(n9989), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n13268), .ROA16(n13267), .ROA15(n13266), 
            .ROA14(n13265), .ROA13(n13264), .ROA12(n13263), .ROA11(n13262), 
            .ROA10(n13261), .ROA9(n13260), .ROA8(n13259), .ROA7(n13258), 
            .ROA6(n13257), .ROA5(n13256), .ROA4(n13255), .ROA3(n13254), 
            .ROA2(n13253), .ROA1(n13252), .ROA0(n13251), .ROB17(n13286), 
            .ROB16(n13285), .ROB15(n13284), .ROB14(n13283), .ROB13(n13282), 
            .ROB12(n13281), .ROB11(n13280), .ROB10(n13279), .ROB9(n13278), 
            .ROB8(n13277), .ROB7(n13276), .ROB6(n13275), .ROB5(n13274), 
            .ROB4(n13273), .ROB3(n13272), .ROB2(n13271), .ROB1(n13270), 
            .ROB0(n13269), .P35(n13323), .P34(n13322), .P33(n13321), 
            .P32(n13320), .P31(n13319), .P30(n13318), .P29(n13317), 
            .P28(n13316), .P27(n13315), .P26(n13314), .P25(n13313), 
            .P24(n13312), .P23(n13311), .P22(n13310), .P21(n13309), 
            .P20(n13308), .P19(n13307), .P18(n13306), .P17(n13305), 
            .P16(n13304), .P15(n13303), .P14(n13302), .P13(n13301), 
            .P12(n13300), .P11(n13299), .P10(n13298), .P9(n13297), .P8(n13296), 
            .P7(n13295), .P6(n13294), .P5(n13293), .P4(n13292), .P3(n13291), 
            .P2(n13290), .P1(n13289), .P0(n13288), .SIGNEDP(n13287));
    defparam lat_mult_0.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTA_CE = "CE0";
    defparam lat_mult_0.REG_INPUTA_RST = "RST0";
    defparam lat_mult_0.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTB_CE = "CE0";
    defparam lat_mult_0.REG_INPUTB_RST = "RST0";
    defparam lat_mult_0.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTC_CE = "CE0";
    defparam lat_mult_0.REG_INPUTC_RST = "RST0";
    defparam lat_mult_0.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_0.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_0.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_0.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_0.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_0.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_0.CLK0_DIV = "ENABLED";
    defparam lat_mult_0.CLK1_DIV = "ENABLED";
    defparam lat_mult_0.CLK2_DIV = "ENABLED";
    defparam lat_mult_0.CLK3_DIV = "ENABLED";
    defparam lat_mult_0.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_0.GSR = "DISABLED";
    defparam lat_mult_0.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_0.MULT_BYPASS = "DISABLED";
    defparam lat_mult_0.RESETMODE = "SYNC";
    MULT18X18D mult_966 (.A17(\rom16_w_i[8] ), .A16(\rom16_w_i[8] ), .A15(\rom16_w_i[8] ), 
            .A14(\rom16_w_i[8] ), .A13(\rom16_w_i[8] ), .A12(\rom16_w_i[8] ), 
            .A11(\rom16_w_i[8] ), .A10(\rom16_w_i[8] ), .A9(\rom16_w_i[8] ), 
            .A8(\rom16_w_i[8] ), .A7(\rom16_w_i[7] ), .A6(\rom16_w_i[6] ), 
            .A5(\rom16_w_i[5] ), .A4(\rom16_w_i[4] ), .A3(\rom16_w_i[3] ), 
            .A2(\rom16_w_i[2] ), .A1(\rom16_w_i[1] ), .A0(\rom16_w_i[0] ), 
            .B17(n10006), .B16(n10005), .B15(n10004), .B14(n10003), 
            .B13(n10002), .B12(n10001), .B11(n10000), .B10(n9999), .B9(n9998), 
            .B8(n9997), .B7(n9996), .B6(n9995), .B5(n9994), .B4(n9993), 
            .B3(n9992), .B2(n9991), .B1(n9990), .B0(n9989), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n13195), .ROA16(n13194), .ROA15(n13193), 
            .ROA14(n13192), .ROA13(n13191), .ROA12(n13190), .ROA11(n13189), 
            .ROA10(n13188), .ROA9(n13187), .ROA8(n13186), .ROA7(n13185), 
            .ROA6(n13184), .ROA5(n13183), .ROA4(n13182), .ROA3(n13181), 
            .ROA2(n13180), .ROA1(n13179), .ROA0(n13178), .ROB17(n13213), 
            .ROB16(n13212), .ROB15(n13211), .ROB14(n13210), .ROB13(n13209), 
            .ROB12(n13208), .ROB11(n13207), .ROB10(n13206), .ROB9(n13205), 
            .ROB8(n13204), .ROB7(n13203), .ROB6(n13202), .ROB5(n13201), 
            .ROB4(n13200), .ROB3(n13199), .ROB2(n13198), .ROB1(n13197), 
            .ROB0(n13196), .P35(n13250), .P34(n13249), .P33(n13248), 
            .P32(n13247), .P31(n13246), .P30(n13245), .P29(n13244), 
            .P28(n13243), .P27(n13242), .P26(n13241), .P25(n13240), 
            .P24(n13239), .P23(n13238), .P22(n13237), .P21(n13236), 
            .P20(n13235), .P19(n13234), .P18(n13233), .P17(n13232), 
            .P16(n13231), .P15(n13230), .P14(n13229), .P13(n13228), 
            .P12(n13227), .P11(n13226), .P10(n13225), .P9(n13224), .P8(n13223), 
            .P7(n13222), .P6(n13221), .P5(n13220), .P4(n13219), .P3(n13218), 
            .P2(n13217), .P1(n13216), .P0(n13215), .SIGNEDP(n13214));
    defparam mult_966.REG_INPUTA_CLK = "NONE";
    defparam mult_966.REG_INPUTA_CE = "CE0";
    defparam mult_966.REG_INPUTA_RST = "RST0";
    defparam mult_966.REG_INPUTB_CLK = "NONE";
    defparam mult_966.REG_INPUTB_CE = "CE0";
    defparam mult_966.REG_INPUTB_RST = "RST0";
    defparam mult_966.REG_INPUTC_CLK = "NONE";
    defparam mult_966.REG_INPUTC_CE = "CE0";
    defparam mult_966.REG_INPUTC_RST = "RST0";
    defparam mult_966.REG_PIPELINE_CLK = "NONE";
    defparam mult_966.REG_PIPELINE_CE = "CE0";
    defparam mult_966.REG_PIPELINE_RST = "RST0";
    defparam mult_966.REG_OUTPUT_CLK = "NONE";
    defparam mult_966.REG_OUTPUT_CE = "CE0";
    defparam mult_966.REG_OUTPUT_RST = "RST0";
    defparam mult_966.CLK0_DIV = "ENABLED";
    defparam mult_966.CLK1_DIV = "ENABLED";
    defparam mult_966.CLK2_DIV = "ENABLED";
    defparam mult_966.CLK3_DIV = "ENABLED";
    defparam mult_966.HIGHSPEED_CLK = "NONE";
    defparam mult_966.GSR = "DISABLED";
    defparam mult_966.CAS_MATCH_REG = "FALSE";
    defparam mult_966.SOURCEB_MODE = "B_SHIFT";
    defparam mult_966.MULT_BYPASS = "DISABLED";
    defparam mult_966.RESETMODE = "SYNC";
    MULT18X18D mult_8 (.A17(\shift_16_dout_i[17] ), .A16(\shift_16_dout_i[16] ), 
            .A15(\shift_16_dout_i[15] ), .A14(\shift_16_dout_i[14] ), .A13(\shift_16_dout_i[13] ), 
            .A12(\shift_16_dout_i[12] ), .A11(\shift_16_dout_i[11] ), .A10(\shift_16_dout_i[10] ), 
            .A9(\shift_16_dout_i[9] ), .A8(\shift_16_dout_i[8] ), .A7(op_i_23__N_1154[7]), 
            .A6(op_i_23__N_1154[6]), .A5(op_i_23__N_1154[5]), .A4(op_i_23__N_1154[4]), 
            .A3(op_i_23__N_1154[3]), .A2(op_i_23__N_1154[2]), .A1(op_i_23__N_1154[1]), 
            .A0(op_i_23__N_1154[0]), .B17(n12368), .B16(n12368), .B15(n12368), 
            .B14(n12368), .B13(n12368), .B12(n12368), .B11(n12368), 
            .B10(n12368), .B9(n12353), .B8(n12352), .B7(n12351), .B6(n12350), 
            .B5(n12349), .B4(n12348), .B3(n12347), .B2(n12346), .B1(n12345), 
            .B0(n12344), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18107), 
            .ROA16(n18106), .ROA15(n18105), .ROA14(n18104), .ROA13(n18103), 
            .ROA12(n18102), .ROA11(n18101), .ROA10(n18100), .ROA9(n18099), 
            .ROA8(n18098), .ROA7(n18097), .ROA6(n18096), .ROA5(n18095), 
            .ROA4(n18094), .ROA3(n18093), .ROA2(n18092), .ROA1(n18091), 
            .ROA0(n18090), .ROB17(n18125), .ROB16(n18124), .ROB15(n18123), 
            .ROB14(n18122), .ROB13(n18121), .ROB12(n18120), .ROB11(n18119), 
            .ROB10(n18118), .ROB9(n18117), .ROB8(n18116), .ROB7(n18115), 
            .ROB6(n18114), .ROB5(n18113), .ROB4(n18112), .ROB3(n18111), 
            .ROB2(n18110), .ROB1(n18109), .ROB0(n18108), .P35(n18162), 
            .P34(n18161), .P33(n18160), .P32(n18159), .P31(n18158), 
            .P30(n18157), .P29(n18156), .P28(n18155), .P27(n18154), 
            .P26(n18153), .P25(n18152), .P24(n18151), .P23(n18150), 
            .P22(n18149), .P21(n18148), .P20(n18147), .P19(n18146), 
            .P18(n18145), .P17(n18144), .P16(n18143), .P15(n18142), 
            .P14(n18141), .P13(n18140), .P12(n18139), .P11(n18138), 
            .P10(n18137), .P9(n18136), .P8(n18135), .P7(n18134), .P6(n18133), 
            .P5(n18132), .P4(n18131), .P3(n18130), .P2(n18129), .P1(n18128), 
            .P0(n18127), .SIGNEDP(n18126));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam mult_8.REG_INPUTA_CLK = "NONE";
    defparam mult_8.REG_INPUTA_CE = "CE0";
    defparam mult_8.REG_INPUTA_RST = "RST0";
    defparam mult_8.REG_INPUTB_CLK = "NONE";
    defparam mult_8.REG_INPUTB_CE = "CE0";
    defparam mult_8.REG_INPUTB_RST = "RST0";
    defparam mult_8.REG_INPUTC_CLK = "NONE";
    defparam mult_8.REG_INPUTC_CE = "CE0";
    defparam mult_8.REG_INPUTC_RST = "RST0";
    defparam mult_8.REG_PIPELINE_CLK = "NONE";
    defparam mult_8.REG_PIPELINE_CE = "CE0";
    defparam mult_8.REG_PIPELINE_RST = "RST0";
    defparam mult_8.REG_OUTPUT_CLK = "NONE";
    defparam mult_8.REG_OUTPUT_CE = "CE0";
    defparam mult_8.REG_OUTPUT_RST = "RST0";
    defparam mult_8.CLK0_DIV = "ENABLED";
    defparam mult_8.CLK1_DIV = "ENABLED";
    defparam mult_8.CLK2_DIV = "ENABLED";
    defparam mult_8.CLK3_DIV = "ENABLED";
    defparam mult_8.HIGHSPEED_CLK = "NONE";
    defparam mult_8.GSR = "DISABLED";
    defparam mult_8.CAS_MATCH_REG = "FALSE";
    defparam mult_8.SOURCEB_MODE = "B_SHIFT";
    defparam mult_8.MULT_BYPASS = "DISABLED";
    defparam mult_8.RESETMODE = "SYNC";
    MULT18X18D lat_mult_70 (.A17(\shift_16_dout_i[23] ), .A16(\shift_16_dout_i[23] ), 
            .A15(\shift_16_dout_i[23] ), .A14(\shift_16_dout_i[23] ), .A13(\shift_16_dout_i[23] ), 
            .A12(\shift_16_dout_i[23] ), .A11(\shift_16_dout_i[23] ), .A10(\shift_16_dout_i[23] ), 
            .A9(\shift_16_dout_i[23] ), .A8(\shift_16_dout_i[23] ), .A7(\shift_16_dout_i[23] ), 
            .A6(\shift_16_dout_i[23] ), .A5(\shift_16_dout_i[23] ), .A4(\shift_16_dout_i[22] ), 
            .A3(\shift_16_dout_i[21] ), .A2(\shift_16_dout_i[20] ), .A1(\shift_16_dout_i[19] ), 
            .A0(\shift_16_dout_i[18] ), .B17(n12368), .B16(n12368), .B15(n12368), 
            .B14(n12368), .B13(n12368), .B12(n12368), .B11(n12368), 
            .B10(n12368), .B9(n12353), .B8(n12352), .B7(n12351), .B6(n12350), 
            .B5(n12349), .B4(n12348), .B3(n12347), .B2(n12346), .B1(n12345), 
            .B0(n12344), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18180), 
            .ROA16(n18179), .ROA15(n18178), .ROA14(n18177), .ROA13(n18176), 
            .ROA12(n18175), .ROA11(n18174), .ROA10(n18173), .ROA9(n18172), 
            .ROA8(n18171), .ROA7(n18170), .ROA6(n18169), .ROA5(n18168), 
            .ROA4(n18167), .ROA3(n18166), .ROA2(n18165), .ROA1(n18164), 
            .ROA0(n18163), .ROB17(n18198), .ROB16(n18197), .ROB15(n18196), 
            .ROB14(n18195), .ROB13(n18194), .ROB12(n18193), .ROB11(n18192), 
            .ROB10(n18191), .ROB9(n18190), .ROB8(n18189), .ROB7(n18188), 
            .ROB6(n18187), .ROB5(n18186), .ROB4(n18185), .ROB3(n18184), 
            .ROB2(n18183), .ROB1(n18182), .ROB0(n18181), .P35(n18235), 
            .P34(n18234), .P33(n18233), .P32(n18232), .P31(n18231), 
            .P30(n18230), .P29(n18229), .P28(n18228), .P27(n18227), 
            .P26(n18226), .P25(n18225), .P24(n18224), .P23(n18223), 
            .P22(n18222), .P21(n18221), .P20(n18220), .P19(n18219), 
            .P18(n18218), .P17(n18217), .P16(n18216), .P15(n18215), 
            .P14(n18214), .P13(n18213), .P12(n18212), .P11(n18211), 
            .P10(n18210), .P9(n18209), .P8(n18208), .P7(n18207), .P6(n18206), 
            .P5(n18205), .P4(n18204), .P3(n18203), .P2(n18202), .P1(n18201), 
            .P0(n18200), .SIGNEDP(n18199));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_70.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_70.REG_INPUTA_CE = "CE0";
    defparam lat_mult_70.REG_INPUTA_RST = "RST0";
    defparam lat_mult_70.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_70.REG_INPUTB_CE = "CE0";
    defparam lat_mult_70.REG_INPUTB_RST = "RST0";
    defparam lat_mult_70.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_70.REG_INPUTC_CE = "CE0";
    defparam lat_mult_70.REG_INPUTC_RST = "RST0";
    defparam lat_mult_70.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_70.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_70.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_70.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_70.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_70.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_70.CLK0_DIV = "ENABLED";
    defparam lat_mult_70.CLK1_DIV = "ENABLED";
    defparam lat_mult_70.CLK2_DIV = "ENABLED";
    defparam lat_mult_70.CLK3_DIV = "ENABLED";
    defparam lat_mult_70.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_70.GSR = "DISABLED";
    defparam lat_mult_70.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_70.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_70.MULT_BYPASS = "DISABLED";
    defparam lat_mult_70.RESETMODE = "SYNC";
    MULT18X18D lat_mult_71 (.A17(\shift_16_dout_i[17] ), .A16(\shift_16_dout_i[16] ), 
            .A15(\shift_16_dout_i[15] ), .A14(\shift_16_dout_i[14] ), .A13(\shift_16_dout_i[13] ), 
            .A12(\shift_16_dout_i[12] ), .A11(\shift_16_dout_i[11] ), .A10(\shift_16_dout_i[10] ), 
            .A9(\shift_16_dout_i[9] ), .A8(\shift_16_dout_i[8] ), .A7(op_i_23__N_1154[7]), 
            .A6(op_i_23__N_1154[6]), .A5(op_i_23__N_1154[5]), .A4(op_i_23__N_1154[4]), 
            .A3(op_i_23__N_1154[3]), .A2(op_i_23__N_1154[2]), .A1(op_i_23__N_1154[1]), 
            .A0(op_i_23__N_1154[0]), .B17(n12368), .B16(n12368), .B15(n12368), 
            .B14(n12368), .B13(n12368), .B12(n12368), .B11(n12368), 
            .B10(n12368), .B9(n12368), .B8(n12368), .B7(n12368), .B6(n12368), 
            .B5(n12368), .B4(n12368), .B3(n12368), .B2(n12368), .B1(n12368), 
            .B0(n12368), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18253), 
            .ROA16(n18252), .ROA15(n18251), .ROA14(n18250), .ROA13(n18249), 
            .ROA12(n18248), .ROA11(n18247), .ROA10(n18246), .ROA9(n18245), 
            .ROA8(n18244), .ROA7(n18243), .ROA6(n18242), .ROA5(n18241), 
            .ROA4(n18240), .ROA3(n18239), .ROA2(n18238), .ROA1(n18237), 
            .ROA0(n18236), .ROB17(n18271), .ROB16(n18270), .ROB15(n18269), 
            .ROB14(n18268), .ROB13(n18267), .ROB12(n18266), .ROB11(n18265), 
            .ROB10(n18264), .ROB9(n18263), .ROB8(n18262), .ROB7(n18261), 
            .ROB6(n18260), .ROB5(n18259), .ROB4(n18258), .ROB3(n18257), 
            .ROB2(n18256), .ROB1(n18255), .ROB0(n18254), .P35(n18308), 
            .P34(n18307), .P33(n18306), .P32(n18305), .P31(n18304), 
            .P30(n18303), .P29(n18302), .P28(n18301), .P27(n18300), 
            .P26(n18299), .P25(n18298), .P24(n18297), .P23(n18296), 
            .P22(n18295), .P21(n18294), .P20(n18293), .P19(n18292), 
            .P18(n18291), .P17(n18290), .P16(n18289), .P15(n18288), 
            .P14(n18287), .P13(n18286), .P12(n18285), .P11(n18284), 
            .P10(n18283), .P9(n18282), .P8(n18281), .P7(n18280), .P6(n18279), 
            .P5(n18278), .P4(n18277), .P3(n18276), .P2(n18275), .P1(n18274), 
            .P0(n18273), .SIGNEDP(n18272));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_71.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_71.REG_INPUTA_CE = "CE0";
    defparam lat_mult_71.REG_INPUTA_RST = "RST0";
    defparam lat_mult_71.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_71.REG_INPUTB_CE = "CE0";
    defparam lat_mult_71.REG_INPUTB_RST = "RST0";
    defparam lat_mult_71.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_71.REG_INPUTC_CE = "CE0";
    defparam lat_mult_71.REG_INPUTC_RST = "RST0";
    defparam lat_mult_71.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_71.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_71.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_71.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_71.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_71.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_71.CLK0_DIV = "ENABLED";
    defparam lat_mult_71.CLK1_DIV = "ENABLED";
    defparam lat_mult_71.CLK2_DIV = "ENABLED";
    defparam lat_mult_71.CLK3_DIV = "ENABLED";
    defparam lat_mult_71.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_71.GSR = "DISABLED";
    defparam lat_mult_71.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_71.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_71.MULT_BYPASS = "DISABLED";
    defparam lat_mult_71.RESETMODE = "SYNC";
    MULT18X18D lat_mult_72 (.A17(\shift_16_dout_i[23] ), .A16(\shift_16_dout_i[23] ), 
            .A15(\shift_16_dout_i[23] ), .A14(\shift_16_dout_i[23] ), .A13(\shift_16_dout_i[23] ), 
            .A12(\shift_16_dout_i[23] ), .A11(\shift_16_dout_i[23] ), .A10(\shift_16_dout_i[23] ), 
            .A9(\shift_16_dout_i[23] ), .A8(\shift_16_dout_i[23] ), .A7(\shift_16_dout_i[23] ), 
            .A6(\shift_16_dout_i[23] ), .A5(\shift_16_dout_i[23] ), .A4(\shift_16_dout_i[22] ), 
            .A3(\shift_16_dout_i[21] ), .A2(\shift_16_dout_i[20] ), .A1(\shift_16_dout_i[19] ), 
            .A0(\shift_16_dout_i[18] ), .B17(n12368), .B16(n12368), .B15(n12368), 
            .B14(n12368), .B13(n12368), .B12(n12368), .B11(n12368), 
            .B10(n12368), .B9(n12368), .B8(n12368), .B7(n12368), .B6(n12368), 
            .B5(n12368), .B4(n12368), .B3(n12368), .B2(n12368), .B1(n12368), 
            .B0(n12368), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n18326), 
            .ROA16(n18325), .ROA15(n18324), .ROA14(n18323), .ROA13(n18322), 
            .ROA12(n18321), .ROA11(n18320), .ROA10(n18319), .ROA9(n18318), 
            .ROA8(n18317), .ROA7(n18316), .ROA6(n18315), .ROA5(n18314), 
            .ROA4(n18313), .ROA3(n18312), .ROA2(n18311), .ROA1(n18310), 
            .ROA0(n18309), .ROB17(n18344), .ROB16(n18343), .ROB15(n18342), 
            .ROB14(n18341), .ROB13(n18340), .ROB12(n18339), .ROB11(n18338), 
            .ROB10(n18337), .ROB9(n18336), .ROB8(n18335), .ROB7(n18334), 
            .ROB6(n18333), .ROB5(n18332), .ROB4(n18331), .ROB3(n18330), 
            .ROB2(n18329), .ROB1(n18328), .ROB0(n18327), .P35(n18381), 
            .P34(n18380), .P33(n18379), .P32(n18378), .P31(n18377), 
            .P30(n18376), .P29(n18375), .P28(n18374), .P27(n18373), 
            .P26(n18372), .P25(n18371), .P24(n18370), .P23(n18369), 
            .P22(n18368), .P21(n18367), .P20(n18366), .P19(n18365), 
            .P18(n18364), .P17(n18363), .P16(n18362), .P15(n18361), 
            .P14(n18360), .P13(n18359), .P12(n18358), .P11(n18357), 
            .P10(n18356), .P9(n18355), .P8(n18354), .P7(n18353), .P6(n18352), 
            .P5(n18351), .P4(n18350), .P3(n18349), .P2(n18348), .P1(n18347), 
            .P0(n18346), .SIGNEDP(n18345));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_72.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_72.REG_INPUTA_CE = "CE0";
    defparam lat_mult_72.REG_INPUTA_RST = "RST0";
    defparam lat_mult_72.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_72.REG_INPUTB_CE = "CE0";
    defparam lat_mult_72.REG_INPUTB_RST = "RST0";
    defparam lat_mult_72.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_72.REG_INPUTC_CE = "CE0";
    defparam lat_mult_72.REG_INPUTC_RST = "RST0";
    defparam lat_mult_72.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_72.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_72.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_72.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_72.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_72.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_72.CLK0_DIV = "ENABLED";
    defparam lat_mult_72.CLK1_DIV = "ENABLED";
    defparam lat_mult_72.CLK2_DIV = "ENABLED";
    defparam lat_mult_72.CLK3_DIV = "ENABLED";
    defparam lat_mult_72.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_72.GSR = "DISABLED";
    defparam lat_mult_72.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_72.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_72.MULT_BYPASS = "DISABLED";
    defparam lat_mult_72.RESETMODE = "SYNC";
    LUT4 mux_399_i23_3_lut_4_lut (.A(op_r_23__N_1106[22]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[22] ), .Z(n7539)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i23_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13829_3_lut_4_lut (.A(op_r_23__N_1106[22]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[30] ), .Z(n31574)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13829_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i24_3_lut_4_lut (.A(op_r_23__N_1106[23]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[23] ), .Z(n7538)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i24_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13827_3_lut_4_lut (.A(op_r_23__N_1106[23]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[31] ), .Z(n31572)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13827_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i23_3_lut_4_lut (.A(op_i_23__N_1154[22]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[22] ), .Z(n7486)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i23_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13633_3_lut_4_lut (.A(op_i_23__N_1154[22]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[30] ), .Z(n31378)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13633_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i24_3_lut_4_lut (.A(op_i_23__N_1154[23]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[23] ), .Z(n7485)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i24_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13631_3_lut_4_lut (.A(op_i_23__N_1154[23]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[31] ), .Z(n31376)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13631_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i21_3_lut_4_lut (.A(op_r_23__N_1106[20]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[20] ), .Z(n7541)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i21_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13833_3_lut_4_lut (.A(op_r_23__N_1106[20]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[28] ), .Z(n31578)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13833_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i22_3_lut_4_lut (.A(op_r_23__N_1106[21]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[21] ), .Z(n7540)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i22_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13831_3_lut_4_lut (.A(op_r_23__N_1106[21]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[29] ), .Z(n31576)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13831_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i21_3_lut_4_lut (.A(op_i_23__N_1154[20]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[20] ), .Z(n7488)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i21_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13637_3_lut_4_lut (.A(op_i_23__N_1154[20]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[28] ), .Z(n31382)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13637_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i22_3_lut_4_lut (.A(op_i_23__N_1154[21]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[21] ), .Z(n7487)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i22_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13635_3_lut_4_lut (.A(op_i_23__N_1154[21]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[29] ), .Z(n31380)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13635_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i19_3_lut_4_lut (.A(op_r_23__N_1106[18]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[18] ), .Z(n7543)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i19_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13837_3_lut_4_lut (.A(op_r_23__N_1106[18]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[26] ), .Z(n31582)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13837_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i20_3_lut_4_lut (.A(op_r_23__N_1106[19]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[19] ), .Z(n7542)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13835_3_lut_4_lut (.A(op_r_23__N_1106[19]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[27] ), .Z(n31580)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13835_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i19_3_lut_4_lut (.A(op_i_23__N_1154[18]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[18] ), .Z(n7490)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i19_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13641_3_lut_4_lut (.A(op_i_23__N_1154[18]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[26] ), .Z(n31386)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13641_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i20_3_lut_4_lut (.A(op_i_23__N_1154[19]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[19] ), .Z(n7489)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13639_3_lut_4_lut (.A(op_i_23__N_1154[19]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[27] ), .Z(n31384)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13639_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i17_3_lut_4_lut (.A(op_r_23__N_1106[16]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[16] ), .Z(n7545)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13841_3_lut_4_lut (.A(op_r_23__N_1106[16]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[24] ), .Z(n31586)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13841_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i18_3_lut_4_lut (.A(op_r_23__N_1106[17]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[17] ), .Z(n7544)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i18_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13839_3_lut_4_lut (.A(op_r_23__N_1106[17]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[25] ), .Z(n31584)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13839_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i17_3_lut_4_lut (.A(op_i_23__N_1154[16]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[16] ), .Z(n7492)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13645_3_lut_4_lut (.A(op_i_23__N_1154[16]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[24] ), .Z(n31390)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13645_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i18_3_lut_4_lut (.A(op_i_23__N_1154[17]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[17] ), .Z(n7491)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i18_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13643_3_lut_4_lut (.A(op_i_23__N_1154[17]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[25] ), .Z(n31388)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13643_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i15_3_lut_4_lut (.A(op_r_23__N_1106[14]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[14] ), .Z(n7547)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i15_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13845_3_lut_4_lut (.A(op_r_23__N_1106[14]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[22] ), .Z(n31590)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13845_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i16_3_lut_4_lut (.A(op_r_23__N_1106[15]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[15] ), .Z(n7546)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i16_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13843_3_lut_4_lut (.A(op_r_23__N_1106[15]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[23] ), .Z(n31588)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13843_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i15_3_lut_4_lut (.A(op_i_23__N_1154[14]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[14] ), .Z(n7494)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i15_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13649_3_lut_4_lut (.A(op_i_23__N_1154[14]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[22] ), .Z(n31394)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13649_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i16_3_lut_4_lut (.A(op_i_23__N_1154[15]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[15] ), .Z(n7493)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i16_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13647_3_lut_4_lut (.A(op_i_23__N_1154[15]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[23] ), .Z(n31392)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13647_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i13_3_lut_4_lut (.A(op_r_23__N_1106[12]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[12] ), .Z(n7549)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13849_3_lut_4_lut (.A(op_r_23__N_1106[12]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[20] ), .Z(n31594)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13849_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i14_3_lut_4_lut (.A(op_r_23__N_1106[13]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[13] ), .Z(n7548)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i14_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13847_3_lut_4_lut (.A(op_r_23__N_1106[13]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[21] ), .Z(n31592)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13847_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i13_3_lut_4_lut (.A(op_i_23__N_1154[12]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[12] ), .Z(n7496)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13653_3_lut_4_lut (.A(op_i_23__N_1154[12]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[20] ), .Z(n31398)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13653_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i14_3_lut_4_lut (.A(op_i_23__N_1154[13]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[13] ), .Z(n7495)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i14_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13651_3_lut_4_lut (.A(op_i_23__N_1154[13]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[21] ), .Z(n31396)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13651_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i11_3_lut_4_lut (.A(op_r_23__N_1106[10]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[10] ), .Z(n7551)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i11_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13853_3_lut_4_lut (.A(op_r_23__N_1106[10]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[18] ), .Z(n31598)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13853_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i12_3_lut_4_lut (.A(op_r_23__N_1106[11]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[11] ), .Z(n7550)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i12_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13851_3_lut_4_lut (.A(op_r_23__N_1106[11]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[19] ), .Z(n31596)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13851_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i11_3_lut_4_lut (.A(op_i_23__N_1154[10]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[10] ), .Z(n7498)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i11_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13657_3_lut_4_lut (.A(op_i_23__N_1154[10]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[18] ), .Z(n31402)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13657_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i12_3_lut_4_lut (.A(op_i_23__N_1154[11]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[11] ), .Z(n7497)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i12_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13655_3_lut_4_lut (.A(op_i_23__N_1154[11]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[19] ), .Z(n31400)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13655_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i9_3_lut_4_lut (.A(op_r_23__N_1106[8]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[8] ), .Z(n7553)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13857_3_lut_4_lut (.A(op_r_23__N_1106[8]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[16] ), .Z(n31602)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13857_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_399_i10_3_lut_4_lut (.A(op_r_23__N_1106[9]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_r[9] ), .Z(n7552)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_399_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13855_3_lut_4_lut (.A(op_r_23__N_1106[9]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_r_23__N_1082[17] ), .Z(n31600)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13855_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i9_3_lut_4_lut (.A(op_i_23__N_1154[8]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[8] ), .Z(n7500)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13661_3_lut_4_lut (.A(op_i_23__N_1154[8]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[16] ), .Z(n31406)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13661_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_395_i10_3_lut_4_lut (.A(op_i_23__N_1154[9]), .B(clk_c_enable_2310), 
         .C(n34755), .D(\shift_8_dout_i[9] ), .Z(n7499)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam mux_395_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13659_3_lut_4_lut (.A(op_i_23__N_1154[9]), .B(clk_c_enable_2310), 
         .C(n34756), .D(\op_i_23__N_1130[17] ), .Z(n31404)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13659_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_369_i9_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[8] ), 
         .D(\delay_r_23__N_1178[8] ), .Z(\dout_r_23__N_2506[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i9_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i10_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[9] ), 
         .D(\delay_r_23__N_1178[9] ), .Z(\dout_r_23__N_2506[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i10_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i11_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[10] ), 
         .D(\delay_r_23__N_1178[10] ), .Z(\dout_r_23__N_2506[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i12_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[11] ), 
         .D(\delay_r_23__N_1178[11] ), .Z(\dout_r_23__N_2506[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i13_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[12] ), 
         .D(\delay_r_23__N_1178[12] ), .Z(\dout_r_23__N_2506[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i13_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i14_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[13] ), 
         .D(\delay_r_23__N_1178[13] ), .Z(\dout_r_23__N_2506[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i14_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i15_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[14] ), 
         .D(\delay_r_23__N_1178[14] ), .Z(\dout_r_23__N_2506[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i15_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i16_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[15] ), 
         .D(\delay_r_23__N_1178[15] ), .Z(\dout_r_23__N_2506[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i16_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i17_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[16] ), 
         .D(\delay_r_23__N_1178[16] ), .Z(\dout_r_23__N_2506[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i17_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i18_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[17] ), 
         .D(\delay_r_23__N_1178[17] ), .Z(\dout_r_23__N_2506[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i18_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i19_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[18] ), 
         .D(\delay_r_23__N_1178[18] ), .Z(\dout_r_23__N_2506[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i19_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i20_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[23] ), 
         .D(\delay_r_23__N_1178[19] ), .Z(\dout_r_23__N_2506[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i20_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i21_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[23] ), 
         .D(\delay_r_23__N_1178[20] ), .Z(\dout_r_23__N_2506[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i21_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i22_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[23] ), 
         .D(\delay_r_23__N_1178[21] ), .Z(\dout_r_23__N_2506[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i22_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i23_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[23] ), 
         .D(\delay_r_23__N_1178[22] ), .Z(\dout_r_23__N_2506[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i23_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_369_i24_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_r_reg[23] ), 
         .D(\delay_r_23__N_1178[23] ), .Z(\dout_r_23__N_2506[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_369_i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i9_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[8] ), 
         .D(\delay_i_23__N_1202[8] ), .Z(\dout_i_23__N_3274[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i9_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i10_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[9] ), 
         .D(\delay_i_23__N_1202[9] ), .Z(\dout_i_23__N_3274[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i10_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i11_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[10] ), 
         .D(\delay_i_23__N_1202[10] ), .Z(\dout_i_23__N_3274[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i12_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[11] ), 
         .D(\delay_i_23__N_1202[11] ), .Z(\dout_i_23__N_3274[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i13_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[12] ), 
         .D(\delay_i_23__N_1202[12] ), .Z(\dout_i_23__N_3274[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i13_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i14_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[13] ), 
         .D(\delay_i_23__N_1202[13] ), .Z(\dout_i_23__N_3274[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i14_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i15_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[14] ), 
         .D(\delay_i_23__N_1202[14] ), .Z(\dout_i_23__N_3274[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i15_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i16_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[15] ), 
         .D(\delay_i_23__N_1202[15] ), .Z(\dout_i_23__N_3274[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i16_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i17_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[16] ), 
         .D(\delay_i_23__N_1202[16] ), .Z(\dout_i_23__N_3274[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i17_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i18_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[17] ), 
         .D(\delay_i_23__N_1202[17] ), .Z(\dout_i_23__N_3274[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i18_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i19_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[18] ), 
         .D(\delay_i_23__N_1202[18] ), .Z(\dout_i_23__N_3274[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i19_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i20_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[23] ), 
         .D(\delay_i_23__N_1202[19] ), .Z(\dout_i_23__N_3274[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i20_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i21_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[23] ), 
         .D(\delay_i_23__N_1202[20] ), .Z(\dout_i_23__N_3274[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i21_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i22_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[23] ), 
         .D(\delay_i_23__N_1202[21] ), .Z(\dout_i_23__N_3274[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i22_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i23_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[23] ), 
         .D(\delay_i_23__N_1202[22] ), .Z(\dout_i_23__N_3274[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i23_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_367_i24_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\din_i_reg[23] ), 
         .D(\delay_i_23__N_1202[23] ), .Z(\dout_i_23__N_3274[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam mux_367_i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i15_2_lut_rep_436 (.A(\count[5] ), .B(\count[4] ), .Z(clk_c_enable_2310)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i15_2_lut_rep_436.init = 16'h6666;
    LUT4 i12838_2_lut_rep_297_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[14]), 
         .Z(n34659)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12838_2_lut_rep_297_3_lut.init = 16'h6060;
    LUT4 i12864_2_lut_rep_290_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[17]), 
         .Z(n34652)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12864_2_lut_rep_290_3_lut.init = 16'h6060;
    LUT4 i12863_2_lut_rep_289_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[16]), 
         .Z(n34651)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12863_2_lut_rep_289_3_lut.init = 16'h6060;
    LUT4 i12841_2_lut_rep_288_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[17]), 
         .Z(n34650)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12841_2_lut_rep_288_3_lut.init = 16'h6060;
    LUT4 i12840_2_lut_rep_287_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[16]), 
         .Z(n34649)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12840_2_lut_rep_287_3_lut.init = 16'h6060;
    LUT4 i12866_2_lut_rep_280_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[19]), 
         .Z(n34642)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12866_2_lut_rep_280_3_lut.init = 16'h6060;
    LUT4 i12865_2_lut_rep_279_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[18]), 
         .Z(n34641)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12865_2_lut_rep_279_3_lut.init = 16'h6060;
    LUT4 i12843_2_lut_rep_278_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[19]), 
         .Z(n34640)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12843_2_lut_rep_278_3_lut.init = 16'h6060;
    LUT4 i12842_2_lut_rep_277_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[18]), 
         .Z(n34639)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12842_2_lut_rep_277_3_lut.init = 16'h6060;
    LUT4 i12868_2_lut_rep_268_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[21]), 
         .Z(n34630)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12868_2_lut_rep_268_3_lut.init = 16'h6060;
    LUT4 i12867_2_lut_rep_267_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[20]), 
         .Z(n34629)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12867_2_lut_rep_267_3_lut.init = 16'h6060;
    LUT4 i12845_2_lut_rep_266_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[21]), 
         .Z(n34628)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12845_2_lut_rep_266_3_lut.init = 16'h6060;
    LUT4 i12844_2_lut_rep_265_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[20]), 
         .Z(n34627)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12844_2_lut_rep_265_3_lut.init = 16'h6060;
    LUT4 i12870_2_lut_rep_256_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[23]), 
         .Z(n34618)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12870_2_lut_rep_256_3_lut.init = 16'h6060;
    LUT4 i12869_2_lut_rep_255_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[22]), 
         .Z(n34617)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12869_2_lut_rep_255_3_lut.init = 16'h6060;
    LUT4 i12847_2_lut_rep_254_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[23]), 
         .Z(n34616)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12847_2_lut_rep_254_3_lut.init = 16'h6060;
    LUT4 i12846_2_lut_rep_253_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[22]), 
         .Z(n34615)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12846_2_lut_rep_253_3_lut.init = 16'h6060;
    LUT4 i12839_2_lut_rep_298_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[15]), 
         .Z(n34660)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12839_2_lut_rep_298_3_lut.init = 16'h6060;
    LUT4 i12861_2_lut_rep_299_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[14]), 
         .Z(n34661)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12861_2_lut_rep_299_3_lut.init = 16'h6060;
    LUT4 i12862_2_lut_rep_300_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[15]), 
         .Z(n34662)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12862_2_lut_rep_300_3_lut.init = 16'h6060;
    LUT4 i12836_2_lut_rep_307_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[12]), 
         .Z(n34669)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12836_2_lut_rep_307_3_lut.init = 16'h6060;
    LUT4 i12837_2_lut_rep_308_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[13]), 
         .Z(n34670)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12837_2_lut_rep_308_3_lut.init = 16'h6060;
    LUT4 i12859_2_lut_rep_309_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[12]), 
         .Z(n34671)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12859_2_lut_rep_309_3_lut.init = 16'h6060;
    LUT4 i12860_2_lut_rep_310_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[13]), 
         .Z(n34672)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12860_2_lut_rep_310_3_lut.init = 16'h6060;
    LUT4 i12834_2_lut_rep_313_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[10]), 
         .Z(n34675)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12834_2_lut_rep_313_3_lut.init = 16'h6060;
    LUT4 i12835_2_lut_rep_314_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[11]), 
         .Z(n34676)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12835_2_lut_rep_314_3_lut.init = 16'h6060;
    LUT4 i12857_2_lut_rep_315_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[10]), 
         .Z(n34677)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12857_2_lut_rep_315_3_lut.init = 16'h6060;
    LUT4 i12858_2_lut_rep_316_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[11]), 
         .Z(n34678)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12858_2_lut_rep_316_3_lut.init = 16'h6060;
    LUT4 i12832_2_lut_rep_321_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[8]), 
         .Z(n34683)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12832_2_lut_rep_321_3_lut.init = 16'h6060;
    LUT4 i12833_2_lut_rep_322_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_r_23__N_1106[9]), 
         .Z(n34684)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12833_2_lut_rep_322_3_lut.init = 16'h6060;
    LUT4 i12855_2_lut_rep_323_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[8]), 
         .Z(n34685)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12855_2_lut_rep_323_3_lut.init = 16'h6060;
    LUT4 i12856_2_lut_rep_324_3_lut (.A(\count[5] ), .B(\count[4] ), .C(op_i_23__N_1154[9]), 
         .Z(n34686)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12856_2_lut_rep_324_3_lut.init = 16'h6060;
    LUT4 i178_2_lut_rep_405_3_lut (.A(\count[5] ), .B(\count[4] ), .C(valid), 
         .Z(clk_c_enable_1419)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i178_2_lut_rep_405_3_lut.init = 16'hf6f6;
    
endmodule
//
// Verilog Description of module radix2_U0
//

module radix2_U0 (\op_r_23__N_1106[14] , n34841, n30179, \delay_r_23__N_1178[14] , 
            \dout_r_23__N_5681[14] , \op_i_23__N_1154[13] , \delay_i_23__N_1202[13] , 
            \dout_i_23__N_5777[13] , \op_r_23__N_1106[21] , \delay_r_23__N_1178[21] , 
            \dout_r_23__N_5681[21] , \op_i_23__N_1154[12] , \delay_i_23__N_1202[12] , 
            \dout_i_23__N_5777[12] , \op_r_23__N_1226[0] , \op_r_23__N_1226[1] , 
            \op_r_23__N_1226[2] , \op_r_23__N_1226[3] , \op_r_23__N_1226[4] , 
            \op_r_23__N_1226[5] , \op_r_23__N_1226[6] , \op_r_23__N_1226[7] , 
            \op_r_23__N_1226[8] , \op_r_23__N_1226[9] , \op_r_23__N_1226[10] , 
            \op_r_23__N_1226[11] , \op_r_23__N_1226[12] , \op_r_23__N_1226[13] , 
            \op_r_23__N_1226[14] , \op_r_23__N_1226[15] , \op_r_23__N_1226[16] , 
            \op_r_23__N_1226[17] , \op_r_23__N_1226[18] , \op_r_23__N_1226[19] , 
            \op_r_23__N_1226[20] , \op_r_23__N_1226[21] , \op_r_23__N_1226[22] , 
            \op_r_23__N_1226[23] , \op_r_23__N_1226[24] , \op_r_23__N_1226[25] , 
            \op_r_23__N_1226[26] , \op_r_23__N_1226[27] , \op_r_23__N_1226[28] , 
            \op_r_23__N_1226[29] , \op_r_23__N_1226[30] , \op_r_23__N_1226[31] , 
            GND_net, VCC_net, n12170, n12171, n12172, n12173, n12174, 
            n12175, n12176, \rom2_w_r[8] , n12152, n12153, n12154, 
            n12155, n12156, n12157, n12158, n12159, n12160, n12161, 
            n12162, n12163, n12164, n12165, n12166, n12167, n12168, 
            n12169, \op_r_23__N_1106[15] , \delay_r_23__N_1178[15] , \dout_r_23__N_5681[15] , 
            \op_r_23__N_1106[13] , \delay_r_23__N_1178[13] , \dout_r_23__N_5681[13] , 
            \op_r_23__N_1106[12] , \delay_r_23__N_1178[12] , \dout_r_23__N_5681[12] , 
            \op_i_23__N_1154[11] , \delay_i_23__N_1202[11] , \dout_i_23__N_5777[11] , 
            \op_r_23__N_1106[20] , \delay_r_23__N_1178[20] , \dout_r_23__N_5681[20] , 
            \op_i_23__N_1154[10] , \delay_i_23__N_1202[10] , \dout_i_23__N_5777[10] , 
            n34795, n114, shift_2_dout_i, \op_r_23__N_1268[0] , \op_r_23__N_1268[1] , 
            \op_r_23__N_1268[2] , \op_r_23__N_1268[3] , \op_r_23__N_1268[4] , 
            \op_r_23__N_1268[5] , \op_r_23__N_1268[6] , \op_r_23__N_1268[7] , 
            \op_r_23__N_1268[8] , \op_r_23__N_1268[9] , \op_r_23__N_1268[10] , 
            \op_r_23__N_1268[11] , \op_r_23__N_1268[12] , \op_r_23__N_1268[13] , 
            \op_r_23__N_1268[14] , \op_r_23__N_1268[15] , \op_r_23__N_1268[16] , 
            \op_r_23__N_1268[17] , \op_r_23__N_1268[18] , \op_r_23__N_1268[19] , 
            \op_r_23__N_1268[20] , \op_r_23__N_1268[21] , \op_r_23__N_1268[22] , 
            \op_r_23__N_1268[23] , \op_r_23__N_1268[24] , \op_r_23__N_1268[25] , 
            \op_r_23__N_1268[26] , \op_r_23__N_1268[27] , \op_r_23__N_1268[28] , 
            \op_r_23__N_1268[29] , \op_r_23__N_1268[30] , \op_r_23__N_1268[31] , 
            n8977, n8976, n8975, n8974, n8973, n8972, n8971, n8970, 
            n8969, n8968, n8967, n8966, n8965, n8964, n8963, n8962, 
            n8961, n8960, n8959, n8958, n8957, n8956, n8955, n8954, 
            n8953, n8952, \op_i_23__N_1154[19] , \delay_i_23__N_1202[19] , 
            \dout_i_23__N_5777[19] , n319, \rom4_w_i[12] , n114_adj_33, 
            n11126, n11127, n11128, n11129, n11130, n11131, n11132, 
            n11133, n11134, n11135, n11136, n11137, n11138, n11139, 
            n11140, n11141, n11142, n11143, n120, n126, \op_i_23__N_1310[0] , 
            n123, n117, n111, \op_i_23__N_1310[2] , \op_i_23__N_1310[3] , 
            \op_i_23__N_1310[4] , \op_i_23__N_1310[5] , n89, n87, n88, 
            n85, n86, n83, n84, n81, n82, n79, n80, n77, n78, 
            n75, n76, n73, n74, n71, n72, n69, n70, n67, n68, 
            n65, n66, \op_i_23__N_1310[1] , n120_adj_34, n126_adj_35, 
            n34777, \op_i_23__N_1310[0]_adj_36 , n123_adj_37, n117_adj_38, 
            n111_adj_39, \op_i_23__N_1310[2]_adj_40 , \op_i_23__N_1310[3]_adj_41 , 
            \op_i_23__N_1310[4]_adj_42 , \op_i_23__N_1310[5]_adj_43 , n89_adj_44, 
            n87_adj_45, n88_adj_46, n85_adj_47, n86_adj_48, n83_adj_49, 
            n84_adj_50, n81_adj_51, n82_adj_52, n79_adj_53, n80_adj_54, 
            n77_adj_55, n78_adj_56, n75_adj_57, n76_adj_58, n73_adj_59, 
            n74_adj_60, n71_adj_61, n72_adj_62, n69_adj_63, n70_adj_64, 
            n67_adj_65, n68_adj_66, n65_adj_67, n66_adj_68, \op_i_23__N_1310[1]_adj_69 , 
            \op_r_23__N_1106[19] , \delay_r_23__N_1178[19] , \dout_r_23__N_5681[19] , 
            \op_r_23__N_1106[11] , \delay_r_23__N_1178[11] , \dout_r_23__N_5681[11] , 
            \op_r_23__N_1106[10] , \delay_r_23__N_1178[10] , \dout_r_23__N_5681[10] , 
            \op_i_23__N_1154[9] , \delay_i_23__N_1202[9] , \dout_i_23__N_5777[9] , 
            \op_r_23__N_1106[18] , \delay_r_23__N_1178[18] , \dout_r_23__N_5681[18] , 
            \op_i_23__N_1154[8] , \delay_i_23__N_1202[8] , \dout_i_23__N_5777[8] , 
            \op_r_23__N_1106[9] , \delay_r_23__N_1178[9] , \dout_r_23__N_5681[9] , 
            \op_r_23__N_1106[8] , \delay_r_23__N_1178[8] , \dout_r_23__N_5681[8] , 
            \op_i_23__N_1154[7] , \delay_i_23__N_1202[7] , \dout_i_23__N_5777[7] , 
            \op_i_23__N_1154[6] , \delay_i_23__N_1202[6] , \dout_i_23__N_5777[6] , 
            \op_i_23__N_1154[17] , \delay_i_23__N_1202[17] , \dout_i_23__N_5777[17] , 
            \op_i_23__N_1154[23] , \delay_i_23__N_1202[23] , \dout_i_23__N_5777[23] , 
            \op_r_23__N_1106[23] , \delay_r_23__N_1178[23] , \dout_r_23__N_5681[23] , 
            \op_r_23__N_1106[22] , \delay_r_23__N_1178[22] , \dout_r_23__N_5681[22] , 
            \op_i_23__N_1154[21] , \delay_i_23__N_1202[21] , \dout_i_23__N_5777[21] , 
            \op_i_23__N_1154[16] , \delay_i_23__N_1202[16] , \dout_i_23__N_5777[16] , 
            \op_i_23__N_1154[20] , \delay_i_23__N_1202[20] , \dout_i_23__N_5777[20] , 
            \op_i_23__N_1154[5] , \delay_i_23__N_1202[5] , \dout_i_23__N_5777[5] , 
            \op_i_23__N_1154[4] , \delay_i_23__N_1202[4] , \dout_i_23__N_5777[4] , 
            \op_i_23__N_1154[3] , \delay_i_23__N_1202[3] , \dout_i_23__N_5777[3] , 
            \op_i_23__N_1154[22] , \delay_i_23__N_1202[22] , \dout_i_23__N_5777[22] , 
            \op_r_23__N_1106[7] , \delay_r_23__N_1178[7] , \dout_r_23__N_5681[7] , 
            \op_r_23__N_1106[6] , \delay_r_23__N_1178[6] , \dout_r_23__N_5681[6] , 
            \op_r_23__N_1106[5] , \delay_r_23__N_1178[5] , \dout_r_23__N_5681[5] , 
            \op_r_23__N_1106[4] , \delay_r_23__N_1178[4] , \dout_r_23__N_5681[4] , 
            \op_r_23__N_1106[17] , \delay_r_23__N_1178[17] , \dout_r_23__N_5681[17] , 
            \op_r_23__N_1106[3] , \delay_r_23__N_1178[3] , \dout_r_23__N_5681[3] , 
            \op_r_23__N_1106[2] , \delay_r_23__N_1178[2] , \dout_r_23__N_5681[2] , 
            \op_r_23__N_1106[16] , \delay_r_23__N_1178[16] , \dout_r_23__N_5681[16] , 
            \op_r_23__N_1106[1] , \delay_r_23__N_1178[1] , \dout_r_23__N_5681[1] , 
            \op_i_23__N_1154[15] , \delay_i_23__N_1202[15] , \dout_i_23__N_5777[15] , 
            \op_i_23__N_1154[14] , \delay_i_23__N_1202[14] , \dout_i_23__N_5777[14] ) /* synthesis syn_module_defined=1 */ ;
    input \op_r_23__N_1106[14] ;
    input n34841;
    input n30179;
    input \delay_r_23__N_1178[14] ;
    output \dout_r_23__N_5681[14] ;
    input \op_i_23__N_1154[13] ;
    input \delay_i_23__N_1202[13] ;
    output \dout_i_23__N_5777[13] ;
    input \op_r_23__N_1106[21] ;
    input \delay_r_23__N_1178[21] ;
    output \dout_r_23__N_5681[21] ;
    input \op_i_23__N_1154[12] ;
    input \delay_i_23__N_1202[12] ;
    output \dout_i_23__N_5777[12] ;
    output \op_r_23__N_1226[0] ;
    output \op_r_23__N_1226[1] ;
    output \op_r_23__N_1226[2] ;
    output \op_r_23__N_1226[3] ;
    output \op_r_23__N_1226[4] ;
    output \op_r_23__N_1226[5] ;
    output \op_r_23__N_1226[6] ;
    output \op_r_23__N_1226[7] ;
    output \op_r_23__N_1226[8] ;
    output \op_r_23__N_1226[9] ;
    output \op_r_23__N_1226[10] ;
    output \op_r_23__N_1226[11] ;
    output \op_r_23__N_1226[12] ;
    output \op_r_23__N_1226[13] ;
    output \op_r_23__N_1226[14] ;
    output \op_r_23__N_1226[15] ;
    output \op_r_23__N_1226[16] ;
    output \op_r_23__N_1226[17] ;
    output \op_r_23__N_1226[18] ;
    output \op_r_23__N_1226[19] ;
    output \op_r_23__N_1226[20] ;
    output \op_r_23__N_1226[21] ;
    output \op_r_23__N_1226[22] ;
    output \op_r_23__N_1226[23] ;
    output \op_r_23__N_1226[24] ;
    output \op_r_23__N_1226[25] ;
    output \op_r_23__N_1226[26] ;
    output \op_r_23__N_1226[27] ;
    output \op_r_23__N_1226[28] ;
    output \op_r_23__N_1226[29] ;
    output \op_r_23__N_1226[30] ;
    output \op_r_23__N_1226[31] ;
    input GND_net;
    input VCC_net;
    input n12170;
    input n12171;
    input n12172;
    input n12173;
    input n12174;
    input n12175;
    input n12176;
    input \rom2_w_r[8] ;
    input n12152;
    input n12153;
    input n12154;
    input n12155;
    input n12156;
    input n12157;
    input n12158;
    input n12159;
    input n12160;
    input n12161;
    input n12162;
    input n12163;
    input n12164;
    input n12165;
    input n12166;
    input n12167;
    input n12168;
    input n12169;
    input \op_r_23__N_1106[15] ;
    input \delay_r_23__N_1178[15] ;
    output \dout_r_23__N_5681[15] ;
    input \op_r_23__N_1106[13] ;
    input \delay_r_23__N_1178[13] ;
    output \dout_r_23__N_5681[13] ;
    input \op_r_23__N_1106[12] ;
    input \delay_r_23__N_1178[12] ;
    output \dout_r_23__N_5681[12] ;
    input \op_i_23__N_1154[11] ;
    input \delay_i_23__N_1202[11] ;
    output \dout_i_23__N_5777[11] ;
    input \op_r_23__N_1106[20] ;
    input \delay_r_23__N_1178[20] ;
    output \dout_r_23__N_5681[20] ;
    input \op_i_23__N_1154[10] ;
    input \delay_i_23__N_1202[10] ;
    output \dout_i_23__N_5777[10] ;
    input n34795;
    input n114;
    input [23:0]shift_2_dout_i;
    output \op_r_23__N_1268[0] ;
    output \op_r_23__N_1268[1] ;
    output \op_r_23__N_1268[2] ;
    output \op_r_23__N_1268[3] ;
    output \op_r_23__N_1268[4] ;
    output \op_r_23__N_1268[5] ;
    output \op_r_23__N_1268[6] ;
    output \op_r_23__N_1268[7] ;
    output \op_r_23__N_1268[8] ;
    output \op_r_23__N_1268[9] ;
    output \op_r_23__N_1268[10] ;
    output \op_r_23__N_1268[11] ;
    output \op_r_23__N_1268[12] ;
    output \op_r_23__N_1268[13] ;
    output \op_r_23__N_1268[14] ;
    output \op_r_23__N_1268[15] ;
    output \op_r_23__N_1268[16] ;
    output \op_r_23__N_1268[17] ;
    output \op_r_23__N_1268[18] ;
    output \op_r_23__N_1268[19] ;
    output \op_r_23__N_1268[20] ;
    output \op_r_23__N_1268[21] ;
    output \op_r_23__N_1268[22] ;
    output \op_r_23__N_1268[23] ;
    output \op_r_23__N_1268[24] ;
    output \op_r_23__N_1268[25] ;
    output \op_r_23__N_1268[26] ;
    output \op_r_23__N_1268[27] ;
    output \op_r_23__N_1268[28] ;
    output \op_r_23__N_1268[29] ;
    output \op_r_23__N_1268[30] ;
    output \op_r_23__N_1268[31] ;
    output n8977;
    output n8976;
    output n8975;
    output n8974;
    output n8973;
    output n8972;
    output n8971;
    output n8970;
    output n8969;
    output n8968;
    output n8967;
    output n8966;
    output n8965;
    output n8964;
    output n8963;
    output n8962;
    output n8961;
    output n8960;
    output n8959;
    output n8958;
    output n8957;
    output n8956;
    output n8955;
    output n8954;
    output n8953;
    output n8952;
    input \op_i_23__N_1154[19] ;
    input \delay_i_23__N_1202[19] ;
    output \dout_i_23__N_5777[19] ;
    input n319;
    input \rom4_w_i[12] ;
    input n114_adj_33;
    input n11126;
    input n11127;
    input n11128;
    input n11129;
    input n11130;
    input n11131;
    input n11132;
    input n11133;
    input n11134;
    input n11135;
    input n11136;
    input n11137;
    input n11138;
    input n11139;
    input n11140;
    input n11141;
    input n11142;
    input n11143;
    input n120;
    input n126;
    output \op_i_23__N_1310[0] ;
    input n123;
    input n117;
    input n111;
    output \op_i_23__N_1310[2] ;
    output \op_i_23__N_1310[3] ;
    output \op_i_23__N_1310[4] ;
    output \op_i_23__N_1310[5] ;
    output n89;
    output n87;
    output n88;
    output n85;
    output n86;
    output n83;
    output n84;
    output n81;
    output n82;
    output n79;
    output n80;
    output n77;
    output n78;
    output n75;
    output n76;
    output n73;
    output n74;
    output n71;
    output n72;
    output n69;
    output n70;
    output n67;
    output n68;
    output n65;
    output n66;
    output \op_i_23__N_1310[1] ;
    input n120_adj_34;
    input n126_adj_35;
    input n34777;
    output \op_i_23__N_1310[0]_adj_36 ;
    input n123_adj_37;
    input n117_adj_38;
    input n111_adj_39;
    output \op_i_23__N_1310[2]_adj_40 ;
    output \op_i_23__N_1310[3]_adj_41 ;
    output \op_i_23__N_1310[4]_adj_42 ;
    output \op_i_23__N_1310[5]_adj_43 ;
    output n89_adj_44;
    output n87_adj_45;
    output n88_adj_46;
    output n85_adj_47;
    output n86_adj_48;
    output n83_adj_49;
    output n84_adj_50;
    output n81_adj_51;
    output n82_adj_52;
    output n79_adj_53;
    output n80_adj_54;
    output n77_adj_55;
    output n78_adj_56;
    output n75_adj_57;
    output n76_adj_58;
    output n73_adj_59;
    output n74_adj_60;
    output n71_adj_61;
    output n72_adj_62;
    output n69_adj_63;
    output n70_adj_64;
    output n67_adj_65;
    output n68_adj_66;
    output n65_adj_67;
    output n66_adj_68;
    output \op_i_23__N_1310[1]_adj_69 ;
    input \op_r_23__N_1106[19] ;
    input \delay_r_23__N_1178[19] ;
    output \dout_r_23__N_5681[19] ;
    input \op_r_23__N_1106[11] ;
    input \delay_r_23__N_1178[11] ;
    output \dout_r_23__N_5681[11] ;
    input \op_r_23__N_1106[10] ;
    input \delay_r_23__N_1178[10] ;
    output \dout_r_23__N_5681[10] ;
    input \op_i_23__N_1154[9] ;
    input \delay_i_23__N_1202[9] ;
    output \dout_i_23__N_5777[9] ;
    input \op_r_23__N_1106[18] ;
    input \delay_r_23__N_1178[18] ;
    output \dout_r_23__N_5681[18] ;
    input \op_i_23__N_1154[8] ;
    input \delay_i_23__N_1202[8] ;
    output \dout_i_23__N_5777[8] ;
    input \op_r_23__N_1106[9] ;
    input \delay_r_23__N_1178[9] ;
    output \dout_r_23__N_5681[9] ;
    input \op_r_23__N_1106[8] ;
    input \delay_r_23__N_1178[8] ;
    output \dout_r_23__N_5681[8] ;
    input \op_i_23__N_1154[7] ;
    input \delay_i_23__N_1202[7] ;
    output \dout_i_23__N_5777[7] ;
    input \op_i_23__N_1154[6] ;
    input \delay_i_23__N_1202[6] ;
    output \dout_i_23__N_5777[6] ;
    input \op_i_23__N_1154[17] ;
    input \delay_i_23__N_1202[17] ;
    output \dout_i_23__N_5777[17] ;
    input \op_i_23__N_1154[23] ;
    input \delay_i_23__N_1202[23] ;
    output \dout_i_23__N_5777[23] ;
    input \op_r_23__N_1106[23] ;
    input \delay_r_23__N_1178[23] ;
    output \dout_r_23__N_5681[23] ;
    input \op_r_23__N_1106[22] ;
    input \delay_r_23__N_1178[22] ;
    output \dout_r_23__N_5681[22] ;
    input \op_i_23__N_1154[21] ;
    input \delay_i_23__N_1202[21] ;
    output \dout_i_23__N_5777[21] ;
    input \op_i_23__N_1154[16] ;
    input \delay_i_23__N_1202[16] ;
    output \dout_i_23__N_5777[16] ;
    input \op_i_23__N_1154[20] ;
    input \delay_i_23__N_1202[20] ;
    output \dout_i_23__N_5777[20] ;
    input \op_i_23__N_1154[5] ;
    input \delay_i_23__N_1202[5] ;
    output \dout_i_23__N_5777[5] ;
    input \op_i_23__N_1154[4] ;
    input \delay_i_23__N_1202[4] ;
    output \dout_i_23__N_5777[4] ;
    input \op_i_23__N_1154[3] ;
    input \delay_i_23__N_1202[3] ;
    output \dout_i_23__N_5777[3] ;
    input \op_i_23__N_1154[22] ;
    input \delay_i_23__N_1202[22] ;
    output \dout_i_23__N_5777[22] ;
    input \op_r_23__N_1106[7] ;
    input \delay_r_23__N_1178[7] ;
    output \dout_r_23__N_5681[7] ;
    input \op_r_23__N_1106[6] ;
    input \delay_r_23__N_1178[6] ;
    output \dout_r_23__N_5681[6] ;
    input \op_r_23__N_1106[5] ;
    input \delay_r_23__N_1178[5] ;
    output \dout_r_23__N_5681[5] ;
    input \op_r_23__N_1106[4] ;
    input \delay_r_23__N_1178[4] ;
    output \dout_r_23__N_5681[4] ;
    input \op_r_23__N_1106[17] ;
    input \delay_r_23__N_1178[17] ;
    output \dout_r_23__N_5681[17] ;
    input \op_r_23__N_1106[3] ;
    input \delay_r_23__N_1178[3] ;
    output \dout_r_23__N_5681[3] ;
    input \op_r_23__N_1106[2] ;
    input \delay_r_23__N_1178[2] ;
    output \dout_r_23__N_5681[2] ;
    input \op_r_23__N_1106[16] ;
    input \delay_r_23__N_1178[16] ;
    output \dout_r_23__N_5681[16] ;
    input \op_r_23__N_1106[1] ;
    input \delay_r_23__N_1178[1] ;
    output \dout_r_23__N_5681[1] ;
    input \op_i_23__N_1154[15] ;
    input \delay_i_23__N_1202[15] ;
    output \dout_i_23__N_5777[15] ;
    input \op_i_23__N_1154[14] ;
    input \delay_i_23__N_1202[14] ;
    output \dout_i_23__N_5777[14] ;
    
    
    wire n15814, n15815, n15816, n15817, n15818, n15819, n15820, 
        n15821, n15822, n15823, n15824, n15825, n15826, n15827, 
        n15828, n15829, n15830, n15831, n15832, n15833, n15834, 
        n15835, n15836, n15837, n15838, n15839, n15840, n15841, 
        n15842, n15843, n15844, n15845, n15846, n15847, n15848, 
        n15849, n15850, n15851, n15852, n15853, n15854, n15855, 
        n15856, n15857, n15858, n15859, n15860, n15861, n15862, 
        n15863, n15864, n15865, n15866, n15867, n15868, n15869, 
        n15870, n15871, n15872, n15873, n15874, n15875, n15876, 
        n15877, n15878, n15879, n15880, n15881, n15882, n15883, 
        n15884, n15885, n15886, n15887, n15888, n15889, n15890, 
        n15891, n15892, n15893, n15894, n15895, n15896, n15897, 
        n15898, n15899, n15900, n15901, n15902, n15903, n15904, 
        n15905, n15906, n15907, n15908, n15909, n15910, n15911, 
        n15912, n15913, n15914, n15915, n15916, n15917, n15918, 
        n15919, n15920, n15921, n15922, n15923, n15924, n15925, 
        n15926, n15927, n15928, n15929, n15930, n15931, n15932, 
        n15933, n15934, n15935, n15936, n15937, n15938, n15939, 
        n15940, n15941, n15942, n15943, n15944, n15945, n15946, 
        n15947, n15948, n15949, n15950, n15951, n15952, n15953, 
        n15954, n15955, n15956, n15957, n15958, n15959, n15960, 
        n15961, n15962, n15963, n15964, n15965, n15966, n15967, 
        n15968, n15969, n15970, n15971, n15972, n15973, n15974, 
        n15975, n15976, n15977, n15978, n15979, n15980, n15981, 
        n15982, n15983, n15984, n15985, n15986, n15987, n15988, 
        n15989, n15990, n15991, n15992, n15993, n15994, n15995, 
        n15996, n15668, n15669, n15670, n15671, n15672, n15673, 
        n15674, n15675, n15676, n15677, n15678, n15679, n15680, 
        n15681, n15682, n15683, n15684, n15685, n15686, n15687, 
        n15688, n15689, n15690, n15691, n15692, n15693, n15694, 
        n15695, n15696, n15697, n15698, n15699, n15700, n15701, 
        n15702, n15703, n15704, n15705, n15706, n15707, n15708, 
        n15709, n15710, n15711, n15712, n15713, n15714, n15715, 
        n15716, n15717, n15718, n15719, n15720, n15721, n15722, 
        n15723, n15724, n15725, n15726, n15727, n15728, n15729, 
        n15730, n15731, n15732, n15733, n15734, n15735, n15736, 
        n15737, n15738, n15739, n15740, n15741, n15742, n15743, 
        n15744, n15745, n15746, n15747, n15748, n15749, n15750, 
        n15751, n15752, n15753, n15754, n15755, n15756, n15757, 
        n15758, n15759, n15760, n15761, n15762, n15763, n15764, 
        n15765, n15766, n15767, n15768, n15769, n15770, n15771, 
        n15772, n15773, n15774, n15775, n15776, n15777, n15778, 
        n15779, n15780, n15781, n15782, n15783, n15784, n15785, 
        n15786, n15787, n15788, n15789, n15790, n15791, n15792, 
        n15793, n15794, n15795, n15796, n15797, n15798, n15799, 
        n15800, n15801, n15802, n15803, n15804, n15805, n15806, 
        n15807, n15808, n15809, n15810, n15811, n15812, n15813, 
        mult_24s_7s_0_mult_4_11_n2, n16579, n16580, n16581, n16582, 
        n16583, n16584, n16585, n16586, n16587, n16588, n16589, 
        n16590, n16591, n16592, n16593, n16594, n16595, n16596, 
        n16597, n16598, n16599, n16600, n16601, n16602, n16603, 
        n16604, n16605, n16606, n16607, n16608, n16609, n16610, 
        n16611, n16612, n16613, n16614, n16615, n16616, n16617, 
        n16618, n16619, n16620, n16621, n16622, n16623, n16624, 
        n16625, n16626, n16627, n16628, n16629, n16630, n16631, 
        n16632, n16633, n16634, n16635, n16636, n16637, n16638, 
        n16639, n16640, n16641, n16642, n16643, n16644, n16645, 
        n16646, n16647, n16648, n16649, n16650, n16651, n16506, 
        n16507, n16508, n16509, n16510, n16511, n16512, n16513, 
        n16514, n16515, n16516, n16517, n16518, n16519, n16520, 
        n16521, n16522, n16523, n16524, n16525, n16526, n16527, 
        n16528, n16529, n16530, n16531, n16532, n16533, n16534, 
        n16535, n16536, n16537, n16538, n16539, n16540, n16541, 
        n16542, n16543, n16544, n16545, n16546, n16547, n16548, 
        n16549, n16550, n16551, n16552, n16553, n16554, n16555, 
        n16556, n16557, n16558, n16559, n16560, n16561, n16562, 
        n16563, n16564, n16565, n16566, n16567, n16568, n16569, 
        n16570, n16571, n16572, n16573, n16574, n16575, n16576, 
        n16577, n16578, n16652, n16653, n16654, n16655, n16656, 
        n16657, n16658, n16659, n16660, n16661, n16662, n16663, 
        n16664, n16665, n16666, n16667, n16668, n16669, n16670, 
        n16671, n16672, n16673, n16674, n16675, n16676, n16677, 
        n16678, n16679, n16680, n16681, n16682, n16683, n16684, 
        n16685, n16686, n16687, n16688, n14413, n14414, n14415, 
        n14416, n14417, n14418, n14419, n14420, n14421, n14422, 
        n14423, n14424, n14425, n14426, n14427, n14428, n14429, 
        n14430, n14431, n14432, n14433, n14434, n14435, n14436, 
        n14437, n14438, n14439, n14440, n14441, n14442, n14443, 
        n14444, n14445, n14446, n14447, n14448, n14449, n14450, 
        n14451, n14452, n14453, n14454, n14455, n14456, n14457, 
        n14458, n14459, n14460, n14461, n14462, n14463, n14464, 
        n14465, n14466, n14467, n14468, n14469, n14470, n14471, 
        n14472, n14473, n14474, n14475, n14476, n14477, n14478, 
        n14479, n14480, n14481, n14482, n14483, n14484, n14485, 
        n14486, n14487, n14488, n14489, n14490, n14491, n14492, 
        n14493, n14494, n14495, n14496, n14497, n14498, n14499, 
        n14500, n14501, n14502, n14503, n14504, n14505, n14506, 
        n14507, n14508, n14509, n14510, n14511, n14512, n14513, 
        n14514, n14515, n14516, n14517, n14518, n14519, n14520, 
        n14521, n14522, n14523, n14524, n14525, n14526, n14527, 
        n14528, n14529, n14530, n14531, n14532, n14533, n14534, 
        n14535, n14536, n14537, n14538, n14539, n14540, n14541, 
        n14542, n14543, n14544, n14545, n14546, n14547, n14548, 
        n14549, n14550, n14551, n14552, n14553, n14554, n14555, 
        n14556, n14557, n14558, n14559, n14560, n14561, n14562, 
        n14563, n14564, n14565, n14566, n14567, n14568, n14569, 
        n14570, n14571, n14572, n14573, n14574, n14575, n14576, 
        n14577, n14578, n14579, n14580, n14581, n14582, n14583, 
        n14584, n14585, n14586, n14587, n14588, n14589, n14590, 
        n14591, n14592, n14593, n14594, n14595, n14267, n14268, 
        n14269, n14270, n14271, n14272, n14273, n14274, n14275, 
        n14276, n14277, n14278, n14279, n14280, n14281, n14282, 
        n14283, n14284, n14285, n14286, n14287, n14288, n14289, 
        n14290, n14291, n14292, n14293, n14294, n14295, n14296, 
        n14297, n14298, n14299, n14300, n14301, n14302, n14303, 
        n14304, n14305, n14306, n14307, n14308, n14309, n14310, 
        n14311, n14312, n14313, n14314, n14315, n14316, n14317, 
        n14318, n14319, n14320, n14321, n14322, n14323, n14324, 
        n14325, n14326, n14327, n14328, n14329, n14330, n14331, 
        n14332, n14333, n14334, n14335, n14336, n14337, n14338, 
        n14339, n14340, n14341, n14342, n14343, n14344, n14345, 
        n14346, n14347, n14348, n14349, n14350, n14351, n14352, 
        n14353, n14354, n14355, n14356, n14357, n14358, n14359, 
        n14360, n14361, n14362, n14363, n14364, n14365, n14366, 
        n14367, n14368, n14369, n14370, n14371, n14372, n14373, 
        n14374, n14375, n14376, n14377, n14378, n14379, n14380, 
        n14381, n14382, n14383, n14384, n14385, n14386, n14387, 
        n14388, n14389, n14390, n14391, n14392, n14393, n14394, 
        n14395, n14396, n14397, n14398, n14399, n14400, n14401, 
        n14402, n14403, n14404, n14405, n14406, n14407, n14408, 
        n14409, n14410, n14411, n14412, mult_24s_7s_0_mult_4_11_n2_adj_6032, 
        n16360, n16361, n16362, n16363, n16364, n16365, n16366, 
        n16367, n16368, n16369, n16370, n16371, n16372, n16373, 
        n16374, n16375, n16376, n16377, n16378, n16379, n16380, 
        n16381, n16382, n16383, n16384, n16385, n16386, n16387, 
        n16388, n16389, n16390, n16391, n16392, n16393, n16394, 
        n16395, n16396, n16397, n16398, n16399, n16400, n16401, 
        n16402, n16403, n16404, n16405, n16406, n16407, n16408, 
        n16409, n16410, n16411, n16412, n16413, n16414, n16415, 
        n16416, n16417, n16418, n16419, n16420, n16421, n16422, 
        n16423, n16424, n16425, n16426, n16427, n16428, n16429, 
        n16430, n16431, n16432, n16433, n16434, n16435, n16436, 
        n16437, n16438, n16439, n16440, n16441, n16442, n16443, 
        n16444, n16445, n16446, n16447, n16448, n16449, n16450, 
        n16451, n16452, n16453, n16454, n16455, n16456, n16457, 
        n16458, n16459, n16460, n16461, n16462, n16463, n16464, 
        n16465, n16466, n16467, n16468, n16469, n16470, n16471, 
        n16472, n16473, n16474, n16475, n16476, n16477, n16478, 
        n16479, n16480, n16481, n16482, n16483, n16484, n16485, 
        n16486, n16487, n16488, n16489, n16490, n16491, n16492, 
        n16493, n16494, n16495, n16496, n16497, n16498, n16499, 
        n16500, n16501, n16502, n16503, n16504, n16505, mult_24s_7s_0_mult_2_11_n2, 
        mult_24s_7s_0_mult_0_11_n3, mult_24s_7s_0_mult_0_11_n1, mult_24s_7s_0_pp_1_2, 
        mult_24s_7s_0_mult_2_11_n1, mult_24s_7s_0_pp_2_4, mult_24s_7s_0_mult_4_11_n1, 
        mult_24s_7s_0_pp_3_6, mult_24s_7s_0_pp_3_7, mult_24s_7s_0_pp_3_8, 
        mult_24s_7s_0_pp_3_9, mult_24s_7s_0_pp_3_10, mult_24s_7s_0_pp_3_11, 
        mult_24s_7s_0_pp_3_12, mult_24s_7s_0_pp_3_13, mult_24s_7s_0_pp_3_14, 
        mult_24s_7s_0_pp_3_15, mult_24s_7s_0_pp_3_16, mult_24s_7s_0_pp_3_17, 
        mult_24s_7s_0_pp_3_18, mult_24s_7s_0_pp_3_19, mult_24s_7s_0_pp_3_20, 
        mult_24s_7s_0_pp_3_21, mult_24s_7s_0_pp_3_22, mult_24s_7s_0_pp_3_23, 
        mult_24s_7s_0_pp_3_24, mult_24s_7s_0_pp_3_25, mult_24s_7s_0_pp_3_26, 
        mult_24s_7s_0_pp_3_27, mult_24s_7s_0_pp_3_28, mult_24s_7s_0_pp_3_29, 
        mult_24s_7s_0_pp_0_25, mfco, mult_24s_7s_0_cin_lr_2, mult_24s_7s_0_pp_1_27, 
        mfco_1, mult_24s_7s_0_cin_lr_4, mult_24s_7s_0_pp_2_29, mfco_2, 
        co_mult_24s_7s_0_0_1, mult_24s_7s_0_pp_0_2, co_mult_24s_7s_0_0_2, 
        s_mult_24s_7s_0_0_4, mult_24s_7s_0_pp_0_4, mult_24s_7s_0_pp_0_3, 
        mult_24s_7s_0_pp_1_4, mult_24s_7s_0_pp_1_3, co_mult_24s_7s_0_0_3, 
        s_mult_24s_7s_0_0_6, s_mult_24s_7s_0_0_5, mult_24s_7s_0_pp_0_6, 
        mult_24s_7s_0_pp_0_5, mult_24s_7s_0_pp_1_6, mult_24s_7s_0_pp_1_5, 
        co_mult_24s_7s_0_0_4, s_mult_24s_7s_0_0_8, s_mult_24s_7s_0_0_7, 
        mult_24s_7s_0_pp_0_8, mult_24s_7s_0_pp_0_7, mult_24s_7s_0_pp_1_8, 
        mult_24s_7s_0_pp_1_7, co_mult_24s_7s_0_0_5, s_mult_24s_7s_0_0_10, 
        s_mult_24s_7s_0_0_9, mult_24s_7s_0_pp_0_10, mult_24s_7s_0_pp_0_9, 
        mult_24s_7s_0_pp_1_10, mult_24s_7s_0_pp_1_9, co_mult_24s_7s_0_0_6, 
        s_mult_24s_7s_0_0_12, s_mult_24s_7s_0_0_11, mult_24s_7s_0_pp_0_12, 
        mult_24s_7s_0_pp_0_11, mult_24s_7s_0_pp_1_12, mult_24s_7s_0_pp_1_11, 
        co_mult_24s_7s_0_0_7, s_mult_24s_7s_0_0_14, s_mult_24s_7s_0_0_13, 
        mult_24s_7s_0_pp_0_14, mult_24s_7s_0_pp_0_13, mult_24s_7s_0_pp_1_14, 
        mult_24s_7s_0_pp_1_13, co_mult_24s_7s_0_0_8, s_mult_24s_7s_0_0_16, 
        s_mult_24s_7s_0_0_15, mult_24s_7s_0_pp_0_16, mult_24s_7s_0_pp_0_15, 
        mult_24s_7s_0_pp_1_16, mult_24s_7s_0_pp_1_15, co_mult_24s_7s_0_0_9, 
        s_mult_24s_7s_0_0_18, s_mult_24s_7s_0_0_17, mult_24s_7s_0_pp_0_18, 
        mult_24s_7s_0_pp_0_17, mult_24s_7s_0_pp_1_18, mult_24s_7s_0_pp_1_17, 
        co_mult_24s_7s_0_0_10, s_mult_24s_7s_0_0_20, s_mult_24s_7s_0_0_19, 
        mult_24s_7s_0_pp_0_20, mult_24s_7s_0_pp_0_19, mult_24s_7s_0_pp_1_20, 
        mult_24s_7s_0_pp_1_19, co_mult_24s_7s_0_0_11, s_mult_24s_7s_0_0_22, 
        s_mult_24s_7s_0_0_21, mult_24s_7s_0_pp_0_22, mult_24s_7s_0_pp_0_21, 
        mult_24s_7s_0_pp_1_22, mult_24s_7s_0_pp_1_21, co_mult_24s_7s_0_0_12, 
        s_mult_24s_7s_0_0_24, s_mult_24s_7s_0_0_23, mult_24s_7s_0_pp_0_24, 
        mult_24s_7s_0_pp_0_23, mult_24s_7s_0_pp_1_24, mult_24s_7s_0_pp_1_23, 
        co_mult_24s_7s_0_0_13, s_mult_24s_7s_0_0_26, s_mult_24s_7s_0_0_25, 
        mult_24s_7s_0_pp_1_26, mult_24s_7s_0_pp_1_25, co_mult_24s_7s_0_0_14, 
        s_mult_24s_7s_0_0_28, s_mult_24s_7s_0_0_27, s_mult_24s_7s_0_0_29, 
        co_mult_24s_7s_0_1_1, s_mult_24s_7s_0_1_6, mult_24s_7s_0_pp_2_6, 
        co_mult_24s_7s_0_1_2, s_mult_24s_7s_0_1_8, s_mult_24s_7s_0_1_7, 
        mult_24s_7s_0_pp_2_8, mult_24s_7s_0_pp_2_7, co_mult_24s_7s_0_1_3, 
        s_mult_24s_7s_0_1_10, s_mult_24s_7s_0_1_9, mult_24s_7s_0_pp_2_10, 
        mult_24s_7s_0_pp_2_9, co_mult_24s_7s_0_1_4, s_mult_24s_7s_0_1_12, 
        s_mult_24s_7s_0_1_11, mult_24s_7s_0_pp_2_12, mult_24s_7s_0_pp_2_11, 
        co_mult_24s_7s_0_1_5, s_mult_24s_7s_0_1_14, s_mult_24s_7s_0_1_13, 
        mult_24s_7s_0_pp_2_14, mult_24s_7s_0_pp_2_13, co_mult_24s_7s_0_1_6, 
        s_mult_24s_7s_0_1_16, s_mult_24s_7s_0_1_15, mult_24s_7s_0_pp_2_16, 
        mult_24s_7s_0_pp_2_15, co_mult_24s_7s_0_1_7, s_mult_24s_7s_0_1_18, 
        s_mult_24s_7s_0_1_17, mult_24s_7s_0_pp_2_18, mult_24s_7s_0_pp_2_17, 
        co_mult_24s_7s_0_1_8, s_mult_24s_7s_0_1_20, s_mult_24s_7s_0_1_19, 
        mult_24s_7s_0_pp_2_20, mult_24s_7s_0_pp_2_19, co_mult_24s_7s_0_1_9, 
        s_mult_24s_7s_0_1_22, s_mult_24s_7s_0_1_21, mult_24s_7s_0_pp_2_22, 
        mult_24s_7s_0_pp_2_21, co_mult_24s_7s_0_1_10, s_mult_24s_7s_0_1_24, 
        s_mult_24s_7s_0_1_23, mult_24s_7s_0_pp_2_24, mult_24s_7s_0_pp_2_23, 
        co_mult_24s_7s_0_1_11, s_mult_24s_7s_0_1_26, s_mult_24s_7s_0_1_25, 
        mult_24s_7s_0_pp_2_26, mult_24s_7s_0_pp_2_25, co_mult_24s_7s_0_1_12, 
        s_mult_24s_7s_0_1_28, s_mult_24s_7s_0_1_27, mult_24s_7s_0_pp_2_28, 
        mult_24s_7s_0_pp_2_27, s_mult_24s_7s_0_1_30, s_mult_24s_7s_0_1_29, 
        co_mult_24s_7s_0_2_1, co_mult_24s_7s_0_2_2, s_mult_24s_7s_0_2_6, 
        mult_24s_7s_0_pp_2_5, co_mult_24s_7s_0_2_3, s_mult_24s_7s_0_2_8, 
        s_mult_24s_7s_0_2_7, co_mult_24s_7s_0_2_4, s_mult_24s_7s_0_2_10, 
        s_mult_24s_7s_0_2_9, co_mult_24s_7s_0_2_5, s_mult_24s_7s_0_2_12, 
        s_mult_24s_7s_0_2_11, co_mult_24s_7s_0_2_6, s_mult_24s_7s_0_2_14, 
        s_mult_24s_7s_0_2_13, co_mult_24s_7s_0_2_7, s_mult_24s_7s_0_2_16, 
        s_mult_24s_7s_0_2_15, co_mult_24s_7s_0_2_8, s_mult_24s_7s_0_2_18, 
        s_mult_24s_7s_0_2_17, co_mult_24s_7s_0_2_9, s_mult_24s_7s_0_2_20, 
        s_mult_24s_7s_0_2_19, co_mult_24s_7s_0_2_10, s_mult_24s_7s_0_2_22, 
        s_mult_24s_7s_0_2_21, co_mult_24s_7s_0_2_11, s_mult_24s_7s_0_2_24, 
        s_mult_24s_7s_0_2_23, co_mult_24s_7s_0_2_12, s_mult_24s_7s_0_2_26, 
        s_mult_24s_7s_0_2_25, co_mult_24s_7s_0_2_13, s_mult_24s_7s_0_2_28, 
        s_mult_24s_7s_0_2_27, s_mult_24s_7s_0_2_30, s_mult_24s_7s_0_2_29, 
        co_t_mult_24s_7s_0_3_1, co_t_mult_24s_7s_0_3_2, co_t_mult_24s_7s_0_3_3, 
        co_t_mult_24s_7s_0_3_4, co_t_mult_24s_7s_0_3_5, co_t_mult_24s_7s_0_3_6, 
        co_t_mult_24s_7s_0_3_7, co_t_mult_24s_7s_0_3_8, co_t_mult_24s_7s_0_3_9, 
        co_t_mult_24s_7s_0_3_10, co_t_mult_24s_7s_0_3_11, co_t_mult_24s_7s_0_3_12, 
        mult_24s_7s_0_cin_lr_0, mco, mco_1, mco_2, mco_3, mco_4, 
        mco_5, mco_6, mco_7, mco_8, mco_9, mco_10, mco_11, mco_12, 
        mco_13, mco_14, mco_15, mco_16, mco_17, mco_18, mco_19, 
        mco_20, mco_21, mco_22, mco_23, mco_24, mco_25, mco_26, 
        mco_27, mco_28, mco_29, mco_30, mco_31, mco_32, mult_24s_7s_0_mult_2_11_n2_adj_6034, 
        mult_24s_7s_0_mult_0_11_n3_adj_6036, mult_24s_7s_0_mult_0_11_n1_adj_6039, 
        mult_24s_7s_0_pp_1_2_adj_6040, mult_24s_7s_0_mult_2_11_n1_adj_6042, 
        mult_24s_7s_0_pp_2_4_adj_6043, mult_24s_7s_0_mult_4_11_n1_adj_6045, 
        mult_24s_7s_0_pp_3_6_adj_6046, mult_24s_7s_0_pp_3_7_adj_6047, mult_24s_7s_0_pp_3_8_adj_6048, 
        mult_24s_7s_0_pp_3_9_adj_6049, mult_24s_7s_0_pp_3_10_adj_6050, mult_24s_7s_0_pp_3_11_adj_6051, 
        mult_24s_7s_0_pp_3_12_adj_6052, mult_24s_7s_0_pp_3_13_adj_6053, 
        mult_24s_7s_0_pp_3_14_adj_6054, mult_24s_7s_0_pp_3_15_adj_6055, 
        mult_24s_7s_0_pp_3_16_adj_6056, mult_24s_7s_0_pp_3_17_adj_6057, 
        mult_24s_7s_0_pp_3_18_adj_6058, mult_24s_7s_0_pp_3_19_adj_6059, 
        mult_24s_7s_0_pp_3_20_adj_6060, mult_24s_7s_0_pp_3_21_adj_6061, 
        mult_24s_7s_0_pp_3_22_adj_6062, mult_24s_7s_0_pp_3_23_adj_6063, 
        mult_24s_7s_0_pp_3_24_adj_6064, mult_24s_7s_0_pp_3_25_adj_6065, 
        mult_24s_7s_0_pp_3_26_adj_6066, mult_24s_7s_0_pp_3_27_adj_6067, 
        mult_24s_7s_0_pp_3_28_adj_6068, mult_24s_7s_0_pp_3_29_adj_6069, 
        mult_24s_7s_0_pp_0_25_adj_6070, mfco_adj_6071, mult_24s_7s_0_cin_lr_2_adj_6072, 
        mult_24s_7s_0_pp_1_27_adj_6073, mfco_1_adj_6074, mult_24s_7s_0_cin_lr_4_adj_6075, 
        mult_24s_7s_0_pp_2_29_adj_6076, mfco_2_adj_6077, co_mult_24s_7s_0_0_1_adj_6079, 
        mult_24s_7s_0_pp_0_2_adj_6080, co_mult_24s_7s_0_0_2_adj_6082, s_mult_24s_7s_0_0_4_adj_6083, 
        mult_24s_7s_0_pp_0_4_adj_6084, mult_24s_7s_0_pp_0_3_adj_6085, mult_24s_7s_0_pp_1_4_adj_6086, 
        mult_24s_7s_0_pp_1_3_adj_6087, co_mult_24s_7s_0_0_3_adj_6088, s_mult_24s_7s_0_0_6_adj_6089, 
        s_mult_24s_7s_0_0_5_adj_6090, mult_24s_7s_0_pp_0_6_adj_6091, mult_24s_7s_0_pp_0_5_adj_6092, 
        mult_24s_7s_0_pp_1_6_adj_6093, mult_24s_7s_0_pp_1_5_adj_6094, co_mult_24s_7s_0_0_4_adj_6095, 
        s_mult_24s_7s_0_0_8_adj_6096, s_mult_24s_7s_0_0_7_adj_6097, mult_24s_7s_0_pp_0_8_adj_6098, 
        mult_24s_7s_0_pp_0_7_adj_6099, mult_24s_7s_0_pp_1_8_adj_6100, mult_24s_7s_0_pp_1_7_adj_6101, 
        co_mult_24s_7s_0_0_5_adj_6102, s_mult_24s_7s_0_0_10_adj_6103, s_mult_24s_7s_0_0_9_adj_6104, 
        mult_24s_7s_0_pp_0_10_adj_6105, mult_24s_7s_0_pp_0_9_adj_6106, mult_24s_7s_0_pp_1_10_adj_6107, 
        mult_24s_7s_0_pp_1_9_adj_6108, co_mult_24s_7s_0_0_6_adj_6109, s_mult_24s_7s_0_0_12_adj_6110, 
        s_mult_24s_7s_0_0_11_adj_6111, mult_24s_7s_0_pp_0_12_adj_6112, mult_24s_7s_0_pp_0_11_adj_6113, 
        mult_24s_7s_0_pp_1_12_adj_6114, mult_24s_7s_0_pp_1_11_adj_6115, 
        co_mult_24s_7s_0_0_7_adj_6116, s_mult_24s_7s_0_0_14_adj_6117, s_mult_24s_7s_0_0_13_adj_6118, 
        mult_24s_7s_0_pp_0_14_adj_6119, mult_24s_7s_0_pp_0_13_adj_6120, 
        mult_24s_7s_0_pp_1_14_adj_6121, mult_24s_7s_0_pp_1_13_adj_6122, 
        co_mult_24s_7s_0_0_8_adj_6123, s_mult_24s_7s_0_0_16_adj_6124, s_mult_24s_7s_0_0_15_adj_6125, 
        mult_24s_7s_0_pp_0_16_adj_6126, mult_24s_7s_0_pp_0_15_adj_6127, 
        mult_24s_7s_0_pp_1_16_adj_6128, mult_24s_7s_0_pp_1_15_adj_6129, 
        co_mult_24s_7s_0_0_9_adj_6130, s_mult_24s_7s_0_0_18_adj_6131, s_mult_24s_7s_0_0_17_adj_6132, 
        mult_24s_7s_0_pp_0_18_adj_6133, mult_24s_7s_0_pp_0_17_adj_6134, 
        mult_24s_7s_0_pp_1_18_adj_6135, mult_24s_7s_0_pp_1_17_adj_6136, 
        co_mult_24s_7s_0_0_10_adj_6137, s_mult_24s_7s_0_0_20_adj_6138, s_mult_24s_7s_0_0_19_adj_6139, 
        mult_24s_7s_0_pp_0_20_adj_6140, mult_24s_7s_0_pp_0_19_adj_6141, 
        mult_24s_7s_0_pp_1_20_adj_6142, mult_24s_7s_0_pp_1_19_adj_6143, 
        co_mult_24s_7s_0_0_11_adj_6144, s_mult_24s_7s_0_0_22_adj_6145, s_mult_24s_7s_0_0_21_adj_6146, 
        mult_24s_7s_0_pp_0_22_adj_6147, mult_24s_7s_0_pp_0_21_adj_6148, 
        mult_24s_7s_0_pp_1_22_adj_6149, mult_24s_7s_0_pp_1_21_adj_6150, 
        co_mult_24s_7s_0_0_12_adj_6151, s_mult_24s_7s_0_0_24_adj_6152, s_mult_24s_7s_0_0_23_adj_6153, 
        mult_24s_7s_0_pp_0_24_adj_6154, mult_24s_7s_0_pp_0_23_adj_6155, 
        mult_24s_7s_0_pp_1_24_adj_6156, mult_24s_7s_0_pp_1_23_adj_6157, 
        co_mult_24s_7s_0_0_13_adj_6158, s_mult_24s_7s_0_0_26_adj_6159, s_mult_24s_7s_0_0_25_adj_6160, 
        mult_24s_7s_0_pp_1_26_adj_6161, mult_24s_7s_0_pp_1_25_adj_6162, 
        co_mult_24s_7s_0_0_14_adj_6163, s_mult_24s_7s_0_0_28_adj_6164, s_mult_24s_7s_0_0_27_adj_6165, 
        s_mult_24s_7s_0_0_29_adj_6166, co_mult_24s_7s_0_1_1_adj_6167, s_mult_24s_7s_0_1_6_adj_6168, 
        mult_24s_7s_0_pp_2_6_adj_6169, co_mult_24s_7s_0_1_2_adj_6170, s_mult_24s_7s_0_1_8_adj_6171, 
        s_mult_24s_7s_0_1_7_adj_6172, mult_24s_7s_0_pp_2_8_adj_6173, mult_24s_7s_0_pp_2_7_adj_6174, 
        co_mult_24s_7s_0_1_3_adj_6175, s_mult_24s_7s_0_1_10_adj_6176, s_mult_24s_7s_0_1_9_adj_6177, 
        mult_24s_7s_0_pp_2_10_adj_6178, mult_24s_7s_0_pp_2_9_adj_6179, co_mult_24s_7s_0_1_4_adj_6180, 
        s_mult_24s_7s_0_1_12_adj_6181, s_mult_24s_7s_0_1_11_adj_6182, mult_24s_7s_0_pp_2_12_adj_6183, 
        mult_24s_7s_0_pp_2_11_adj_6184, co_mult_24s_7s_0_1_5_adj_6185, s_mult_24s_7s_0_1_14_adj_6186, 
        s_mult_24s_7s_0_1_13_adj_6187, mult_24s_7s_0_pp_2_14_adj_6188, mult_24s_7s_0_pp_2_13_adj_6189, 
        co_mult_24s_7s_0_1_6_adj_6190, s_mult_24s_7s_0_1_16_adj_6191, s_mult_24s_7s_0_1_15_adj_6192, 
        mult_24s_7s_0_pp_2_16_adj_6193, mult_24s_7s_0_pp_2_15_adj_6194, 
        co_mult_24s_7s_0_1_7_adj_6195, s_mult_24s_7s_0_1_18_adj_6196, s_mult_24s_7s_0_1_17_adj_6197, 
        mult_24s_7s_0_pp_2_18_adj_6198, mult_24s_7s_0_pp_2_17_adj_6199, 
        co_mult_24s_7s_0_1_8_adj_6200, s_mult_24s_7s_0_1_20_adj_6201, s_mult_24s_7s_0_1_19_adj_6202, 
        mult_24s_7s_0_pp_2_20_adj_6203, mult_24s_7s_0_pp_2_19_adj_6204, 
        co_mult_24s_7s_0_1_9_adj_6205, s_mult_24s_7s_0_1_22_adj_6206, s_mult_24s_7s_0_1_21_adj_6207, 
        mult_24s_7s_0_pp_2_22_adj_6208, mult_24s_7s_0_pp_2_21_adj_6209, 
        co_mult_24s_7s_0_1_10_adj_6210, s_mult_24s_7s_0_1_24_adj_6211, s_mult_24s_7s_0_1_23_adj_6212, 
        mult_24s_7s_0_pp_2_24_adj_6213, mult_24s_7s_0_pp_2_23_adj_6214, 
        co_mult_24s_7s_0_1_11_adj_6215, s_mult_24s_7s_0_1_26_adj_6216, s_mult_24s_7s_0_1_25_adj_6217, 
        mult_24s_7s_0_pp_2_26_adj_6218, mult_24s_7s_0_pp_2_25_adj_6219, 
        co_mult_24s_7s_0_1_12_adj_6220, s_mult_24s_7s_0_1_28_adj_6221, s_mult_24s_7s_0_1_27_adj_6222, 
        mult_24s_7s_0_pp_2_28_adj_6223, mult_24s_7s_0_pp_2_27_adj_6224, 
        s_mult_24s_7s_0_1_30_adj_6225, s_mult_24s_7s_0_1_29_adj_6226, co_mult_24s_7s_0_2_1_adj_6228, 
        co_mult_24s_7s_0_2_2_adj_6230, s_mult_24s_7s_0_2_6_adj_6231, mult_24s_7s_0_pp_2_5_adj_6232, 
        co_mult_24s_7s_0_2_3_adj_6233, s_mult_24s_7s_0_2_8_adj_6234, s_mult_24s_7s_0_2_7_adj_6235, 
        co_mult_24s_7s_0_2_4_adj_6236, s_mult_24s_7s_0_2_10_adj_6237, s_mult_24s_7s_0_2_9_adj_6238, 
        co_mult_24s_7s_0_2_5_adj_6239, s_mult_24s_7s_0_2_12_adj_6240, s_mult_24s_7s_0_2_11_adj_6241, 
        co_mult_24s_7s_0_2_6_adj_6242, s_mult_24s_7s_0_2_14_adj_6243, s_mult_24s_7s_0_2_13_adj_6244, 
        co_mult_24s_7s_0_2_7_adj_6245, s_mult_24s_7s_0_2_16_adj_6246, s_mult_24s_7s_0_2_15_adj_6247, 
        co_mult_24s_7s_0_2_8_adj_6248, s_mult_24s_7s_0_2_18_adj_6249, s_mult_24s_7s_0_2_17_adj_6250, 
        co_mult_24s_7s_0_2_9_adj_6251, s_mult_24s_7s_0_2_20_adj_6252, s_mult_24s_7s_0_2_19_adj_6253, 
        co_mult_24s_7s_0_2_10_adj_6254, s_mult_24s_7s_0_2_22_adj_6255, s_mult_24s_7s_0_2_21_adj_6256, 
        co_mult_24s_7s_0_2_11_adj_6257, s_mult_24s_7s_0_2_24_adj_6258, s_mult_24s_7s_0_2_23_adj_6259, 
        co_mult_24s_7s_0_2_12_adj_6260, s_mult_24s_7s_0_2_26_adj_6261, s_mult_24s_7s_0_2_25_adj_6262, 
        co_mult_24s_7s_0_2_13_adj_6263, s_mult_24s_7s_0_2_28_adj_6264, s_mult_24s_7s_0_2_27_adj_6265, 
        s_mult_24s_7s_0_2_30_adj_6266, s_mult_24s_7s_0_2_29_adj_6267, co_t_mult_24s_7s_0_3_1_adj_6269, 
        co_t_mult_24s_7s_0_3_2_adj_6272, co_t_mult_24s_7s_0_3_3_adj_6275, 
        co_t_mult_24s_7s_0_3_4_adj_6278, co_t_mult_24s_7s_0_3_5_adj_6281, 
        co_t_mult_24s_7s_0_3_6_adj_6284, co_t_mult_24s_7s_0_3_7_adj_6287, 
        co_t_mult_24s_7s_0_3_8_adj_6290, co_t_mult_24s_7s_0_3_9_adj_6293, 
        co_t_mult_24s_7s_0_3_10_adj_6296, co_t_mult_24s_7s_0_3_11_adj_6299, 
        co_t_mult_24s_7s_0_3_12_adj_6302, mult_24s_7s_0_cin_lr_0_adj_6306, 
        mco_adj_6307, mco_1_adj_6308, mco_2_adj_6309, mco_3_adj_6310, 
        mco_4_adj_6311, mco_5_adj_6312, mco_6_adj_6313, mco_7_adj_6314, 
        mco_8_adj_6315, mco_9_adj_6316, mco_10_adj_6317, mco_11_adj_6318, 
        mco_12_adj_6319, mco_13_adj_6320, mco_14_adj_6321, mco_15_adj_6322, 
        mco_16_adj_6323, mco_17_adj_6324, mco_18_adj_6325, mco_19_adj_6326, 
        mco_20_adj_6327, mco_21_adj_6328, mco_22_adj_6329, mco_23_adj_6330, 
        mco_24_adj_6331, mco_25_adj_6332, mco_26_adj_6333, mco_27_adj_6334, 
        mco_28_adj_6335, mco_29_adj_6336, mco_30_adj_6337, mco_31_adj_6338, 
        mco_32_adj_6339;
    
    LUT4 i20_3_lut_4_lut (.A(\op_r_23__N_1106[14] ), .B(n34841), .C(n30179), 
         .D(\delay_r_23__N_1178[14] ), .Z(\dout_r_23__N_5681[14] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_28 (.A(\op_i_23__N_1154[13] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[13] ), .Z(\dout_i_23__N_5777[13] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_28.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_29 (.A(\op_r_23__N_1106[21] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[21] ), .Z(\dout_r_23__N_5681[21] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_29.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_30 (.A(\op_i_23__N_1154[12] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[12] ), .Z(\dout_i_23__N_5777[12] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_30.init = 16'h8f80;
    ALU54B lat_alu_39 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n15850), .SIGNEDIB(n15923), .SIGNEDCIN(n15996), .A35(n15849), 
           .A34(n15848), .A33(n15847), .A32(n15846), .A31(n15845), .A30(n15844), 
           .A29(n15843), .A28(n15842), .A27(n15841), .A26(n15840), .A25(n15839), 
           .A24(n15838), .A23(n15837), .A22(n15836), .A21(n15835), .A20(n15834), 
           .A19(n15833), .A18(n15832), .A17(n15831), .A16(n15830), .A15(n15829), 
           .A14(n15828), .A13(n15827), .A12(n15826), .A11(n15825), .A10(n15824), 
           .A9(n15823), .A8(n15822), .A7(n15821), .A6(n15820), .A5(n15819), 
           .A4(n15818), .A3(n15817), .A2(n15816), .A1(n15815), .A0(n15814), 
           .B35(n15922), .B34(n15921), .B33(n15920), .B32(n15919), .B31(n15918), 
           .B30(n15917), .B29(n15916), .B28(n15915), .B27(n15914), .B26(n15913), 
           .B25(n15912), .B24(n15911), .B23(n15910), .B22(n15909), .B21(n15908), 
           .B20(n15907), .B19(n15906), .B18(n15905), .B17(n15904), .B16(n15903), 
           .B15(n15902), .B14(n15901), .B13(n15900), .B12(n15899), .B11(n15898), 
           .B10(n15897), .B9(n15896), .B8(n15895), .B7(n15894), .B6(n15893), 
           .B5(n15892), .B4(n15891), .B3(n15890), .B2(n15889), .B1(n15888), 
           .B0(n15887), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n15886), .MA34(n15885), .MA33(n15884), .MA32(n15883), 
           .MA31(n15882), .MA30(n15881), .MA29(n15880), .MA28(n15879), 
           .MA27(n15878), .MA26(n15877), .MA25(n15876), .MA24(n15875), 
           .MA23(n15874), .MA22(n15873), .MA21(n15872), .MA20(n15871), 
           .MA19(n15870), .MA18(n15869), .MA17(n15868), .MA16(n15867), 
           .MA15(n15866), .MA14(n15865), .MA13(n15864), .MA12(n15863), 
           .MA11(n15862), .MA10(n15861), .MA9(n15860), .MA8(n15859), 
           .MA7(n15858), .MA6(n15857), .MA5(n15856), .MA4(n15855), .MA3(n15854), 
           .MA2(n15853), .MA1(n15852), .MA0(n15851), .MB35(n15959), 
           .MB34(n15958), .MB33(n15957), .MB32(n15956), .MB31(n15955), 
           .MB30(n15954), .MB29(n15953), .MB28(n15952), .MB27(n15951), 
           .MB26(n15950), .MB25(n15949), .MB24(n15948), .MB23(n15947), 
           .MB22(n15946), .MB21(n15945), .MB20(n15944), .MB19(n15943), 
           .MB18(n15942), .MB17(n15941), .MB16(n15940), .MB15(n15939), 
           .MB14(n15938), .MB13(n15937), .MB12(n15936), .MB11(n15935), 
           .MB10(n15934), .MB9(n15933), .MB8(n15932), .MB7(n15931), 
           .MB6(n15930), .MB5(n15929), .MB4(n15928), .MB3(n15927), .MB2(n15926), 
           .MB1(n15925), .MB0(n15924), .CIN53(n15995), .CIN52(n15994), 
           .CIN51(n15993), .CIN50(n15992), .CIN49(n15991), .CIN48(n15990), 
           .CIN47(n15989), .CIN46(n15988), .CIN45(n15987), .CIN44(n15986), 
           .CIN43(n15985), .CIN42(n15984), .CIN41(n15983), .CIN40(n15982), 
           .CIN39(n15981), .CIN38(n15980), .CIN37(n15979), .CIN36(n15978), 
           .CIN35(n15977), .CIN34(n15976), .CIN33(n15975), .CIN32(n15974), 
           .CIN31(n15973), .CIN30(n15972), .CIN29(n15971), .CIN28(n15970), 
           .CIN27(n15969), .CIN26(n15968), .CIN25(n15967), .CIN24(n15966), 
           .CIN23(n15965), .CIN22(n15964), .CIN21(n15963), .CIN20(n15962), 
           .CIN19(n15961), .CIN18(n15960), .CIN17(\op_r_23__N_1226[17] ), 
           .CIN16(\op_r_23__N_1226[16] ), .CIN15(\op_r_23__N_1226[15] ), 
           .CIN14(\op_r_23__N_1226[14] ), .CIN13(\op_r_23__N_1226[13] ), 
           .CIN12(\op_r_23__N_1226[12] ), .CIN11(\op_r_23__N_1226[11] ), 
           .CIN10(\op_r_23__N_1226[10] ), .CIN9(\op_r_23__N_1226[9] ), .CIN8(\op_r_23__N_1226[8] ), 
           .CIN7(\op_r_23__N_1226[7] ), .CIN6(\op_r_23__N_1226[6] ), .CIN5(\op_r_23__N_1226[5] ), 
           .CIN4(\op_r_23__N_1226[4] ), .CIN3(\op_r_23__N_1226[3] ), .CIN2(\op_r_23__N_1226[2] ), 
           .CIN1(\op_r_23__N_1226[1] ), .CIN0(\op_r_23__N_1226[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1226[31] ), 
           .R12(\op_r_23__N_1226[30] ), .R11(\op_r_23__N_1226[29] ), .R10(\op_r_23__N_1226[28] ), 
           .R9(\op_r_23__N_1226[27] ), .R8(\op_r_23__N_1226[26] ), .R7(\op_r_23__N_1226[25] ), 
           .R6(\op_r_23__N_1226[24] ), .R5(\op_r_23__N_1226[23] ), .R4(\op_r_23__N_1226[22] ), 
           .R3(\op_r_23__N_1226[21] ), .R2(\op_r_23__N_1226[20] ), .R1(\op_r_23__N_1226[19] ), 
           .R0(\op_r_23__N_1226[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_39.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_39.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_39.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_39.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_39.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_39.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_39.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_39.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_39.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_39.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_39.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_39.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_39.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_39.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_39.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_39.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_39.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_39.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_39.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_39.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_39.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_39.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_39.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_39.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_39.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_39.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_39.REG_FLAG_CLK = "NONE";
    defparam lat_alu_39.REG_FLAG_CE = "CE0";
    defparam lat_alu_39.REG_FLAG_RST = "RST0";
    defparam lat_alu_39.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_39.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_39.MASK01 = "0x00000000000000";
    defparam lat_alu_39.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_39.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_39.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_39.CLK0_DIV = "ENABLED";
    defparam lat_alu_39.CLK1_DIV = "ENABLED";
    defparam lat_alu_39.CLK2_DIV = "ENABLED";
    defparam lat_alu_39.CLK3_DIV = "ENABLED";
    defparam lat_alu_39.MCPAT = "0x00000000000000";
    defparam lat_alu_39.MASKPAT = "0x00000000000000";
    defparam lat_alu_39.RNDPAT = "0x00000000000000";
    defparam lat_alu_39.GSR = "DISABLED";
    defparam lat_alu_39.RESETMODE = "SYNC";
    defparam lat_alu_39.MULT9_MODE = "DISABLED";
    defparam lat_alu_39.LEGACY = "DISABLED";
    ALU54B lat_alu_38 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n15704), .SIGNEDIB(n15777), .SIGNEDCIN(GND_net), 
           .A35(n15703), .A34(n15702), .A33(n15701), .A32(n15700), .A31(n15699), 
           .A30(n15698), .A29(n15697), .A28(n15696), .A27(n15695), .A26(n15694), 
           .A25(n15693), .A24(n15692), .A23(n15691), .A22(n15690), .A21(n15689), 
           .A20(n15688), .A19(n15687), .A18(n15686), .A17(n15685), .A16(n15684), 
           .A15(n15683), .A14(n15682), .A13(n15681), .A12(n15680), .A11(n15679), 
           .A10(n15678), .A9(n15677), .A8(n15676), .A7(n15675), .A6(n15674), 
           .A5(n15673), .A4(n15672), .A3(n15671), .A2(n15670), .A1(n15669), 
           .A0(n15668), .B35(n15776), .B34(n15775), .B33(n15774), .B32(n15773), 
           .B31(n15772), .B30(n15771), .B29(n15770), .B28(n15769), .B27(n15768), 
           .B26(n15767), .B25(n15766), .B24(n15765), .B23(n15764), .B22(n15763), 
           .B21(n15762), .B20(n15761), .B19(n15760), .B18(n15759), .B17(n15758), 
           .B16(n15757), .B15(n15756), .B14(n15755), .B13(n15754), .B12(n15753), 
           .B11(n15752), .B10(n15751), .B9(n15750), .B8(n15749), .B7(n15748), 
           .B6(n15747), .B5(n15746), .B4(n15745), .B3(n15744), .B2(n15743), 
           .B1(n15742), .B0(n15741), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n15740), .MA34(n15739), .MA33(n15738), .MA32(n15737), 
           .MA31(n15736), .MA30(n15735), .MA29(n15734), .MA28(n15733), 
           .MA27(n15732), .MA26(n15731), .MA25(n15730), .MA24(n15729), 
           .MA23(n15728), .MA22(n15727), .MA21(n15726), .MA20(n15725), 
           .MA19(n15724), .MA18(n15723), .MA17(n15722), .MA16(n15721), 
           .MA15(n15720), .MA14(n15719), .MA13(n15718), .MA12(n15717), 
           .MA11(n15716), .MA10(n15715), .MA9(n15714), .MA8(n15713), 
           .MA7(n15712), .MA6(n15711), .MA5(n15710), .MA4(n15709), .MA3(n15708), 
           .MA2(n15707), .MA1(n15706), .MA0(n15705), .MB35(n15813), 
           .MB34(n15812), .MB33(n15811), .MB32(n15810), .MB31(n15809), 
           .MB30(n15808), .MB29(n15807), .MB28(n15806), .MB27(n15805), 
           .MB26(n15804), .MB25(n15803), .MB24(n15802), .MB23(n15801), 
           .MB22(n15800), .MB21(n15799), .MB20(n15798), .MB19(n15797), 
           .MB18(n15796), .MB17(n15795), .MB16(n15794), .MB15(n15793), 
           .MB14(n15792), .MB13(n15791), .MB12(n15790), .MB11(n15789), 
           .MB10(n15788), .MB9(n15787), .MB8(n15786), .MB7(n15785), 
           .MB6(n15784), .MB5(n15783), .MB4(n15782), .MB3(n15781), .MB2(n15780), 
           .MB1(n15779), .MB0(n15778), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n15995), 
           .R52(n15994), .R51(n15993), .R50(n15992), .R49(n15991), .R48(n15990), 
           .R47(n15989), .R46(n15988), .R45(n15987), .R44(n15986), .R43(n15985), 
           .R42(n15984), .R41(n15983), .R40(n15982), .R39(n15981), .R38(n15980), 
           .R37(n15979), .R36(n15978), .R35(n15977), .R34(n15976), .R33(n15975), 
           .R32(n15974), .R31(n15973), .R30(n15972), .R29(n15971), .R28(n15970), 
           .R27(n15969), .R26(n15968), .R25(n15967), .R24(n15966), .R23(n15965), 
           .R22(n15964), .R21(n15963), .R20(n15962), .R19(n15961), .R18(n15960), 
           .R17(\op_r_23__N_1226[17] ), .R16(\op_r_23__N_1226[16] ), .R15(\op_r_23__N_1226[15] ), 
           .R14(\op_r_23__N_1226[14] ), .R13(\op_r_23__N_1226[13] ), .R12(\op_r_23__N_1226[12] ), 
           .R11(\op_r_23__N_1226[11] ), .R10(\op_r_23__N_1226[10] ), .R9(\op_r_23__N_1226[9] ), 
           .R8(\op_r_23__N_1226[8] ), .R7(\op_r_23__N_1226[7] ), .R6(\op_r_23__N_1226[6] ), 
           .R5(\op_r_23__N_1226[5] ), .R4(\op_r_23__N_1226[4] ), .R3(\op_r_23__N_1226[3] ), 
           .R2(\op_r_23__N_1226[2] ), .R1(\op_r_23__N_1226[1] ), .R0(\op_r_23__N_1226[0] ), 
           .SIGNEDR(n15996));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_38.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_38.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_38.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_38.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_38.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_38.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_38.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_38.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_38.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_38.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_38.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_38.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_38.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_38.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_38.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_38.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_38.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_38.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_38.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_38.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_38.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_38.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_38.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_38.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_38.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_38.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_38.REG_FLAG_CLK = "NONE";
    defparam lat_alu_38.REG_FLAG_CE = "CE0";
    defparam lat_alu_38.REG_FLAG_RST = "RST0";
    defparam lat_alu_38.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_38.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_38.MASK01 = "0x00000000000000";
    defparam lat_alu_38.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_38.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_38.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_38.CLK0_DIV = "ENABLED";
    defparam lat_alu_38.CLK1_DIV = "ENABLED";
    defparam lat_alu_38.CLK2_DIV = "ENABLED";
    defparam lat_alu_38.CLK3_DIV = "ENABLED";
    defparam lat_alu_38.MCPAT = "0x00000000000000";
    defparam lat_alu_38.MASKPAT = "0x00000000000000";
    defparam lat_alu_38.RNDPAT = "0x00000000000000";
    defparam lat_alu_38.GSR = "DISABLED";
    defparam lat_alu_38.RESETMODE = "SYNC";
    defparam lat_alu_38.MULT9_MODE = "DISABLED";
    defparam lat_alu_38.LEGACY = "DISABLED";
    MULT18X18D lat_mult_37 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12176), 
            .B16(n12176), .B15(n12176), .B14(n12176), .B13(n12176), 
            .B12(n12176), .B11(n12176), .B10(n12176), .B9(n12176), .B8(n12176), 
            .B7(n12176), .B6(n12176), .B5(n12175), .B4(n12174), .B3(n12173), 
            .B2(n12172), .B1(n12171), .B0(n12170), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15904), .ROA16(n15903), .ROA15(n15902), .ROA14(n15901), 
            .ROA13(n15900), .ROA12(n15899), .ROA11(n15898), .ROA10(n15897), 
            .ROA9(n15896), .ROA8(n15895), .ROA7(n15894), .ROA6(n15893), 
            .ROA5(n15892), .ROA4(n15891), .ROA3(n15890), .ROA2(n15889), 
            .ROA1(n15888), .ROA0(n15887), .ROB17(n15922), .ROB16(n15921), 
            .ROB15(n15920), .ROB14(n15919), .ROB13(n15918), .ROB12(n15917), 
            .ROB11(n15916), .ROB10(n15915), .ROB9(n15914), .ROB8(n15913), 
            .ROB7(n15912), .ROB6(n15911), .ROB5(n15910), .ROB4(n15909), 
            .ROB3(n15908), .ROB2(n15907), .ROB1(n15906), .ROB0(n15905), 
            .P35(n15959), .P34(n15958), .P33(n15957), .P32(n15956), 
            .P31(n15955), .P30(n15954), .P29(n15953), .P28(n15952), 
            .P27(n15951), .P26(n15950), .P25(n15949), .P24(n15948), 
            .P23(n15947), .P22(n15946), .P21(n15945), .P20(n15944), 
            .P19(n15943), .P18(n15942), .P17(n15941), .P16(n15940), 
            .P15(n15939), .P14(n15938), .P13(n15937), .P12(n15936), 
            .P11(n15935), .P10(n15934), .P9(n15933), .P8(n15932), .P7(n15931), 
            .P6(n15930), .P5(n15929), .P4(n15928), .P3(n15927), .P2(n15926), 
            .P1(n15925), .P0(n15924), .SIGNEDP(n15923));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_37.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_37.REG_INPUTA_CE = "CE0";
    defparam lat_mult_37.REG_INPUTA_RST = "RST0";
    defparam lat_mult_37.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_37.REG_INPUTB_CE = "CE0";
    defparam lat_mult_37.REG_INPUTB_RST = "RST0";
    defparam lat_mult_37.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_37.REG_INPUTC_CE = "CE0";
    defparam lat_mult_37.REG_INPUTC_RST = "RST0";
    defparam lat_mult_37.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_37.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_37.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_37.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_37.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_37.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_37.CLK0_DIV = "ENABLED";
    defparam lat_mult_37.CLK1_DIV = "ENABLED";
    defparam lat_mult_37.CLK2_DIV = "ENABLED";
    defparam lat_mult_37.CLK3_DIV = "ENABLED";
    defparam lat_mult_37.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_37.GSR = "DISABLED";
    defparam lat_mult_37.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_37.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_37.MULT_BYPASS = "DISABLED";
    defparam lat_mult_37.RESETMODE = "SYNC";
    MULT18X18D lat_mult_36 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(\rom2_w_r[8] ), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12176), 
            .B16(n12176), .B15(n12176), .B14(n12176), .B13(n12176), 
            .B12(n12176), .B11(n12176), .B10(n12176), .B9(n12176), .B8(n12176), 
            .B7(n12176), .B6(n12176), .B5(n12175), .B4(n12174), .B3(n12173), 
            .B2(n12172), .B1(n12171), .B0(n12170), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15831), .ROA16(n15830), .ROA15(n15829), .ROA14(n15828), 
            .ROA13(n15827), .ROA12(n15826), .ROA11(n15825), .ROA10(n15824), 
            .ROA9(n15823), .ROA8(n15822), .ROA7(n15821), .ROA6(n15820), 
            .ROA5(n15819), .ROA4(n15818), .ROA3(n15817), .ROA2(n15816), 
            .ROA1(n15815), .ROA0(n15814), .ROB17(n15849), .ROB16(n15848), 
            .ROB15(n15847), .ROB14(n15846), .ROB13(n15845), .ROB12(n15844), 
            .ROB11(n15843), .ROB10(n15842), .ROB9(n15841), .ROB8(n15840), 
            .ROB7(n15839), .ROB6(n15838), .ROB5(n15837), .ROB4(n15836), 
            .ROB3(n15835), .ROB2(n15834), .ROB1(n15833), .ROB0(n15832), 
            .P35(n15886), .P34(n15885), .P33(n15884), .P32(n15883), 
            .P31(n15882), .P30(n15881), .P29(n15880), .P28(n15879), 
            .P27(n15878), .P26(n15877), .P25(n15876), .P24(n15875), 
            .P23(n15874), .P22(n15873), .P21(n15872), .P20(n15871), 
            .P19(n15870), .P18(n15869), .P17(n15868), .P16(n15867), 
            .P15(n15866), .P14(n15865), .P13(n15864), .P12(n15863), 
            .P11(n15862), .P10(n15861), .P9(n15860), .P8(n15859), .P7(n15858), 
            .P6(n15857), .P5(n15856), .P4(n15855), .P3(n15854), .P2(n15853), 
            .P1(n15852), .P0(n15851), .SIGNEDP(n15850));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_36.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_36.REG_INPUTA_CE = "CE0";
    defparam lat_mult_36.REG_INPUTA_RST = "RST0";
    defparam lat_mult_36.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_36.REG_INPUTB_CE = "CE0";
    defparam lat_mult_36.REG_INPUTB_RST = "RST0";
    defparam lat_mult_36.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_36.REG_INPUTC_CE = "CE0";
    defparam lat_mult_36.REG_INPUTC_RST = "RST0";
    defparam lat_mult_36.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_36.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_36.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_36.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_36.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_36.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_36.CLK0_DIV = "ENABLED";
    defparam lat_mult_36.CLK1_DIV = "ENABLED";
    defparam lat_mult_36.CLK2_DIV = "ENABLED";
    defparam lat_mult_36.CLK3_DIV = "ENABLED";
    defparam lat_mult_36.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_36.GSR = "DISABLED";
    defparam lat_mult_36.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_36.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_36.MULT_BYPASS = "DISABLED";
    defparam lat_mult_36.RESETMODE = "SYNC";
    MULT18X18D lat_mult_35 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12169), 
            .B16(n12168), .B15(n12167), .B14(n12166), .B13(n12165), 
            .B12(n12164), .B11(n12163), .B10(n12162), .B9(n12161), .B8(n12160), 
            .B7(n12159), .B6(n12158), .B5(n12157), .B4(n12156), .B3(n12155), 
            .B2(n12154), .B1(n12153), .B0(n12152), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15758), .ROA16(n15757), .ROA15(n15756), .ROA14(n15755), 
            .ROA13(n15754), .ROA12(n15753), .ROA11(n15752), .ROA10(n15751), 
            .ROA9(n15750), .ROA8(n15749), .ROA7(n15748), .ROA6(n15747), 
            .ROA5(n15746), .ROA4(n15745), .ROA3(n15744), .ROA2(n15743), 
            .ROA1(n15742), .ROA0(n15741), .ROB17(n15776), .ROB16(n15775), 
            .ROB15(n15774), .ROB14(n15773), .ROB13(n15772), .ROB12(n15771), 
            .ROB11(n15770), .ROB10(n15769), .ROB9(n15768), .ROB8(n15767), 
            .ROB7(n15766), .ROB6(n15765), .ROB5(n15764), .ROB4(n15763), 
            .ROB3(n15762), .ROB2(n15761), .ROB1(n15760), .ROB0(n15759), 
            .P35(n15813), .P34(n15812), .P33(n15811), .P32(n15810), 
            .P31(n15809), .P30(n15808), .P29(n15807), .P28(n15806), 
            .P27(n15805), .P26(n15804), .P25(n15803), .P24(n15802), 
            .P23(n15801), .P22(n15800), .P21(n15799), .P20(n15798), 
            .P19(n15797), .P18(n15796), .P17(n15795), .P16(n15794), 
            .P15(n15793), .P14(n15792), .P13(n15791), .P12(n15790), 
            .P11(n15789), .P10(n15788), .P9(n15787), .P8(n15786), .P7(n15785), 
            .P6(n15784), .P5(n15783), .P4(n15782), .P3(n15781), .P2(n15780), 
            .P1(n15779), .P0(n15778), .SIGNEDP(n15777));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_35.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_35.REG_INPUTA_CE = "CE0";
    defparam lat_mult_35.REG_INPUTA_RST = "RST0";
    defparam lat_mult_35.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_35.REG_INPUTB_CE = "CE0";
    defparam lat_mult_35.REG_INPUTB_RST = "RST0";
    defparam lat_mult_35.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_35.REG_INPUTC_CE = "CE0";
    defparam lat_mult_35.REG_INPUTC_RST = "RST0";
    defparam lat_mult_35.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_35.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_35.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_35.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_35.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_35.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_35.CLK0_DIV = "ENABLED";
    defparam lat_mult_35.CLK1_DIV = "ENABLED";
    defparam lat_mult_35.CLK2_DIV = "ENABLED";
    defparam lat_mult_35.CLK3_DIV = "ENABLED";
    defparam lat_mult_35.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_35.GSR = "DISABLED";
    defparam lat_mult_35.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_35.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_35.MULT_BYPASS = "DISABLED";
    defparam lat_mult_35.RESETMODE = "SYNC";
    MULT18X18D mult_10_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(\rom2_w_r[8] ), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12169), 
            .B16(n12168), .B15(n12167), .B14(n12166), .B13(n12165), 
            .B12(n12164), .B11(n12163), .B10(n12162), .B9(n12161), .B8(n12160), 
            .B7(n12159), .B6(n12158), .B5(n12157), .B4(n12156), .B3(n12155), 
            .B2(n12154), .B1(n12153), .B0(n12152), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15685), .ROA16(n15684), .ROA15(n15683), .ROA14(n15682), 
            .ROA13(n15681), .ROA12(n15680), .ROA11(n15679), .ROA10(n15678), 
            .ROA9(n15677), .ROA8(n15676), .ROA7(n15675), .ROA6(n15674), 
            .ROA5(n15673), .ROA4(n15672), .ROA3(n15671), .ROA2(n15670), 
            .ROA1(n15669), .ROA0(n15668), .ROB17(n15703), .ROB16(n15702), 
            .ROB15(n15701), .ROB14(n15700), .ROB13(n15699), .ROB12(n15698), 
            .ROB11(n15697), .ROB10(n15696), .ROB9(n15695), .ROB8(n15694), 
            .ROB7(n15693), .ROB6(n15692), .ROB5(n15691), .ROB4(n15690), 
            .ROB3(n15689), .ROB2(n15688), .ROB1(n15687), .ROB0(n15686), 
            .P35(n15740), .P34(n15739), .P33(n15738), .P32(n15737), 
            .P31(n15736), .P30(n15735), .P29(n15734), .P28(n15733), 
            .P27(n15732), .P26(n15731), .P25(n15730), .P24(n15729), 
            .P23(n15728), .P22(n15727), .P21(n15726), .P20(n15725), 
            .P19(n15724), .P18(n15723), .P17(n15722), .P16(n15721), 
            .P15(n15720), .P14(n15719), .P13(n15718), .P12(n15717), 
            .P11(n15716), .P10(n15715), .P9(n15714), .P8(n15713), .P7(n15712), 
            .P6(n15711), .P5(n15710), .P4(n15709), .P3(n15708), .P2(n15707), 
            .P1(n15706), .P0(n15705), .SIGNEDP(n15704));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam mult_10_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_10_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_10_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_10_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_10_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_10_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_10_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_10_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_10_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_10_mult_2.GSR = "DISABLED";
    defparam mult_10_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_10_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_10_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_10_mult_2.RESETMODE = "SYNC";
    LUT4 i20_3_lut_4_lut_adj_31 (.A(\op_r_23__N_1106[15] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[15] ), .Z(\dout_r_23__N_5681[15] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_31.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_32 (.A(\op_r_23__N_1106[13] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[13] ), .Z(\dout_r_23__N_5681[13] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_32.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_33 (.A(\op_r_23__N_1106[12] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[12] ), .Z(\dout_r_23__N_5681[12] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_33.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_34 (.A(\op_i_23__N_1154[11] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[11] ), .Z(\dout_i_23__N_5777[11] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_34.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_35 (.A(\op_r_23__N_1106[20] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[20] ), .Z(\dout_r_23__N_5681[20] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_35.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_36 (.A(\op_i_23__N_1154[10] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[10] ), .Z(\dout_i_23__N_5777[10] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_36.init = 16'h8f80;
    ND2 ND2_t25 (.A(n34795), .B(n114), .Z(mult_24s_7s_0_mult_4_11_n2)) /* synthesis syn_instantiated=1 */ ;
    MULT18X18D lat_mult_47 (.A17(shift_2_dout_i[23]), .A16(shift_2_dout_i[23]), 
            .A15(shift_2_dout_i[23]), .A14(shift_2_dout_i[23]), .A13(shift_2_dout_i[23]), 
            .A12(shift_2_dout_i[23]), .A11(shift_2_dout_i[23]), .A10(shift_2_dout_i[23]), 
            .A9(shift_2_dout_i[23]), .A8(shift_2_dout_i[23]), .A7(shift_2_dout_i[23]), 
            .A6(shift_2_dout_i[23]), .A5(shift_2_dout_i[23]), .A4(shift_2_dout_i[22]), 
            .A3(shift_2_dout_i[21]), .A2(shift_2_dout_i[20]), .A1(shift_2_dout_i[19]), 
            .A0(shift_2_dout_i[18]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(GND_net), .B7(GND_net), 
            .B6(GND_net), .B5(GND_net), .B4(GND_net), .B3(GND_net), 
            .B2(GND_net), .B1(GND_net), .B0(GND_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n16596), .ROA16(n16595), .ROA15(n16594), 
            .ROA14(n16593), .ROA13(n16592), .ROA12(n16591), .ROA11(n16590), 
            .ROA10(n16589), .ROA9(n16588), .ROA8(n16587), .ROA7(n16586), 
            .ROA6(n16585), .ROA5(n16584), .ROA4(n16583), .ROA3(n16582), 
            .ROA2(n16581), .ROA1(n16580), .ROA0(n16579), .ROB17(n16614), 
            .ROB16(n16613), .ROB15(n16612), .ROB14(n16611), .ROB13(n16610), 
            .ROB12(n16609), .ROB11(n16608), .ROB10(n16607), .ROB9(n16606), 
            .ROB8(n16605), .ROB7(n16604), .ROB6(n16603), .ROB5(n16602), 
            .ROB4(n16601), .ROB3(n16600), .ROB2(n16599), .ROB1(n16598), 
            .ROB0(n16597), .P35(n16651), .P34(n16650), .P33(n16649), 
            .P32(n16648), .P31(n16647), .P30(n16646), .P29(n16645), 
            .P28(n16644), .P27(n16643), .P26(n16642), .P25(n16641), 
            .P24(n16640), .P23(n16639), .P22(n16638), .P21(n16637), 
            .P20(n16636), .P19(n16635), .P18(n16634), .P17(n16633), 
            .P16(n16632), .P15(n16631), .P14(n16630), .P13(n16629), 
            .P12(n16628), .P11(n16627), .P10(n16626), .P9(n16625), .P8(n16624), 
            .P7(n16623), .P6(n16622), .P5(n16621), .P4(n16620), .P3(n16619), 
            .P2(n16618), .P1(n16617), .P0(n16616), .SIGNEDP(n16615));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_47.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_47.REG_INPUTA_CE = "CE0";
    defparam lat_mult_47.REG_INPUTA_RST = "RST0";
    defparam lat_mult_47.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_47.REG_INPUTB_CE = "CE0";
    defparam lat_mult_47.REG_INPUTB_RST = "RST0";
    defparam lat_mult_47.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_47.REG_INPUTC_CE = "CE0";
    defparam lat_mult_47.REG_INPUTC_RST = "RST0";
    defparam lat_mult_47.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_47.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_47.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_47.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_47.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_47.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_47.CLK0_DIV = "ENABLED";
    defparam lat_mult_47.CLK1_DIV = "ENABLED";
    defparam lat_mult_47.CLK2_DIV = "ENABLED";
    defparam lat_mult_47.CLK3_DIV = "ENABLED";
    defparam lat_mult_47.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_47.GSR = "DISABLED";
    defparam lat_mult_47.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_47.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_47.MULT_BYPASS = "DISABLED";
    defparam lat_mult_47.RESETMODE = "SYNC";
    ALU54B lat_alu_49 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n16542), .SIGNEDIB(n16615), .SIGNEDCIN(n16688), .A35(n16541), 
           .A34(n16540), .A33(n16539), .A32(n16538), .A31(n16537), .A30(n16536), 
           .A29(n16535), .A28(n16534), .A27(n16533), .A26(n16532), .A25(n16531), 
           .A24(n16530), .A23(n16529), .A22(n16528), .A21(n16527), .A20(n16526), 
           .A19(n16525), .A18(n16524), .A17(n16523), .A16(n16522), .A15(n16521), 
           .A14(n16520), .A13(n16519), .A12(n16518), .A11(n16517), .A10(n16516), 
           .A9(n16515), .A8(n16514), .A7(n16513), .A6(n16512), .A5(n16511), 
           .A4(n16510), .A3(n16509), .A2(n16508), .A1(n16507), .A0(n16506), 
           .B35(n16614), .B34(n16613), .B33(n16612), .B32(n16611), .B31(n16610), 
           .B30(n16609), .B29(n16608), .B28(n16607), .B27(n16606), .B26(n16605), 
           .B25(n16604), .B24(n16603), .B23(n16602), .B22(n16601), .B21(n16600), 
           .B20(n16599), .B19(n16598), .B18(n16597), .B17(n16596), .B16(n16595), 
           .B15(n16594), .B14(n16593), .B13(n16592), .B12(n16591), .B11(n16590), 
           .B10(n16589), .B9(n16588), .B8(n16587), .B7(n16586), .B6(n16585), 
           .B5(n16584), .B4(n16583), .B3(n16582), .B2(n16581), .B1(n16580), 
           .B0(n16579), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n16578), .MA34(n16577), .MA33(n16576), .MA32(n16575), 
           .MA31(n16574), .MA30(n16573), .MA29(n16572), .MA28(n16571), 
           .MA27(n16570), .MA26(n16569), .MA25(n16568), .MA24(n16567), 
           .MA23(n16566), .MA22(n16565), .MA21(n16564), .MA20(n16563), 
           .MA19(n16562), .MA18(n16561), .MA17(n16560), .MA16(n16559), 
           .MA15(n16558), .MA14(n16557), .MA13(n16556), .MA12(n16555), 
           .MA11(n16554), .MA10(n16553), .MA9(n16552), .MA8(n16551), 
           .MA7(n16550), .MA6(n16549), .MA5(n16548), .MA4(n16547), .MA3(n16546), 
           .MA2(n16545), .MA1(n16544), .MA0(n16543), .MB35(n16651), 
           .MB34(n16650), .MB33(n16649), .MB32(n16648), .MB31(n16647), 
           .MB30(n16646), .MB29(n16645), .MB28(n16644), .MB27(n16643), 
           .MB26(n16642), .MB25(n16641), .MB24(n16640), .MB23(n16639), 
           .MB22(n16638), .MB21(n16637), .MB20(n16636), .MB19(n16635), 
           .MB18(n16634), .MB17(n16633), .MB16(n16632), .MB15(n16631), 
           .MB14(n16630), .MB13(n16629), .MB12(n16628), .MB11(n16627), 
           .MB10(n16626), .MB9(n16625), .MB8(n16624), .MB7(n16623), 
           .MB6(n16622), .MB5(n16621), .MB4(n16620), .MB3(n16619), .MB2(n16618), 
           .MB1(n16617), .MB0(n16616), .CIN53(n16687), .CIN52(n16686), 
           .CIN51(n16685), .CIN50(n16684), .CIN49(n16683), .CIN48(n16682), 
           .CIN47(n16681), .CIN46(n16680), .CIN45(n16679), .CIN44(n16678), 
           .CIN43(n16677), .CIN42(n16676), .CIN41(n16675), .CIN40(n16674), 
           .CIN39(n16673), .CIN38(n16672), .CIN37(n16671), .CIN36(n16670), 
           .CIN35(n16669), .CIN34(n16668), .CIN33(n16667), .CIN32(n16666), 
           .CIN31(n16665), .CIN30(n16664), .CIN29(n16663), .CIN28(n16662), 
           .CIN27(n16661), .CIN26(n16660), .CIN25(n16659), .CIN24(n16658), 
           .CIN23(n16657), .CIN22(n16656), .CIN21(n16655), .CIN20(n16654), 
           .CIN19(n16653), .CIN18(n16652), .CIN17(\op_r_23__N_1268[17] ), 
           .CIN16(\op_r_23__N_1268[16] ), .CIN15(\op_r_23__N_1268[15] ), 
           .CIN14(\op_r_23__N_1268[14] ), .CIN13(\op_r_23__N_1268[13] ), 
           .CIN12(\op_r_23__N_1268[12] ), .CIN11(\op_r_23__N_1268[11] ), 
           .CIN10(\op_r_23__N_1268[10] ), .CIN9(\op_r_23__N_1268[9] ), .CIN8(\op_r_23__N_1268[8] ), 
           .CIN7(\op_r_23__N_1268[7] ), .CIN6(\op_r_23__N_1268[6] ), .CIN5(\op_r_23__N_1268[5] ), 
           .CIN4(\op_r_23__N_1268[4] ), .CIN3(\op_r_23__N_1268[3] ), .CIN2(\op_r_23__N_1268[2] ), 
           .CIN1(\op_r_23__N_1268[1] ), .CIN0(\op_r_23__N_1268[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1268[31] ), 
           .R12(\op_r_23__N_1268[30] ), .R11(\op_r_23__N_1268[29] ), .R10(\op_r_23__N_1268[28] ), 
           .R9(\op_r_23__N_1268[27] ), .R8(\op_r_23__N_1268[26] ), .R7(\op_r_23__N_1268[25] ), 
           .R6(\op_r_23__N_1268[24] ), .R5(\op_r_23__N_1268[23] ), .R4(\op_r_23__N_1268[22] ), 
           .R3(\op_r_23__N_1268[21] ), .R2(\op_r_23__N_1268[20] ), .R1(\op_r_23__N_1268[19] ), 
           .R0(\op_r_23__N_1268[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_49.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_49.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_49.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_49.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_49.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_49.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_49.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_49.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_49.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_49.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_49.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_49.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_49.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_49.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_49.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_49.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_49.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_49.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_49.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_49.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_49.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_49.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_49.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_49.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_49.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_49.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_49.REG_FLAG_CLK = "NONE";
    defparam lat_alu_49.REG_FLAG_CE = "CE0";
    defparam lat_alu_49.REG_FLAG_RST = "RST0";
    defparam lat_alu_49.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_49.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_49.MASK01 = "0x00000000000000";
    defparam lat_alu_49.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_49.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_49.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_49.CLK0_DIV = "ENABLED";
    defparam lat_alu_49.CLK1_DIV = "ENABLED";
    defparam lat_alu_49.CLK2_DIV = "ENABLED";
    defparam lat_alu_49.CLK3_DIV = "ENABLED";
    defparam lat_alu_49.MCPAT = "0x00000000000000";
    defparam lat_alu_49.MASKPAT = "0x00000000000000";
    defparam lat_alu_49.RNDPAT = "0x00000000000000";
    defparam lat_alu_49.GSR = "DISABLED";
    defparam lat_alu_49.RESETMODE = "SYNC";
    defparam lat_alu_49.MULT9_MODE = "DISABLED";
    defparam lat_alu_49.LEGACY = "DISABLED";
    ALU54B lat_alu_19 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n14449), .SIGNEDIB(n14522), .SIGNEDCIN(n14595), .A35(n14448), 
           .A34(n14447), .A33(n14446), .A32(n14445), .A31(n14444), .A30(n14443), 
           .A29(n14442), .A28(n14441), .A27(n14440), .A26(n14439), .A25(n14438), 
           .A24(n14437), .A23(n14436), .A22(n14435), .A21(n14434), .A20(n14433), 
           .A19(n14432), .A18(n14431), .A17(n14430), .A16(n14429), .A15(n14428), 
           .A14(n14427), .A13(n14426), .A12(n14425), .A11(n14424), .A10(n14423), 
           .A9(n14422), .A8(n14421), .A7(n14420), .A6(n14419), .A5(n14418), 
           .A4(n14417), .A3(n14416), .A2(n14415), .A1(n14414), .A0(n14413), 
           .B35(n14521), .B34(n14520), .B33(n14519), .B32(n14518), .B31(n14517), 
           .B30(n14516), .B29(n14515), .B28(n14514), .B27(n14513), .B26(n14512), 
           .B25(n14511), .B24(n14510), .B23(n14509), .B22(n14508), .B21(n14507), 
           .B20(n14506), .B19(n14505), .B18(n14504), .B17(n14503), .B16(n14502), 
           .B15(n14501), .B14(n14500), .B13(n14499), .B12(n14498), .B11(n14497), 
           .B10(n14496), .B9(n14495), .B8(n14494), .B7(n14493), .B6(n14492), 
           .B5(n14491), .B4(n14490), .B3(n14489), .B2(n14488), .B1(n14487), 
           .B0(n14486), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n14485), .MA34(n14484), .MA33(n14483), .MA32(n14482), 
           .MA31(n14481), .MA30(n14480), .MA29(n14479), .MA28(n14478), 
           .MA27(n14477), .MA26(n14476), .MA25(n14475), .MA24(n14474), 
           .MA23(n14473), .MA22(n14472), .MA21(n14471), .MA20(n14470), 
           .MA19(n14469), .MA18(n14468), .MA17(n14467), .MA16(n14466), 
           .MA15(n14465), .MA14(n14464), .MA13(n14463), .MA12(n14462), 
           .MA11(n14461), .MA10(n14460), .MA9(n14459), .MA8(n14458), 
           .MA7(n14457), .MA6(n14456), .MA5(n14455), .MA4(n14454), .MA3(n14453), 
           .MA2(n14452), .MA1(n14451), .MA0(n14450), .MB35(n14558), 
           .MB34(n14557), .MB33(n14556), .MB32(n14555), .MB31(n14554), 
           .MB30(n14553), .MB29(n14552), .MB28(n14551), .MB27(n14550), 
           .MB26(n14549), .MB25(n14548), .MB24(n14547), .MB23(n14546), 
           .MB22(n14545), .MB21(n14544), .MB20(n14543), .MB19(n14542), 
           .MB18(n14541), .MB17(n14540), .MB16(n14539), .MB15(n14538), 
           .MB14(n14537), .MB13(n14536), .MB12(n14535), .MB11(n14534), 
           .MB10(n14533), .MB9(n14532), .MB8(n14531), .MB7(n14530), 
           .MB6(n14529), .MB5(n14528), .MB4(n14527), .MB3(n14526), .MB2(n14525), 
           .MB1(n14524), .MB0(n14523), .CIN53(n14594), .CIN52(n14593), 
           .CIN51(n14592), .CIN50(n14591), .CIN49(n14590), .CIN48(n14589), 
           .CIN47(n14588), .CIN46(n14587), .CIN45(n14586), .CIN44(n14585), 
           .CIN43(n14584), .CIN42(n14583), .CIN41(n14582), .CIN40(n14581), 
           .CIN39(n14580), .CIN38(n14579), .CIN37(n14578), .CIN36(n14577), 
           .CIN35(n14576), .CIN34(n14575), .CIN33(n14574), .CIN32(n14573), 
           .CIN31(n14572), .CIN30(n14571), .CIN29(n14570), .CIN28(n14569), 
           .CIN27(n14568), .CIN26(n14567), .CIN25(n14566), .CIN24(n14565), 
           .CIN23(n14564), .CIN22(n14563), .CIN21(n14562), .CIN20(n14561), 
           .CIN19(n14560), .CIN18(n14559), .CIN17(n8960), .CIN16(n8961), 
           .CIN15(n8962), .CIN14(n8963), .CIN13(n8964), .CIN12(n8965), 
           .CIN11(n8966), .CIN10(n8967), .CIN9(n8968), .CIN8(n8969), 
           .CIN7(n8970), .CIN6(n8971), .CIN5(n8972), .CIN4(n8973), .CIN3(n8974), 
           .CIN2(n8975), .CIN1(n8976), .CIN0(n8977), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R7(n8952), .R6(n8953), .R5(n8954), 
           .R4(n8955), .R3(n8956), .R2(n8957), .R1(n8958), .R0(n8959));
    defparam lat_alu_19.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_19.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_19.REG_FLAG_CLK = "NONE";
    defparam lat_alu_19.REG_FLAG_CE = "CE0";
    defparam lat_alu_19.REG_FLAG_RST = "RST0";
    defparam lat_alu_19.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASK01 = "0x00000000000000";
    defparam lat_alu_19.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_19.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_19.CLK0_DIV = "ENABLED";
    defparam lat_alu_19.CLK1_DIV = "ENABLED";
    defparam lat_alu_19.CLK2_DIV = "ENABLED";
    defparam lat_alu_19.CLK3_DIV = "ENABLED";
    defparam lat_alu_19.MCPAT = "0x00000000000000";
    defparam lat_alu_19.MASKPAT = "0x00000000000000";
    defparam lat_alu_19.RNDPAT = "0x00000000000000";
    defparam lat_alu_19.GSR = "DISABLED";
    defparam lat_alu_19.RESETMODE = "SYNC";
    defparam lat_alu_19.MULT9_MODE = "DISABLED";
    defparam lat_alu_19.LEGACY = "DISABLED";
    ALU54B lat_alu_18 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n14303), .SIGNEDIB(n14376), .SIGNEDCIN(GND_net), 
           .A35(n14302), .A34(n14301), .A33(n14300), .A32(n14299), .A31(n14298), 
           .A30(n14297), .A29(n14296), .A28(n14295), .A27(n14294), .A26(n14293), 
           .A25(n14292), .A24(n14291), .A23(n14290), .A22(n14289), .A21(n14288), 
           .A20(n14287), .A19(n14286), .A18(n14285), .A17(n14284), .A16(n14283), 
           .A15(n14282), .A14(n14281), .A13(n14280), .A12(n14279), .A11(n14278), 
           .A10(n14277), .A9(n14276), .A8(n14275), .A7(n14274), .A6(n14273), 
           .A5(n14272), .A4(n14271), .A3(n14270), .A2(n14269), .A1(n14268), 
           .A0(n14267), .B35(n14375), .B34(n14374), .B33(n14373), .B32(n14372), 
           .B31(n14371), .B30(n14370), .B29(n14369), .B28(n14368), .B27(n14367), 
           .B26(n14366), .B25(n14365), .B24(n14364), .B23(n14363), .B22(n14362), 
           .B21(n14361), .B20(n14360), .B19(n14359), .B18(n14358), .B17(n14357), 
           .B16(n14356), .B15(n14355), .B14(n14354), .B13(n14353), .B12(n14352), 
           .B11(n14351), .B10(n14350), .B9(n14349), .B8(n14348), .B7(n14347), 
           .B6(n14346), .B5(n14345), .B4(n14344), .B3(n14343), .B2(n14342), 
           .B1(n14341), .B0(n14340), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n14339), .MA34(n14338), .MA33(n14337), .MA32(n14336), 
           .MA31(n14335), .MA30(n14334), .MA29(n14333), .MA28(n14332), 
           .MA27(n14331), .MA26(n14330), .MA25(n14329), .MA24(n14328), 
           .MA23(n14327), .MA22(n14326), .MA21(n14325), .MA20(n14324), 
           .MA19(n14323), .MA18(n14322), .MA17(n14321), .MA16(n14320), 
           .MA15(n14319), .MA14(n14318), .MA13(n14317), .MA12(n14316), 
           .MA11(n14315), .MA10(n14314), .MA9(n14313), .MA8(n14312), 
           .MA7(n14311), .MA6(n14310), .MA5(n14309), .MA4(n14308), .MA3(n14307), 
           .MA2(n14306), .MA1(n14305), .MA0(n14304), .MB35(n14412), 
           .MB34(n14411), .MB33(n14410), .MB32(n14409), .MB31(n14408), 
           .MB30(n14407), .MB29(n14406), .MB28(n14405), .MB27(n14404), 
           .MB26(n14403), .MB25(n14402), .MB24(n14401), .MB23(n14400), 
           .MB22(n14399), .MB21(n14398), .MB20(n14397), .MB19(n14396), 
           .MB18(n14395), .MB17(n14394), .MB16(n14393), .MB15(n14392), 
           .MB14(n14391), .MB13(n14390), .MB12(n14389), .MB11(n14388), 
           .MB10(n14387), .MB9(n14386), .MB8(n14385), .MB7(n14384), 
           .MB6(n14383), .MB5(n14382), .MB4(n14381), .MB3(n14380), .MB2(n14379), 
           .MB1(n14378), .MB0(n14377), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n14594), 
           .R52(n14593), .R51(n14592), .R50(n14591), .R49(n14590), .R48(n14589), 
           .R47(n14588), .R46(n14587), .R45(n14586), .R44(n14585), .R43(n14584), 
           .R42(n14583), .R41(n14582), .R40(n14581), .R39(n14580), .R38(n14579), 
           .R37(n14578), .R36(n14577), .R35(n14576), .R34(n14575), .R33(n14574), 
           .R32(n14573), .R31(n14572), .R30(n14571), .R29(n14570), .R28(n14569), 
           .R27(n14568), .R26(n14567), .R25(n14566), .R24(n14565), .R23(n14564), 
           .R22(n14563), .R21(n14562), .R20(n14561), .R19(n14560), .R18(n14559), 
           .R17(n8960), .R16(n8961), .R15(n8962), .R14(n8963), .R13(n8964), 
           .R12(n8965), .R11(n8966), .R10(n8967), .R9(n8968), .R8(n8969), 
           .R7(n8970), .R6(n8971), .R5(n8972), .R4(n8973), .R3(n8974), 
           .R2(n8975), .R1(n8976), .R0(n8977), .SIGNEDR(n14595));
    defparam lat_alu_18.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_18.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_18.REG_FLAG_CLK = "NONE";
    defparam lat_alu_18.REG_FLAG_CE = "CE0";
    defparam lat_alu_18.REG_FLAG_RST = "RST0";
    defparam lat_alu_18.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASK01 = "0x00000000000000";
    defparam lat_alu_18.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_18.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_18.CLK0_DIV = "ENABLED";
    defparam lat_alu_18.CLK1_DIV = "ENABLED";
    defparam lat_alu_18.CLK2_DIV = "ENABLED";
    defparam lat_alu_18.CLK3_DIV = "ENABLED";
    defparam lat_alu_18.MCPAT = "0x00000000000000";
    defparam lat_alu_18.MASKPAT = "0x00000000000000";
    defparam lat_alu_18.RNDPAT = "0x00000000000000";
    defparam lat_alu_18.GSR = "DISABLED";
    defparam lat_alu_18.RESETMODE = "SYNC";
    defparam lat_alu_18.MULT9_MODE = "DISABLED";
    defparam lat_alu_18.LEGACY = "DISABLED";
    LUT4 i20_3_lut_4_lut_adj_37 (.A(\op_i_23__N_1154[19] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[19] ), .Z(\dout_i_23__N_5777[19] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_37.init = 16'h8f80;
    MULT18X18D lat_mult_17 (.A17(n34795), .A16(n34795), .A15(n34795), 
            .A14(n34795), .A13(n34795), .A12(n34795), .A11(n34795), 
            .A10(n34795), .A9(n34795), .A8(n34795), .A7(n34795), .A6(n34795), 
            .A5(n34795), .A4(n34795), .A3(n34795), .A2(n34795), .A1(n34795), 
            .A0(n34795), .B17(n319), .B16(n319), .B15(n319), .B14(n319), 
            .B13(n319), .B12(n319), .B11(n319), .B10(n319), .B9(n319), 
            .B8(n319), .B7(n319), .B6(n319), .B5(n319), .B4(n319), 
            .B3(n319), .B2(n319), .B1(n319), .B0(n319), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n14503), .ROA16(n14502), .ROA15(n14501), 
            .ROA14(n14500), .ROA13(n14499), .ROA12(n14498), .ROA11(n14497), 
            .ROA10(n14496), .ROA9(n14495), .ROA8(n14494), .ROA7(n14493), 
            .ROA6(n14492), .ROA5(n14491), .ROA4(n14490), .ROA3(n14489), 
            .ROA2(n14488), .ROA1(n14487), .ROA0(n14486), .ROB17(n14521), 
            .ROB16(n14520), .ROB15(n14519), .ROB14(n14518), .ROB13(n14517), 
            .ROB12(n14516), .ROB11(n14515), .ROB10(n14514), .ROB9(n14513), 
            .ROB8(n14512), .ROB7(n14511), .ROB6(n14510), .ROB5(n14509), 
            .ROB4(n14508), .ROB3(n14507), .ROB2(n14506), .ROB1(n14505), 
            .ROB0(n14504), .P35(n14558), .P34(n14557), .P33(n14556), 
            .P32(n14555), .P31(n14554), .P30(n14553), .P29(n14552), 
            .P28(n14551), .P27(n14550), .P26(n14549), .P25(n14548), 
            .P24(n14547), .P23(n14546), .P22(n14545), .P21(n14544), 
            .P20(n14543), .P19(n14542), .P18(n14541), .P17(n14540), 
            .P16(n14539), .P15(n14538), .P14(n14537), .P13(n14536), 
            .P12(n14535), .P11(n14534), .P10(n14533), .P9(n14532), .P8(n14531), 
            .P7(n14530), .P6(n14529), .P5(n14528), .P4(n14527), .P3(n14526), 
            .P2(n14525), .P1(n14524), .P0(n14523), .SIGNEDP(n14522));
    defparam lat_mult_17.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTA_CE = "CE0";
    defparam lat_mult_17.REG_INPUTA_RST = "RST0";
    defparam lat_mult_17.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTB_CE = "CE0";
    defparam lat_mult_17.REG_INPUTB_RST = "RST0";
    defparam lat_mult_17.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTC_CE = "CE0";
    defparam lat_mult_17.REG_INPUTC_RST = "RST0";
    defparam lat_mult_17.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_17.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_17.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_17.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_17.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_17.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_17.CLK0_DIV = "ENABLED";
    defparam lat_mult_17.CLK1_DIV = "ENABLED";
    defparam lat_mult_17.CLK2_DIV = "ENABLED";
    defparam lat_mult_17.CLK3_DIV = "ENABLED";
    defparam lat_mult_17.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_17.GSR = "DISABLED";
    defparam lat_mult_17.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_17.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_17.MULT_BYPASS = "DISABLED";
    defparam lat_mult_17.RESETMODE = "SYNC";
    ND2 ND2_t25_adj_38 (.A(\rom4_w_i[12] ), .B(n114_adj_33), .Z(mult_24s_7s_0_mult_4_11_n2_adj_6032)) /* synthesis syn_instantiated=1 */ ;
    MULT18X18D lat_mult_16 (.A17(n34795), .A16(n34795), .A15(n34795), 
            .A14(n34795), .A13(n34795), .A12(n34795), .A11(n34795), 
            .A10(n34795), .A9(n34795), .A8(n34795), .A7(GND_net), .A6(GND_net), 
            .A5(GND_net), .A4(GND_net), .A3(GND_net), .A2(GND_net), 
            .A1(GND_net), .A0(GND_net), .B17(n319), .B16(n319), .B15(n319), 
            .B14(n319), .B13(n319), .B12(n319), .B11(n319), .B10(n319), 
            .B9(n319), .B8(n319), .B7(n319), .B6(n319), .B5(n319), 
            .B4(n319), .B3(n319), .B2(n319), .B1(n319), .B0(n319), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14430), .ROA16(n14429), 
            .ROA15(n14428), .ROA14(n14427), .ROA13(n14426), .ROA12(n14425), 
            .ROA11(n14424), .ROA10(n14423), .ROA9(n14422), .ROA8(n14421), 
            .ROA7(n14420), .ROA6(n14419), .ROA5(n14418), .ROA4(n14417), 
            .ROA3(n14416), .ROA2(n14415), .ROA1(n14414), .ROA0(n14413), 
            .ROB17(n14448), .ROB16(n14447), .ROB15(n14446), .ROB14(n14445), 
            .ROB13(n14444), .ROB12(n14443), .ROB11(n14442), .ROB10(n14441), 
            .ROB9(n14440), .ROB8(n14439), .ROB7(n14438), .ROB6(n14437), 
            .ROB5(n14436), .ROB4(n14435), .ROB3(n14434), .ROB2(n14433), 
            .ROB1(n14432), .ROB0(n14431), .P35(n14485), .P34(n14484), 
            .P33(n14483), .P32(n14482), .P31(n14481), .P30(n14480), 
            .P29(n14479), .P28(n14478), .P27(n14477), .P26(n14476), 
            .P25(n14475), .P24(n14474), .P23(n14473), .P22(n14472), 
            .P21(n14471), .P20(n14470), .P19(n14469), .P18(n14468), 
            .P17(n14467), .P16(n14466), .P15(n14465), .P14(n14464), 
            .P13(n14463), .P12(n14462), .P11(n14461), .P10(n14460), 
            .P9(n14459), .P8(n14458), .P7(n14457), .P6(n14456), .P5(n14455), 
            .P4(n14454), .P3(n14453), .P2(n14452), .P1(n14451), .P0(n14450), 
            .SIGNEDP(n14449));
    defparam lat_mult_16.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTA_CE = "CE0";
    defparam lat_mult_16.REG_INPUTA_RST = "RST0";
    defparam lat_mult_16.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTB_CE = "CE0";
    defparam lat_mult_16.REG_INPUTB_RST = "RST0";
    defparam lat_mult_16.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTC_CE = "CE0";
    defparam lat_mult_16.REG_INPUTC_RST = "RST0";
    defparam lat_mult_16.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_16.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_16.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_16.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_16.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_16.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_16.CLK0_DIV = "ENABLED";
    defparam lat_mult_16.CLK1_DIV = "ENABLED";
    defparam lat_mult_16.CLK2_DIV = "ENABLED";
    defparam lat_mult_16.CLK3_DIV = "ENABLED";
    defparam lat_mult_16.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_16.GSR = "DISABLED";
    defparam lat_mult_16.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_16.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_16.MULT_BYPASS = "DISABLED";
    defparam lat_mult_16.RESETMODE = "SYNC";
    MULT18X18D lat_mult_15 (.A17(n34795), .A16(n34795), .A15(n34795), 
            .A14(n34795), .A13(n34795), .A12(n34795), .A11(n34795), 
            .A10(n34795), .A9(n34795), .A8(n34795), .A7(n34795), .A6(n34795), 
            .A5(n34795), .A4(n34795), .A3(n34795), .A2(n34795), .A1(n34795), 
            .A0(n34795), .B17(n11143), .B16(n11142), .B15(n11141), .B14(n11140), 
            .B13(n11139), .B12(n11138), .B11(n11137), .B10(n11136), 
            .B9(n11135), .B8(n11134), .B7(n11133), .B6(n11132), .B5(n11131), 
            .B4(n11130), .B3(n11129), .B2(n11128), .B1(n11127), .B0(n11126), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14357), .ROA16(n14356), 
            .ROA15(n14355), .ROA14(n14354), .ROA13(n14353), .ROA12(n14352), 
            .ROA11(n14351), .ROA10(n14350), .ROA9(n14349), .ROA8(n14348), 
            .ROA7(n14347), .ROA6(n14346), .ROA5(n14345), .ROA4(n14344), 
            .ROA3(n14343), .ROA2(n14342), .ROA1(n14341), .ROA0(n14340), 
            .ROB17(n14375), .ROB16(n14374), .ROB15(n14373), .ROB14(n14372), 
            .ROB13(n14371), .ROB12(n14370), .ROB11(n14369), .ROB10(n14368), 
            .ROB9(n14367), .ROB8(n14366), .ROB7(n14365), .ROB6(n14364), 
            .ROB5(n14363), .ROB4(n14362), .ROB3(n14361), .ROB2(n14360), 
            .ROB1(n14359), .ROB0(n14358), .P35(n14412), .P34(n14411), 
            .P33(n14410), .P32(n14409), .P31(n14408), .P30(n14407), 
            .P29(n14406), .P28(n14405), .P27(n14404), .P26(n14403), 
            .P25(n14402), .P24(n14401), .P23(n14400), .P22(n14399), 
            .P21(n14398), .P20(n14397), .P19(n14396), .P18(n14395), 
            .P17(n14394), .P16(n14393), .P15(n14392), .P14(n14391), 
            .P13(n14390), .P12(n14389), .P11(n14388), .P10(n14387), 
            .P9(n14386), .P8(n14385), .P7(n14384), .P6(n14383), .P5(n14382), 
            .P4(n14381), .P3(n14380), .P2(n14379), .P1(n14378), .P0(n14377), 
            .SIGNEDP(n14376));
    defparam lat_mult_15.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTA_CE = "CE0";
    defparam lat_mult_15.REG_INPUTA_RST = "RST0";
    defparam lat_mult_15.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTB_CE = "CE0";
    defparam lat_mult_15.REG_INPUTB_RST = "RST0";
    defparam lat_mult_15.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTC_CE = "CE0";
    defparam lat_mult_15.REG_INPUTC_RST = "RST0";
    defparam lat_mult_15.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_15.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_15.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_15.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_15.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_15.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_15.CLK0_DIV = "ENABLED";
    defparam lat_mult_15.CLK1_DIV = "ENABLED";
    defparam lat_mult_15.CLK2_DIV = "ENABLED";
    defparam lat_mult_15.CLK3_DIV = "ENABLED";
    defparam lat_mult_15.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_15.GSR = "DISABLED";
    defparam lat_mult_15.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_15.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_15.MULT_BYPASS = "DISABLED";
    defparam lat_mult_15.RESETMODE = "SYNC";
    ALU54B lat_alu_48 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n16396), .SIGNEDIB(n16469), .SIGNEDCIN(GND_net), 
           .A35(n16395), .A34(n16394), .A33(n16393), .A32(n16392), .A31(n16391), 
           .A30(n16390), .A29(n16389), .A28(n16388), .A27(n16387), .A26(n16386), 
           .A25(n16385), .A24(n16384), .A23(n16383), .A22(n16382), .A21(n16381), 
           .A20(n16380), .A19(n16379), .A18(n16378), .A17(n16377), .A16(n16376), 
           .A15(n16375), .A14(n16374), .A13(n16373), .A12(n16372), .A11(n16371), 
           .A10(n16370), .A9(n16369), .A8(n16368), .A7(n16367), .A6(n16366), 
           .A5(n16365), .A4(n16364), .A3(n16363), .A2(n16362), .A1(n16361), 
           .A0(n16360), .B35(n16468), .B34(n16467), .B33(n16466), .B32(n16465), 
           .B31(n16464), .B30(n16463), .B29(n16462), .B28(n16461), .B27(n16460), 
           .B26(n16459), .B25(n16458), .B24(n16457), .B23(n16456), .B22(n16455), 
           .B21(n16454), .B20(n16453), .B19(n16452), .B18(n16451), .B17(n16450), 
           .B16(n16449), .B15(n16448), .B14(n16447), .B13(n16446), .B12(n16445), 
           .B11(n16444), .B10(n16443), .B9(n16442), .B8(n16441), .B7(n16440), 
           .B6(n16439), .B5(n16438), .B4(n16437), .B3(n16436), .B2(n16435), 
           .B1(n16434), .B0(n16433), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n16432), .MA34(n16431), .MA33(n16430), .MA32(n16429), 
           .MA31(n16428), .MA30(n16427), .MA29(n16426), .MA28(n16425), 
           .MA27(n16424), .MA26(n16423), .MA25(n16422), .MA24(n16421), 
           .MA23(n16420), .MA22(n16419), .MA21(n16418), .MA20(n16417), 
           .MA19(n16416), .MA18(n16415), .MA17(n16414), .MA16(n16413), 
           .MA15(n16412), .MA14(n16411), .MA13(n16410), .MA12(n16409), 
           .MA11(n16408), .MA10(n16407), .MA9(n16406), .MA8(n16405), 
           .MA7(n16404), .MA6(n16403), .MA5(n16402), .MA4(n16401), .MA3(n16400), 
           .MA2(n16399), .MA1(n16398), .MA0(n16397), .MB35(n16505), 
           .MB34(n16504), .MB33(n16503), .MB32(n16502), .MB31(n16501), 
           .MB30(n16500), .MB29(n16499), .MB28(n16498), .MB27(n16497), 
           .MB26(n16496), .MB25(n16495), .MB24(n16494), .MB23(n16493), 
           .MB22(n16492), .MB21(n16491), .MB20(n16490), .MB19(n16489), 
           .MB18(n16488), .MB17(n16487), .MB16(n16486), .MB15(n16485), 
           .MB14(n16484), .MB13(n16483), .MB12(n16482), .MB11(n16481), 
           .MB10(n16480), .MB9(n16479), .MB8(n16478), .MB7(n16477), 
           .MB6(n16476), .MB5(n16475), .MB4(n16474), .MB3(n16473), .MB2(n16472), 
           .MB1(n16471), .MB0(n16470), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n16687), 
           .R52(n16686), .R51(n16685), .R50(n16684), .R49(n16683), .R48(n16682), 
           .R47(n16681), .R46(n16680), .R45(n16679), .R44(n16678), .R43(n16677), 
           .R42(n16676), .R41(n16675), .R40(n16674), .R39(n16673), .R38(n16672), 
           .R37(n16671), .R36(n16670), .R35(n16669), .R34(n16668), .R33(n16667), 
           .R32(n16666), .R31(n16665), .R30(n16664), .R29(n16663), .R28(n16662), 
           .R27(n16661), .R26(n16660), .R25(n16659), .R24(n16658), .R23(n16657), 
           .R22(n16656), .R21(n16655), .R20(n16654), .R19(n16653), .R18(n16652), 
           .R17(\op_r_23__N_1268[17] ), .R16(\op_r_23__N_1268[16] ), .R15(\op_r_23__N_1268[15] ), 
           .R14(\op_r_23__N_1268[14] ), .R13(\op_r_23__N_1268[13] ), .R12(\op_r_23__N_1268[12] ), 
           .R11(\op_r_23__N_1268[11] ), .R10(\op_r_23__N_1268[10] ), .R9(\op_r_23__N_1268[9] ), 
           .R8(\op_r_23__N_1268[8] ), .R7(\op_r_23__N_1268[7] ), .R6(\op_r_23__N_1268[6] ), 
           .R5(\op_r_23__N_1268[5] ), .R4(\op_r_23__N_1268[4] ), .R3(\op_r_23__N_1268[3] ), 
           .R2(\op_r_23__N_1268[2] ), .R1(\op_r_23__N_1268[1] ), .R0(\op_r_23__N_1268[0] ), 
           .SIGNEDR(n16688));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_48.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_48.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_48.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_48.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_48.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_48.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_48.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_48.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_48.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_48.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_48.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_48.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_48.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_48.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_48.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_48.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_48.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_48.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_48.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_48.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_48.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_48.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_48.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_48.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_48.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_48.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_48.REG_FLAG_CLK = "NONE";
    defparam lat_alu_48.REG_FLAG_CE = "CE0";
    defparam lat_alu_48.REG_FLAG_RST = "RST0";
    defparam lat_alu_48.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_48.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_48.MASK01 = "0x00000000000000";
    defparam lat_alu_48.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_48.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_48.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_48.CLK0_DIV = "ENABLED";
    defparam lat_alu_48.CLK1_DIV = "ENABLED";
    defparam lat_alu_48.CLK2_DIV = "ENABLED";
    defparam lat_alu_48.CLK3_DIV = "ENABLED";
    defparam lat_alu_48.MCPAT = "0x00000000000000";
    defparam lat_alu_48.MASKPAT = "0x00000000000000";
    defparam lat_alu_48.RNDPAT = "0x00000000000000";
    defparam lat_alu_48.GSR = "DISABLED";
    defparam lat_alu_48.RESETMODE = "SYNC";
    defparam lat_alu_48.MULT9_MODE = "DISABLED";
    defparam lat_alu_48.LEGACY = "DISABLED";
    MULT18X18D mult_975 (.A17(n34795), .A16(n34795), .A15(n34795), .A14(n34795), 
            .A13(n34795), .A12(n34795), .A11(n34795), .A10(n34795), 
            .A9(n34795), .A8(n34795), .A7(GND_net), .A6(GND_net), .A5(GND_net), 
            .A4(GND_net), .A3(GND_net), .A2(GND_net), .A1(GND_net), 
            .A0(GND_net), .B17(n11143), .B16(n11142), .B15(n11141), 
            .B14(n11140), .B13(n11139), .B12(n11138), .B11(n11137), 
            .B10(n11136), .B9(n11135), .B8(n11134), .B7(n11133), .B6(n11132), 
            .B5(n11131), .B4(n11130), .B3(n11129), .B2(n11128), .B1(n11127), 
            .B0(n11126), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14284), 
            .ROA16(n14283), .ROA15(n14282), .ROA14(n14281), .ROA13(n14280), 
            .ROA12(n14279), .ROA11(n14278), .ROA10(n14277), .ROA9(n14276), 
            .ROA8(n14275), .ROA7(n14274), .ROA6(n14273), .ROA5(n14272), 
            .ROA4(n14271), .ROA3(n14270), .ROA2(n14269), .ROA1(n14268), 
            .ROA0(n14267), .ROB17(n14302), .ROB16(n14301), .ROB15(n14300), 
            .ROB14(n14299), .ROB13(n14298), .ROB12(n14297), .ROB11(n14296), 
            .ROB10(n14295), .ROB9(n14294), .ROB8(n14293), .ROB7(n14292), 
            .ROB6(n14291), .ROB5(n14290), .ROB4(n14289), .ROB3(n14288), 
            .ROB2(n14287), .ROB1(n14286), .ROB0(n14285), .P35(n14339), 
            .P34(n14338), .P33(n14337), .P32(n14336), .P31(n14335), 
            .P30(n14334), .P29(n14333), .P28(n14332), .P27(n14331), 
            .P26(n14330), .P25(n14329), .P24(n14328), .P23(n14327), 
            .P22(n14326), .P21(n14325), .P20(n14324), .P19(n14323), 
            .P18(n14322), .P17(n14321), .P16(n14320), .P15(n14319), 
            .P14(n14318), .P13(n14317), .P12(n14316), .P11(n14315), 
            .P10(n14314), .P9(n14313), .P8(n14312), .P7(n14311), .P6(n14310), 
            .P5(n14309), .P4(n14308), .P3(n14307), .P2(n14306), .P1(n14305), 
            .P0(n14304), .SIGNEDP(n14303));
    defparam mult_975.REG_INPUTA_CLK = "NONE";
    defparam mult_975.REG_INPUTA_CE = "CE0";
    defparam mult_975.REG_INPUTA_RST = "RST0";
    defparam mult_975.REG_INPUTB_CLK = "NONE";
    defparam mult_975.REG_INPUTB_CE = "CE0";
    defparam mult_975.REG_INPUTB_RST = "RST0";
    defparam mult_975.REG_INPUTC_CLK = "NONE";
    defparam mult_975.REG_INPUTC_CE = "CE0";
    defparam mult_975.REG_INPUTC_RST = "RST0";
    defparam mult_975.REG_PIPELINE_CLK = "NONE";
    defparam mult_975.REG_PIPELINE_CE = "CE0";
    defparam mult_975.REG_PIPELINE_RST = "RST0";
    defparam mult_975.REG_OUTPUT_CLK = "NONE";
    defparam mult_975.REG_OUTPUT_CE = "CE0";
    defparam mult_975.REG_OUTPUT_RST = "RST0";
    defparam mult_975.CLK0_DIV = "ENABLED";
    defparam mult_975.CLK1_DIV = "ENABLED";
    defparam mult_975.CLK2_DIV = "ENABLED";
    defparam mult_975.CLK3_DIV = "ENABLED";
    defparam mult_975.HIGHSPEED_CLK = "NONE";
    defparam mult_975.GSR = "DISABLED";
    defparam mult_975.CAS_MATCH_REG = "FALSE";
    defparam mult_975.SOURCEB_MODE = "B_SHIFT";
    defparam mult_975.MULT_BYPASS = "DISABLED";
    defparam mult_975.RESETMODE = "SYNC";
    MULT18X18D lat_mult_46 (.A17(shift_2_dout_i[17]), .A16(shift_2_dout_i[16]), 
            .A15(shift_2_dout_i[15]), .A14(shift_2_dout_i[14]), .A13(shift_2_dout_i[13]), 
            .A12(shift_2_dout_i[12]), .A11(shift_2_dout_i[11]), .A10(shift_2_dout_i[10]), 
            .A9(shift_2_dout_i[9]), .A8(shift_2_dout_i[8]), .A7(shift_2_dout_i[7]), 
            .A6(shift_2_dout_i[6]), .A5(shift_2_dout_i[5]), .A4(shift_2_dout_i[4]), 
            .A3(shift_2_dout_i[3]), .A2(shift_2_dout_i[2]), .A1(shift_2_dout_i[1]), 
            .A0(shift_2_dout_i[0]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(GND_net), .B7(GND_net), 
            .B6(GND_net), .B5(GND_net), .B4(GND_net), .B3(GND_net), 
            .B2(GND_net), .B1(GND_net), .B0(GND_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n16523), .ROA16(n16522), .ROA15(n16521), 
            .ROA14(n16520), .ROA13(n16519), .ROA12(n16518), .ROA11(n16517), 
            .ROA10(n16516), .ROA9(n16515), .ROA8(n16514), .ROA7(n16513), 
            .ROA6(n16512), .ROA5(n16511), .ROA4(n16510), .ROA3(n16509), 
            .ROA2(n16508), .ROA1(n16507), .ROA0(n16506), .ROB17(n16541), 
            .ROB16(n16540), .ROB15(n16539), .ROB14(n16538), .ROB13(n16537), 
            .ROB12(n16536), .ROB11(n16535), .ROB10(n16534), .ROB9(n16533), 
            .ROB8(n16532), .ROB7(n16531), .ROB6(n16530), .ROB5(n16529), 
            .ROB4(n16528), .ROB3(n16527), .ROB2(n16526), .ROB1(n16525), 
            .ROB0(n16524), .P35(n16578), .P34(n16577), .P33(n16576), 
            .P32(n16575), .P31(n16574), .P30(n16573), .P29(n16572), 
            .P28(n16571), .P27(n16570), .P26(n16569), .P25(n16568), 
            .P24(n16567), .P23(n16566), .P22(n16565), .P21(n16564), 
            .P20(n16563), .P19(n16562), .P18(n16561), .P17(n16560), 
            .P16(n16559), .P15(n16558), .P14(n16557), .P13(n16556), 
            .P12(n16555), .P11(n16554), .P10(n16553), .P9(n16552), .P8(n16551), 
            .P7(n16550), .P6(n16549), .P5(n16548), .P4(n16547), .P3(n16546), 
            .P2(n16545), .P1(n16544), .P0(n16543), .SIGNEDP(n16542));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_46.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_46.REG_INPUTA_CE = "CE0";
    defparam lat_mult_46.REG_INPUTA_RST = "RST0";
    defparam lat_mult_46.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_46.REG_INPUTB_CE = "CE0";
    defparam lat_mult_46.REG_INPUTB_RST = "RST0";
    defparam lat_mult_46.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_46.REG_INPUTC_CE = "CE0";
    defparam lat_mult_46.REG_INPUTC_RST = "RST0";
    defparam lat_mult_46.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_46.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_46.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_46.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_46.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_46.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_46.CLK0_DIV = "ENABLED";
    defparam lat_mult_46.CLK1_DIV = "ENABLED";
    defparam lat_mult_46.CLK2_DIV = "ENABLED";
    defparam lat_mult_46.CLK3_DIV = "ENABLED";
    defparam lat_mult_46.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_46.GSR = "DISABLED";
    defparam lat_mult_46.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_46.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_46.MULT_BYPASS = "DISABLED";
    defparam lat_mult_46.RESETMODE = "SYNC";
    MULT18X18D lat_mult_45 (.A17(shift_2_dout_i[23]), .A16(shift_2_dout_i[23]), 
            .A15(shift_2_dout_i[23]), .A14(shift_2_dout_i[23]), .A13(shift_2_dout_i[23]), 
            .A12(shift_2_dout_i[23]), .A11(shift_2_dout_i[23]), .A10(shift_2_dout_i[23]), 
            .A9(shift_2_dout_i[23]), .A8(shift_2_dout_i[23]), .A7(shift_2_dout_i[23]), 
            .A6(shift_2_dout_i[23]), .A5(shift_2_dout_i[23]), .A4(shift_2_dout_i[22]), 
            .A3(shift_2_dout_i[21]), .A2(shift_2_dout_i[20]), .A1(shift_2_dout_i[19]), 
            .A0(shift_2_dout_i[18]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(VCC_net), .B7(GND_net), 
            .B6(GND_net), .B5(GND_net), .B4(GND_net), .B3(GND_net), 
            .B2(GND_net), .B1(GND_net), .B0(GND_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n16450), .ROA16(n16449), .ROA15(n16448), 
            .ROA14(n16447), .ROA13(n16446), .ROA12(n16445), .ROA11(n16444), 
            .ROA10(n16443), .ROA9(n16442), .ROA8(n16441), .ROA7(n16440), 
            .ROA6(n16439), .ROA5(n16438), .ROA4(n16437), .ROA3(n16436), 
            .ROA2(n16435), .ROA1(n16434), .ROA0(n16433), .ROB17(n16468), 
            .ROB16(n16467), .ROB15(n16466), .ROB14(n16465), .ROB13(n16464), 
            .ROB12(n16463), .ROB11(n16462), .ROB10(n16461), .ROB9(n16460), 
            .ROB8(n16459), .ROB7(n16458), .ROB6(n16457), .ROB5(n16456), 
            .ROB4(n16455), .ROB3(n16454), .ROB2(n16453), .ROB1(n16452), 
            .ROB0(n16451), .P35(n16505), .P34(n16504), .P33(n16503), 
            .P32(n16502), .P31(n16501), .P30(n16500), .P29(n16499), 
            .P28(n16498), .P27(n16497), .P26(n16496), .P25(n16495), 
            .P24(n16494), .P23(n16493), .P22(n16492), .P21(n16491), 
            .P20(n16490), .P19(n16489), .P18(n16488), .P17(n16487), 
            .P16(n16486), .P15(n16485), .P14(n16484), .P13(n16483), 
            .P12(n16482), .P11(n16481), .P10(n16480), .P9(n16479), .P8(n16478), 
            .P7(n16477), .P6(n16476), .P5(n16475), .P4(n16474), .P3(n16473), 
            .P2(n16472), .P1(n16471), .P0(n16470), .SIGNEDP(n16469));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_45.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_45.REG_INPUTA_CE = "CE0";
    defparam lat_mult_45.REG_INPUTA_RST = "RST0";
    defparam lat_mult_45.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_45.REG_INPUTB_CE = "CE0";
    defparam lat_mult_45.REG_INPUTB_RST = "RST0";
    defparam lat_mult_45.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_45.REG_INPUTC_CE = "CE0";
    defparam lat_mult_45.REG_INPUTC_RST = "RST0";
    defparam lat_mult_45.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_45.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_45.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_45.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_45.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_45.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_45.CLK0_DIV = "ENABLED";
    defparam lat_mult_45.CLK1_DIV = "ENABLED";
    defparam lat_mult_45.CLK2_DIV = "ENABLED";
    defparam lat_mult_45.CLK3_DIV = "ENABLED";
    defparam lat_mult_45.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_45.GSR = "DISABLED";
    defparam lat_mult_45.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_45.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_45.MULT_BYPASS = "DISABLED";
    defparam lat_mult_45.RESETMODE = "SYNC";
    MULT18X18D mult_8 (.A17(shift_2_dout_i[17]), .A16(shift_2_dout_i[16]), 
            .A15(shift_2_dout_i[15]), .A14(shift_2_dout_i[14]), .A13(shift_2_dout_i[13]), 
            .A12(shift_2_dout_i[12]), .A11(shift_2_dout_i[11]), .A10(shift_2_dout_i[10]), 
            .A9(shift_2_dout_i[9]), .A8(shift_2_dout_i[8]), .A7(shift_2_dout_i[7]), 
            .A6(shift_2_dout_i[6]), .A5(shift_2_dout_i[5]), .A4(shift_2_dout_i[4]), 
            .A3(shift_2_dout_i[3]), .A2(shift_2_dout_i[2]), .A1(shift_2_dout_i[1]), 
            .A0(shift_2_dout_i[0]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(VCC_net), .B7(GND_net), 
            .B6(GND_net), .B5(GND_net), .B4(GND_net), .B3(GND_net), 
            .B2(GND_net), .B1(GND_net), .B0(GND_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n16377), .ROA16(n16376), .ROA15(n16375), 
            .ROA14(n16374), .ROA13(n16373), .ROA12(n16372), .ROA11(n16371), 
            .ROA10(n16370), .ROA9(n16369), .ROA8(n16368), .ROA7(n16367), 
            .ROA6(n16366), .ROA5(n16365), .ROA4(n16364), .ROA3(n16363), 
            .ROA2(n16362), .ROA1(n16361), .ROA0(n16360), .ROB17(n16395), 
            .ROB16(n16394), .ROB15(n16393), .ROB14(n16392), .ROB13(n16391), 
            .ROB12(n16390), .ROB11(n16389), .ROB10(n16388), .ROB9(n16387), 
            .ROB8(n16386), .ROB7(n16385), .ROB6(n16384), .ROB5(n16383), 
            .ROB4(n16382), .ROB3(n16381), .ROB2(n16380), .ROB1(n16379), 
            .ROB0(n16378), .P35(n16432), .P34(n16431), .P33(n16430), 
            .P32(n16429), .P31(n16428), .P30(n16427), .P29(n16426), 
            .P28(n16425), .P27(n16424), .P26(n16423), .P25(n16422), 
            .P24(n16421), .P23(n16420), .P22(n16419), .P21(n16418), 
            .P20(n16417), .P19(n16416), .P18(n16415), .P17(n16414), 
            .P16(n16413), .P15(n16412), .P14(n16411), .P13(n16410), 
            .P12(n16409), .P11(n16408), .P10(n16407), .P9(n16406), .P8(n16405), 
            .P7(n16404), .P6(n16403), .P5(n16402), .P4(n16401), .P3(n16400), 
            .P2(n16399), .P1(n16398), .P0(n16397), .SIGNEDP(n16396));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam mult_8.REG_INPUTA_CLK = "NONE";
    defparam mult_8.REG_INPUTA_CE = "CE0";
    defparam mult_8.REG_INPUTA_RST = "RST0";
    defparam mult_8.REG_INPUTB_CLK = "NONE";
    defparam mult_8.REG_INPUTB_CE = "CE0";
    defparam mult_8.REG_INPUTB_RST = "RST0";
    defparam mult_8.REG_INPUTC_CLK = "NONE";
    defparam mult_8.REG_INPUTC_CE = "CE0";
    defparam mult_8.REG_INPUTC_RST = "RST0";
    defparam mult_8.REG_PIPELINE_CLK = "NONE";
    defparam mult_8.REG_PIPELINE_CE = "CE0";
    defparam mult_8.REG_PIPELINE_RST = "RST0";
    defparam mult_8.REG_OUTPUT_CLK = "NONE";
    defparam mult_8.REG_OUTPUT_CE = "CE0";
    defparam mult_8.REG_OUTPUT_RST = "RST0";
    defparam mult_8.CLK0_DIV = "ENABLED";
    defparam mult_8.CLK1_DIV = "ENABLED";
    defparam mult_8.CLK2_DIV = "ENABLED";
    defparam mult_8.CLK3_DIV = "ENABLED";
    defparam mult_8.HIGHSPEED_CLK = "NONE";
    defparam mult_8.GSR = "DISABLED";
    defparam mult_8.CAS_MATCH_REG = "FALSE";
    defparam mult_8.SOURCEB_MODE = "B_SHIFT";
    defparam mult_8.MULT_BYPASS = "DISABLED";
    defparam mult_8.RESETMODE = "SYNC";
    ND2 ND2_t28 (.A(n34795), .B(n120), .Z(mult_24s_7s_0_mult_2_11_n2)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t31 (.A(n34795), .B(n126), .Z(mult_24s_7s_0_mult_0_11_n3)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t32 (.A(GND_net), .B(n126), .Z(\op_i_23__N_1310[0] )) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(297[10:65])
    ND2 ND2_t30 (.A(n34795), .B(n123), .Z(mult_24s_7s_0_mult_0_11_n1)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t29 (.A(GND_net), .B(n120), .Z(mult_24s_7s_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(303[10:65])
    ND2 ND2_t27 (.A(n34795), .B(n117), .Z(mult_24s_7s_0_mult_2_11_n1)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t26 (.A(GND_net), .B(n114), .Z(mult_24s_7s_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(309[10:65])
    ND2 ND2_t24 (.A(n34795), .B(n111), .Z(mult_24s_7s_0_mult_4_11_n1)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t23 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t22 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_7)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t21 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t20 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_9)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t19 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t18 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_11)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t17 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t16 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_13)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t15 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t14 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_15)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t13 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t12 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_17)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t11 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t10 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_19)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t9 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t8 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_21)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t7 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t6 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_23)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t5 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t4 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_25)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t3 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t2 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_27)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t1 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t0 (.A(n34795), .B(GND_net), .Z(mult_24s_7s_0_pp_3_29)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(361[10:66])
    CCU2C mult_24s_7s_0_Cadd_0_12 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco), .S0(mult_24s_7s_0_pp_0_25)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(375[11] 377[80])
    defparam mult_24s_7s_0_Cadd_0_12.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_0_12.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_0_12.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_Cadd_0_12.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_cin_lr_add_2 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(mult_24s_7s_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(383[11] 385[77])
    defparam mult_24s_7s_0_cin_lr_add_2.INIT0 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_2.INIT1 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_cin_lr_add_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_Cadd_2_12 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_1), .S0(mult_24s_7s_0_pp_1_27)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(391[11] 394[17])
    defparam mult_24s_7s_0_Cadd_2_12.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_2_12.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_2_12.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_Cadd_2_12.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_cin_lr_add_4 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(mult_24s_7s_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(400[11] 402[77])
    defparam mult_24s_7s_0_cin_lr_add_4.INIT0 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_4.INIT1 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_cin_lr_add_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_Cadd_4_12 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_2), .S0(mult_24s_7s_0_pp_2_29)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(408[11] 411[17])
    defparam mult_24s_7s_0_Cadd_4_12.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_4_12.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_4_12.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_Cadd_4_12.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_0_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_2), .B1(mult_24s_7s_0_pp_1_2), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_mult_24s_7s_0_0_1), .S1(\op_i_23__N_1310[2] )) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(417[11] 420[37])
    defparam Cadd_mult_24s_7s_0_0_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_1.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_0_1.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_2 (.A0(mult_24s_7s_0_pp_0_3), .B0(mult_24s_7s_0_pp_1_3), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_4), .B1(mult_24s_7s_0_pp_1_4), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_1), .COUT(co_mult_24s_7s_0_0_2), 
          .S0(\op_i_23__N_1310[3] ), .S1(s_mult_24s_7s_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(426[11] 429[89])
    defparam mult_24s_7s_0_add_0_2.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_2.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_3 (.A0(mult_24s_7s_0_pp_0_5), .B0(mult_24s_7s_0_pp_1_5), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_6), .B1(mult_24s_7s_0_pp_1_6), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_2), .COUT(co_mult_24s_7s_0_0_3), 
          .S0(s_mult_24s_7s_0_0_5), .S1(s_mult_24s_7s_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(435[11] 438[89])
    defparam mult_24s_7s_0_add_0_3.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_3.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_3.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_3.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_4 (.A0(mult_24s_7s_0_pp_0_7), .B0(mult_24s_7s_0_pp_1_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_8), .B1(mult_24s_7s_0_pp_1_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_3), .COUT(co_mult_24s_7s_0_0_4), 
          .S0(s_mult_24s_7s_0_0_7), .S1(s_mult_24s_7s_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(444[11] 447[89])
    defparam mult_24s_7s_0_add_0_4.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_4.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_5 (.A0(mult_24s_7s_0_pp_0_9), .B0(mult_24s_7s_0_pp_1_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_10), .B1(mult_24s_7s_0_pp_1_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_4), .COUT(co_mult_24s_7s_0_0_5), 
          .S0(s_mult_24s_7s_0_0_9), .S1(s_mult_24s_7s_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(453[11] 456[90])
    defparam mult_24s_7s_0_add_0_5.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_5.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_5.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_5.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_6 (.A0(mult_24s_7s_0_pp_0_11), .B0(mult_24s_7s_0_pp_1_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_12), .B1(mult_24s_7s_0_pp_1_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_5), .COUT(co_mult_24s_7s_0_0_6), 
          .S0(s_mult_24s_7s_0_0_11), .S1(s_mult_24s_7s_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(462[11] 465[91])
    defparam mult_24s_7s_0_add_0_6.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_6.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_6.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_6.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_7 (.A0(mult_24s_7s_0_pp_0_13), .B0(mult_24s_7s_0_pp_1_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_14), .B1(mult_24s_7s_0_pp_1_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_6), .COUT(co_mult_24s_7s_0_0_7), 
          .S0(s_mult_24s_7s_0_0_13), .S1(s_mult_24s_7s_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(471[11] 474[91])
    defparam mult_24s_7s_0_add_0_7.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_7.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_7.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_7.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_8 (.A0(mult_24s_7s_0_pp_0_15), .B0(mult_24s_7s_0_pp_1_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_16), .B1(mult_24s_7s_0_pp_1_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_7), .COUT(co_mult_24s_7s_0_0_8), 
          .S0(s_mult_24s_7s_0_0_15), .S1(s_mult_24s_7s_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(480[11] 483[91])
    defparam mult_24s_7s_0_add_0_8.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_8.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_8.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_8.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_9 (.A0(mult_24s_7s_0_pp_0_17), .B0(mult_24s_7s_0_pp_1_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_18), .B1(mult_24s_7s_0_pp_1_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_8), .COUT(co_mult_24s_7s_0_0_9), 
          .S0(s_mult_24s_7s_0_0_17), .S1(s_mult_24s_7s_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(489[11] 492[91])
    defparam mult_24s_7s_0_add_0_9.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_9.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_9.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_9.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_10 (.A0(mult_24s_7s_0_pp_0_19), .B0(mult_24s_7s_0_pp_1_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_20), .B1(mult_24s_7s_0_pp_1_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_9), .COUT(co_mult_24s_7s_0_0_10), 
          .S0(s_mult_24s_7s_0_0_19), .S1(s_mult_24s_7s_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(498[11] 501[92])
    defparam mult_24s_7s_0_add_0_10.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_10.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_10.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_10.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_11 (.A0(mult_24s_7s_0_pp_0_21), .B0(mult_24s_7s_0_pp_1_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_22), .B1(mult_24s_7s_0_pp_1_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_10), .COUT(co_mult_24s_7s_0_0_11), 
          .S0(s_mult_24s_7s_0_0_21), .S1(s_mult_24s_7s_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(507[11] 510[92])
    defparam mult_24s_7s_0_add_0_11.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_11.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_11.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_11.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_12 (.A0(mult_24s_7s_0_pp_0_23), .B0(mult_24s_7s_0_pp_1_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_24), .B1(mult_24s_7s_0_pp_1_24), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_11), .COUT(co_mult_24s_7s_0_0_12), 
          .S0(s_mult_24s_7s_0_0_23), .S1(s_mult_24s_7s_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(516[11] 519[92])
    defparam mult_24s_7s_0_add_0_12.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_12.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_12.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_12.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_13 (.A0(mult_24s_7s_0_pp_0_25), .B0(mult_24s_7s_0_pp_1_25), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(mult_24s_7s_0_pp_1_26), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_12), .COUT(co_mult_24s_7s_0_0_13), 
          .S0(s_mult_24s_7s_0_0_25), .S1(s_mult_24s_7s_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(525[11] 528[92])
    defparam mult_24s_7s_0_add_0_13.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_13.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_13.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_13.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_14 (.A0(GND_net), .B0(mult_24s_7s_0_pp_1_27), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_13), .COUT(co_mult_24s_7s_0_0_14), 
          .S0(s_mult_24s_7s_0_0_27), .S1(s_mult_24s_7s_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(534[11] 537[65])
    defparam mult_24s_7s_0_add_0_14.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_14.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_14.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_14.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_0_15 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_mult_24s_7s_0_0_14), .S0(s_mult_24s_7s_0_0_29)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(543[11] 546[24])
    defparam Cadd_mult_24s_7s_0_0_15.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_15.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_15.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_0_15.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_1_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_6), .B1(mult_24s_7s_0_pp_3_6), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_mult_24s_7s_0_1_1), .S1(s_mult_24s_7s_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(552[11] 555[37])
    defparam Cadd_mult_24s_7s_0_1_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_1_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_1_1.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_1_1.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_2 (.A0(mult_24s_7s_0_pp_2_7), .B0(mult_24s_7s_0_pp_3_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_8), .B1(mult_24s_7s_0_pp_3_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_1), .COUT(co_mult_24s_7s_0_1_2), 
          .S0(s_mult_24s_7s_0_1_7), .S1(s_mult_24s_7s_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(561[11] 564[89])
    defparam mult_24s_7s_0_add_1_2.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_2.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_3 (.A0(mult_24s_7s_0_pp_2_9), .B0(mult_24s_7s_0_pp_3_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_10), .B1(mult_24s_7s_0_pp_3_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_2), .COUT(co_mult_24s_7s_0_1_3), 
          .S0(s_mult_24s_7s_0_1_9), .S1(s_mult_24s_7s_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(570[11] 573[90])
    defparam mult_24s_7s_0_add_1_3.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_3.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_3.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_3.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_4 (.A0(mult_24s_7s_0_pp_2_11), .B0(mult_24s_7s_0_pp_3_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_12), .B1(mult_24s_7s_0_pp_3_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_3), .COUT(co_mult_24s_7s_0_1_4), 
          .S0(s_mult_24s_7s_0_1_11), .S1(s_mult_24s_7s_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(579[11] 582[91])
    defparam mult_24s_7s_0_add_1_4.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_4.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_5 (.A0(mult_24s_7s_0_pp_2_13), .B0(mult_24s_7s_0_pp_3_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_14), .B1(mult_24s_7s_0_pp_3_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_4), .COUT(co_mult_24s_7s_0_1_5), 
          .S0(s_mult_24s_7s_0_1_13), .S1(s_mult_24s_7s_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(588[11] 591[91])
    defparam mult_24s_7s_0_add_1_5.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_5.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_5.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_5.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_6 (.A0(mult_24s_7s_0_pp_2_15), .B0(mult_24s_7s_0_pp_3_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_16), .B1(mult_24s_7s_0_pp_3_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_5), .COUT(co_mult_24s_7s_0_1_6), 
          .S0(s_mult_24s_7s_0_1_15), .S1(s_mult_24s_7s_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(597[11] 600[91])
    defparam mult_24s_7s_0_add_1_6.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_6.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_6.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_6.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_7 (.A0(mult_24s_7s_0_pp_2_17), .B0(mult_24s_7s_0_pp_3_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_18), .B1(mult_24s_7s_0_pp_3_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_6), .COUT(co_mult_24s_7s_0_1_7), 
          .S0(s_mult_24s_7s_0_1_17), .S1(s_mult_24s_7s_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(606[11] 609[91])
    defparam mult_24s_7s_0_add_1_7.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_7.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_7.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_7.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_8 (.A0(mult_24s_7s_0_pp_2_19), .B0(mult_24s_7s_0_pp_3_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_20), .B1(mult_24s_7s_0_pp_3_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_7), .COUT(co_mult_24s_7s_0_1_8), 
          .S0(s_mult_24s_7s_0_1_19), .S1(s_mult_24s_7s_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(615[11] 618[91])
    defparam mult_24s_7s_0_add_1_8.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_8.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_8.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_8.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_9 (.A0(mult_24s_7s_0_pp_2_21), .B0(mult_24s_7s_0_pp_3_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_22), .B1(mult_24s_7s_0_pp_3_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_8), .COUT(co_mult_24s_7s_0_1_9), 
          .S0(s_mult_24s_7s_0_1_21), .S1(s_mult_24s_7s_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(624[11] 627[91])
    defparam mult_24s_7s_0_add_1_9.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_9.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_9.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_9.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_10 (.A0(mult_24s_7s_0_pp_2_23), .B0(mult_24s_7s_0_pp_3_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_24), .B1(mult_24s_7s_0_pp_3_24), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_9), .COUT(co_mult_24s_7s_0_1_10), 
          .S0(s_mult_24s_7s_0_1_23), .S1(s_mult_24s_7s_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(633[11] 636[92])
    defparam mult_24s_7s_0_add_1_10.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_10.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_10.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_10.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_11 (.A0(mult_24s_7s_0_pp_2_25), .B0(mult_24s_7s_0_pp_3_25), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_26), .B1(mult_24s_7s_0_pp_3_26), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_10), .COUT(co_mult_24s_7s_0_1_11), 
          .S0(s_mult_24s_7s_0_1_25), .S1(s_mult_24s_7s_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(642[11] 645[92])
    defparam mult_24s_7s_0_add_1_11.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_11.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_11.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_11.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_12 (.A0(mult_24s_7s_0_pp_2_27), .B0(mult_24s_7s_0_pp_3_27), 
          .C0(VCC_net), .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_28), .B1(mult_24s_7s_0_pp_3_28), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_11), .COUT(co_mult_24s_7s_0_1_12), 
          .S0(s_mult_24s_7s_0_1_27), .S1(s_mult_24s_7s_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(651[11] 654[92])
    defparam mult_24s_7s_0_add_1_12.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_12.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_12.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_12.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_13 (.A0(mult_24s_7s_0_pp_2_29), .B0(mult_24s_7s_0_pp_3_29), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_12), .S0(s_mult_24s_7s_0_1_29), 
          .S1(s_mult_24s_7s_0_1_30)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(660[11] 663[65])
    defparam mult_24s_7s_0_add_1_13.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_13.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_13.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_13.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_2_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(s_mult_24s_7s_0_0_4), .B1(mult_24s_7s_0_pp_2_4), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_mult_24s_7s_0_2_1), .S1(\op_i_23__N_1310[4] )) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(669[11] 672[37])
    defparam Cadd_mult_24s_7s_0_2_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_2_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_2_1.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_2_1.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_2 (.A0(s_mult_24s_7s_0_0_5), .B0(mult_24s_7s_0_pp_2_5), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_6), .B1(s_mult_24s_7s_0_1_6), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_1), .COUT(co_mult_24s_7s_0_2_2), 
          .S0(\op_i_23__N_1310[5] ), .S1(s_mult_24s_7s_0_2_6)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(678[11] 681[89])
    defparam mult_24s_7s_0_add_2_2.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_2.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_3 (.A0(s_mult_24s_7s_0_0_7), .B0(s_mult_24s_7s_0_1_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_8), .B1(s_mult_24s_7s_0_1_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_2), .COUT(co_mult_24s_7s_0_2_3), 
          .S0(s_mult_24s_7s_0_2_7), .S1(s_mult_24s_7s_0_2_8)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(687[11] 690[89])
    defparam mult_24s_7s_0_add_2_3.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_3.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_3.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_3.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_4 (.A0(s_mult_24s_7s_0_0_9), .B0(s_mult_24s_7s_0_1_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_10), .B1(s_mult_24s_7s_0_1_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_3), .COUT(co_mult_24s_7s_0_2_4), 
          .S0(s_mult_24s_7s_0_2_9), .S1(s_mult_24s_7s_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(696[11] 699[90])
    defparam mult_24s_7s_0_add_2_4.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_4.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_5 (.A0(s_mult_24s_7s_0_0_11), .B0(s_mult_24s_7s_0_1_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_12), .B1(s_mult_24s_7s_0_1_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_4), .COUT(co_mult_24s_7s_0_2_5), 
          .S0(s_mult_24s_7s_0_2_11), .S1(s_mult_24s_7s_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(705[11] 708[91])
    defparam mult_24s_7s_0_add_2_5.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_5.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_5.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_5.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_6 (.A0(s_mult_24s_7s_0_0_13), .B0(s_mult_24s_7s_0_1_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_14), .B1(s_mult_24s_7s_0_1_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_5), .COUT(co_mult_24s_7s_0_2_6), 
          .S0(s_mult_24s_7s_0_2_13), .S1(s_mult_24s_7s_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(714[11] 717[91])
    defparam mult_24s_7s_0_add_2_6.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_6.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_6.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_6.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_7 (.A0(s_mult_24s_7s_0_0_15), .B0(s_mult_24s_7s_0_1_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_16), .B1(s_mult_24s_7s_0_1_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_6), .COUT(co_mult_24s_7s_0_2_7), 
          .S0(s_mult_24s_7s_0_2_15), .S1(s_mult_24s_7s_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(723[11] 726[91])
    defparam mult_24s_7s_0_add_2_7.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_7.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_7.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_7.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_8 (.A0(s_mult_24s_7s_0_0_17), .B0(s_mult_24s_7s_0_1_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_18), .B1(s_mult_24s_7s_0_1_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_7), .COUT(co_mult_24s_7s_0_2_8), 
          .S0(s_mult_24s_7s_0_2_17), .S1(s_mult_24s_7s_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(732[11] 735[91])
    defparam mult_24s_7s_0_add_2_8.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_8.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_8.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_8.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_9 (.A0(s_mult_24s_7s_0_0_19), .B0(s_mult_24s_7s_0_1_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_20), .B1(s_mult_24s_7s_0_1_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_8), .COUT(co_mult_24s_7s_0_2_9), 
          .S0(s_mult_24s_7s_0_2_19), .S1(s_mult_24s_7s_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(741[11] 744[91])
    defparam mult_24s_7s_0_add_2_9.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_9.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_9.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_9.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_10 (.A0(s_mult_24s_7s_0_0_21), .B0(s_mult_24s_7s_0_1_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_22), .B1(s_mult_24s_7s_0_1_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_9), .COUT(co_mult_24s_7s_0_2_10), 
          .S0(s_mult_24s_7s_0_2_21), .S1(s_mult_24s_7s_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(750[11] 753[92])
    defparam mult_24s_7s_0_add_2_10.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_10.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_10.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_10.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_11 (.A0(s_mult_24s_7s_0_0_23), .B0(s_mult_24s_7s_0_1_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_24), .B1(s_mult_24s_7s_0_1_24), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_10), .COUT(co_mult_24s_7s_0_2_11), 
          .S0(s_mult_24s_7s_0_2_23), .S1(s_mult_24s_7s_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(759[11] 762[92])
    defparam mult_24s_7s_0_add_2_11.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_11.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_11.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_11.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_12 (.A0(s_mult_24s_7s_0_0_25), .B0(s_mult_24s_7s_0_1_25), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_26), .B1(s_mult_24s_7s_0_1_26), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_11), .COUT(co_mult_24s_7s_0_2_12), 
          .S0(s_mult_24s_7s_0_2_25), .S1(s_mult_24s_7s_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(768[11] 771[92])
    defparam mult_24s_7s_0_add_2_12.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_12.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_12.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_12.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_13 (.A0(s_mult_24s_7s_0_0_27), .B0(s_mult_24s_7s_0_1_27), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_0_28), .B1(s_mult_24s_7s_0_1_28), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_12), .COUT(co_mult_24s_7s_0_2_13), 
          .S0(s_mult_24s_7s_0_2_27), .S1(s_mult_24s_7s_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(777[11] 780[92])
    defparam mult_24s_7s_0_add_2_13.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_13.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_13.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_13.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_14 (.A0(s_mult_24s_7s_0_0_29), .B0(s_mult_24s_7s_0_1_29), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(s_mult_24s_7s_0_1_30), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_13), .S0(s_mult_24s_7s_0_2_29), 
          .S1(s_mult_24s_7s_0_2_30)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(786[11] 789[92])
    defparam mult_24s_7s_0_add_2_14.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_14.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_14.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_14.INJECT1_1 = "NO";
    CCU2C Cadd_t_mult_24s_7s_0_3_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(s_mult_24s_7s_0_2_6), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co_t_mult_24s_7s_0_3_1), .S1(n89)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(795[11] 797[97])
    defparam Cadd_t_mult_24s_7s_0_3_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_t_mult_24s_7s_0_3_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_t_mult_24s_7s_0_3_1.INJECT1_0 = "NO";
    defparam Cadd_t_mult_24s_7s_0_3_1.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_2 (.A0(s_mult_24s_7s_0_2_7), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_8), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_1), .COUT(co_t_mult_24s_7s_0_3_2), 
          .S0(n88), .S1(n87)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(803[11] 806[50])
    defparam t_mult_24s_7s_0_add_3_2.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_2.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_2.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_2.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_3 (.A0(s_mult_24s_7s_0_2_9), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_10), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_2), .COUT(co_t_mult_24s_7s_0_3_3), 
          .S0(n86), .S1(n85)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(812[11] 815[51])
    defparam t_mult_24s_7s_0_add_3_3.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_3.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_3.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_3.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_4 (.A0(s_mult_24s_7s_0_2_11), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_12), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_3), .COUT(co_t_mult_24s_7s_0_3_4), 
          .S0(n84), .S1(n83)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(821[11] 824[51])
    defparam t_mult_24s_7s_0_add_3_4.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_4.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_4.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_4.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_5 (.A0(s_mult_24s_7s_0_2_13), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_14), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_4), .COUT(co_t_mult_24s_7s_0_3_5), 
          .S0(n82), .S1(n81)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(830[11] 833[51])
    defparam t_mult_24s_7s_0_add_3_5.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_5.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_5.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_5.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_6 (.A0(s_mult_24s_7s_0_2_15), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_16), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_5), .COUT(co_t_mult_24s_7s_0_3_6), 
          .S0(n80), .S1(n79)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(839[11] 842[51])
    defparam t_mult_24s_7s_0_add_3_6.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_6.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_6.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_6.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_7 (.A0(s_mult_24s_7s_0_2_17), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_18), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_6), .COUT(co_t_mult_24s_7s_0_3_7), 
          .S0(n78), .S1(n77)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(848[11] 851[51])
    defparam t_mult_24s_7s_0_add_3_7.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_7.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_7.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_7.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_8 (.A0(s_mult_24s_7s_0_2_19), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_20), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_7), .COUT(co_t_mult_24s_7s_0_3_8), 
          .S0(n76), .S1(n75)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(857[11] 860[51])
    defparam t_mult_24s_7s_0_add_3_8.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_8.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_8.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_8.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_9 (.A0(s_mult_24s_7s_0_2_21), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_22), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_8), .COUT(co_t_mult_24s_7s_0_3_9), 
          .S0(n74), .S1(n73)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(866[11] 869[51])
    defparam t_mult_24s_7s_0_add_3_9.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_9.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_9.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_9.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_10 (.A0(s_mult_24s_7s_0_2_23), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_24), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_9), .COUT(co_t_mult_24s_7s_0_3_10), 
          .S0(n72), .S1(n71)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(875[11] 878[52])
    defparam t_mult_24s_7s_0_add_3_10.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_10.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_10.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_10.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_11 (.A0(s_mult_24s_7s_0_2_25), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_26), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_10), .COUT(co_t_mult_24s_7s_0_3_11), 
          .S0(n70), .S1(n69)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(884[11] 887[52])
    defparam t_mult_24s_7s_0_add_3_11.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_11.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_11.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_11.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_12 (.A0(s_mult_24s_7s_0_2_27), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_28), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_11), .COUT(co_t_mult_24s_7s_0_3_12), 
          .S0(n68), .S1(n67)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(893[11] 896[52])
    defparam t_mult_24s_7s_0_add_3_12.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_12.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_12.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_12.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_13 (.A0(s_mult_24s_7s_0_2_29), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_30), .B1(GND_net), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_12), .S0(n66), 
          .S1(n65)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(902[11] 905[52])
    defparam t_mult_24s_7s_0_add_3_13.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_13.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_13.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_13.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_0 (.A0(GND_net), .B0(n123), .C0(GND_net), 
          .D0(n126), .A1(GND_net), .B1(n123), .C1(GND_net), .D1(n126), 
          .CIN(mult_24s_7s_0_cin_lr_0), .COUT(mco), .S0(\op_i_23__N_1310[1] ), 
          .S1(mult_24s_7s_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(911[11] 913[74])
    defparam mult_24s_7s_0_mult_0_0.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_0.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_0.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_0.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_1 (.A0(GND_net), .B0(n123), .C0(GND_net), 
          .D0(n126), .A1(GND_net), .B1(n123), .C1(GND_net), .D1(n126), 
          .CIN(mco), .COUT(mco_1), .S0(mult_24s_7s_0_pp_0_3), .S1(mult_24s_7s_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(919[11] 921[49])
    defparam mult_24s_7s_0_mult_0_1.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_1.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_1.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_1.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_2 (.A0(GND_net), .B0(n123), .C0(GND_net), 
          .D0(n126), .A1(GND_net), .B1(n123), .C1(GND_net), .D1(n126), 
          .CIN(mco_1), .COUT(mco_2), .S0(mult_24s_7s_0_pp_0_5), .S1(mult_24s_7s_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(927[11] 929[49])
    defparam mult_24s_7s_0_mult_0_2.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_2.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_3 (.A0(GND_net), .B0(n123), .C0(GND_net), 
          .D0(n126), .A1(GND_net), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_2), .COUT(mco_3), .S0(mult_24s_7s_0_pp_0_7), .S1(mult_24s_7s_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(935[11] 937[49])
    defparam mult_24s_7s_0_mult_0_3.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_3.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_3.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_3.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_4 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_3), .COUT(mco_4), .S0(mult_24s_7s_0_pp_0_9), .S1(mult_24s_7s_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(943[11] 945[50])
    defparam mult_24s_7s_0_mult_0_4.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_4.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_5 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_4), .COUT(mco_5), .S0(mult_24s_7s_0_pp_0_11), .S1(mult_24s_7s_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(951[11] 953[50])
    defparam mult_24s_7s_0_mult_0_5.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_5.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_5.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_5.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_6 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_5), .COUT(mco_6), .S0(mult_24s_7s_0_pp_0_13), .S1(mult_24s_7s_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(959[11] 961[50])
    defparam mult_24s_7s_0_mult_0_6.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_6.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_6.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_6.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_7 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_6), .COUT(mco_7), .S0(mult_24s_7s_0_pp_0_15), .S1(mult_24s_7s_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(967[11] 969[50])
    defparam mult_24s_7s_0_mult_0_7.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_7.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_7.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_7.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_8 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_7), .COUT(mco_8), .S0(mult_24s_7s_0_pp_0_17), .S1(mult_24s_7s_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(975[11] 977[50])
    defparam mult_24s_7s_0_mult_0_8.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_8.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_8.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_8.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_9 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_8), .COUT(mco_9), .S0(mult_24s_7s_0_pp_0_19), .S1(mult_24s_7s_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(983[11] 985[50])
    defparam mult_24s_7s_0_mult_0_9.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_9.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_9.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_9.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_10 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(n34795), .B1(n123), .C1(n34795), .D1(n126), 
          .CIN(mco_9), .COUT(mco_10), .S0(mult_24s_7s_0_pp_0_21), .S1(mult_24s_7s_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(991[11] 993[51])
    defparam mult_24s_7s_0_mult_0_10.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_10.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_10.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_10.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_11 (.A0(n34795), .B0(n123), .C0(n34795), 
          .D0(n126), .A1(mult_24s_7s_0_mult_0_11_n1), .B1(VCC_net), .C1(mult_24s_7s_0_mult_0_11_n3), 
          .D1(VCC_net), .CIN(mco_10), .COUT(mfco), .S0(mult_24s_7s_0_pp_0_23), 
          .S1(mult_24s_7s_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(999[11] 1002[49])
    defparam mult_24s_7s_0_mult_0_11.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_11.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_11.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_11.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_0 (.A0(GND_net), .B0(n117), .C0(GND_net), 
          .D0(n120), .A1(GND_net), .B1(n117), .C1(GND_net), .D1(n120), 
          .CIN(mult_24s_7s_0_cin_lr_2), .COUT(mco_11), .S0(mult_24s_7s_0_pp_1_3), 
          .S1(mult_24s_7s_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1008[11] 1010[77])
    defparam mult_24s_7s_0_mult_2_0.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_0.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_0.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_0.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_1 (.A0(GND_net), .B0(n117), .C0(GND_net), 
          .D0(n120), .A1(GND_net), .B1(n117), .C1(GND_net), .D1(n120), 
          .CIN(mco_11), .COUT(mco_12), .S0(mult_24s_7s_0_pp_1_5), .S1(mult_24s_7s_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1016[11] 1018[50])
    defparam mult_24s_7s_0_mult_2_1.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_1.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_1.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_1.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_2 (.A0(GND_net), .B0(n117), .C0(GND_net), 
          .D0(n120), .A1(GND_net), .B1(n117), .C1(GND_net), .D1(n120), 
          .CIN(mco_12), .COUT(mco_13), .S0(mult_24s_7s_0_pp_1_7), .S1(mult_24s_7s_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1024[11] 1026[50])
    defparam mult_24s_7s_0_mult_2_2.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_2.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_3 (.A0(GND_net), .B0(n117), .C0(GND_net), 
          .D0(n120), .A1(GND_net), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_13), .COUT(mco_14), .S0(mult_24s_7s_0_pp_1_9), .S1(mult_24s_7s_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1032[11] 1034[51])
    defparam mult_24s_7s_0_mult_2_3.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_3.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_3.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_3.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_4 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_14), .COUT(mco_15), .S0(mult_24s_7s_0_pp_1_11), .S1(mult_24s_7s_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1040[11] 1042[51])
    defparam mult_24s_7s_0_mult_2_4.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_4.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_5 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_15), .COUT(mco_16), .S0(mult_24s_7s_0_pp_1_13), .S1(mult_24s_7s_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1048[11] 1050[51])
    defparam mult_24s_7s_0_mult_2_5.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_5.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_5.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_5.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_6 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_16), .COUT(mco_17), .S0(mult_24s_7s_0_pp_1_15), .S1(mult_24s_7s_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1056[11] 1058[51])
    defparam mult_24s_7s_0_mult_2_6.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_6.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_6.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_6.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_7 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_17), .COUT(mco_18), .S0(mult_24s_7s_0_pp_1_17), .S1(mult_24s_7s_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1064[11] 1066[51])
    defparam mult_24s_7s_0_mult_2_7.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_7.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_7.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_7.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_8 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_18), .COUT(mco_19), .S0(mult_24s_7s_0_pp_1_19), .S1(mult_24s_7s_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1072[11] 1074[51])
    defparam mult_24s_7s_0_mult_2_8.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_8.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_8.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_8.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_9 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_19), .COUT(mco_20), .S0(mult_24s_7s_0_pp_1_21), .S1(mult_24s_7s_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1080[11] 1082[51])
    defparam mult_24s_7s_0_mult_2_9.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_9.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_9.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_9.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_10 (.A0(n34795), .B0(n117), .C0(n34795), 
          .D0(n120), .A1(n34795), .B1(n117), .C1(n34795), .D1(n120), 
          .CIN(mco_20), .COUT(mco_21), .S0(mult_24s_7s_0_pp_1_23), .S1(mult_24s_7s_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1088[11] 1090[51])
    defparam mult_24s_7s_0_mult_2_10.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_10.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_10.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_10.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_11 (.A0(n34795), .B0(n117), .C0(mult_24s_7s_0_mult_2_11_n2), 
          .D0(VCC_net), .A1(mult_24s_7s_0_mult_2_11_n1), .B1(VCC_net), 
          .C1(GND_net), .D1(n120), .CIN(mco_21), .COUT(mfco_1), .S0(mult_24s_7s_0_pp_1_25), 
          .S1(mult_24s_7s_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1096[11] 1099[51])
    defparam mult_24s_7s_0_mult_2_11.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_11.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_11.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_11.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_0 (.A0(GND_net), .B0(n111), .C0(GND_net), 
          .D0(n114), .A1(GND_net), .B1(n111), .C1(GND_net), .D1(n114), 
          .CIN(mult_24s_7s_0_cin_lr_4), .COUT(mco_22), .S0(mult_24s_7s_0_pp_2_5), 
          .S1(mult_24s_7s_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1105[11] 1107[77])
    defparam mult_24s_7s_0_mult_4_0.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_0.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_0.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_0.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_1 (.A0(GND_net), .B0(n111), .C0(GND_net), 
          .D0(n114), .A1(GND_net), .B1(n111), .C1(GND_net), .D1(n114), 
          .CIN(mco_22), .COUT(mco_23), .S0(mult_24s_7s_0_pp_2_7), .S1(mult_24s_7s_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1113[11] 1115[50])
    defparam mult_24s_7s_0_mult_4_1.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_1.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_1.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_1.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_2 (.A0(GND_net), .B0(n111), .C0(GND_net), 
          .D0(n114), .A1(GND_net), .B1(n111), .C1(GND_net), .D1(n114), 
          .CIN(mco_23), .COUT(mco_24), .S0(mult_24s_7s_0_pp_2_9), .S1(mult_24s_7s_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1121[11] 1123[51])
    defparam mult_24s_7s_0_mult_4_2.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_2.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_2.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_2.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_3 (.A0(GND_net), .B0(n111), .C0(GND_net), 
          .D0(n114), .A1(GND_net), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_24), .COUT(mco_25), .S0(mult_24s_7s_0_pp_2_11), .S1(mult_24s_7s_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1129[11] 1131[51])
    defparam mult_24s_7s_0_mult_4_3.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_3.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_3.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_3.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_4 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_25), .COUT(mco_26), .S0(mult_24s_7s_0_pp_2_13), .S1(mult_24s_7s_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1137[11] 1139[51])
    defparam mult_24s_7s_0_mult_4_4.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_4.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_4.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_4.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_5 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_26), .COUT(mco_27), .S0(mult_24s_7s_0_pp_2_15), .S1(mult_24s_7s_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1145[11] 1147[51])
    defparam mult_24s_7s_0_mult_4_5.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_5.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_5.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_5.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_6 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_27), .COUT(mco_28), .S0(mult_24s_7s_0_pp_2_17), .S1(mult_24s_7s_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1153[11] 1155[51])
    defparam mult_24s_7s_0_mult_4_6.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_6.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_6.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_6.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_7 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_28), .COUT(mco_29), .S0(mult_24s_7s_0_pp_2_19), .S1(mult_24s_7s_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1161[11] 1163[51])
    defparam mult_24s_7s_0_mult_4_7.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_7.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_7.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_7.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_8 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_29), .COUT(mco_30), .S0(mult_24s_7s_0_pp_2_21), .S1(mult_24s_7s_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1169[11] 1171[51])
    defparam mult_24s_7s_0_mult_4_8.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_8.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_8.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_8.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_9 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_30), .COUT(mco_31), .S0(mult_24s_7s_0_pp_2_23), .S1(mult_24s_7s_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1177[11] 1179[51])
    defparam mult_24s_7s_0_mult_4_9.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_9.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_9.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_9.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_10 (.A0(n34795), .B0(n111), .C0(n34795), 
          .D0(n114), .A1(n34795), .B1(n111), .C1(n34795), .D1(n114), 
          .CIN(mco_31), .COUT(mco_32), .S0(mult_24s_7s_0_pp_2_25), .S1(mult_24s_7s_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1185[11] 1187[51])
    defparam mult_24s_7s_0_mult_4_10.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_10.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_10.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_10.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_11 (.A0(n34795), .B0(n111), .C0(mult_24s_7s_0_mult_4_11_n2), 
          .D0(VCC_net), .A1(mult_24s_7s_0_mult_4_11_n1), .B1(VCC_net), 
          .C1(GND_net), .D1(n114), .CIN(mco_32), .COUT(mfco_2), .S0(mult_24s_7s_0_pp_2_27), 
          .S1(mult_24s_7s_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1197[11] 1200[51])
    defparam mult_24s_7s_0_mult_4_11.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_11.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_11.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_11.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_cin_lr_add_0 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(mult_24s_7s_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(367[11] 369[77])
    defparam mult_24s_7s_0_cin_lr_add_0.INIT0 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_0.INIT1 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_0.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_cin_lr_add_0.INJECT1_1 = "NO";
    ND2 ND2_t28_adj_39 (.A(\rom4_w_i[12] ), .B(n120_adj_34), .Z(mult_24s_7s_0_mult_2_11_n2_adj_6034)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t31_adj_40 (.A(\rom4_w_i[12] ), .B(n126_adj_35), .Z(mult_24s_7s_0_mult_0_11_n3_adj_6036)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t32_adj_41 (.A(n34777), .B(n126_adj_35), .Z(\op_i_23__N_1310[0]_adj_36 )) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(297[10:65])
    ND2 ND2_t30_adj_42 (.A(\rom4_w_i[12] ), .B(n123_adj_37), .Z(mult_24s_7s_0_mult_0_11_n1_adj_6039)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t29_adj_43 (.A(n34777), .B(n120_adj_34), .Z(mult_24s_7s_0_pp_1_2_adj_6040)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(303[10:65])
    ND2 ND2_t27_adj_44 (.A(\rom4_w_i[12] ), .B(n117_adj_38), .Z(mult_24s_7s_0_mult_2_11_n1_adj_6042)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t26_adj_45 (.A(n34777), .B(n114_adj_33), .Z(mult_24s_7s_0_pp_2_4_adj_6043)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(309[10:65])
    ND2 ND2_t24_adj_46 (.A(\rom4_w_i[12] ), .B(n111_adj_39), .Z(mult_24s_7s_0_mult_4_11_n1_adj_6045)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t23_adj_47 (.A(n34777), .B(GND_net), .Z(mult_24s_7s_0_pp_3_6_adj_6046)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t22_adj_48 (.A(n34777), .B(GND_net), .Z(mult_24s_7s_0_pp_3_7_adj_6047)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t21_adj_49 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_8_adj_6048)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t20_adj_50 (.A(n34777), .B(GND_net), .Z(mult_24s_7s_0_pp_3_9_adj_6049)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t19_adj_51 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_10_adj_6050)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t18_adj_52 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_11_adj_6051)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t17_adj_53 (.A(n34777), .B(GND_net), .Z(mult_24s_7s_0_pp_3_12_adj_6052)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t16_adj_54 (.A(GND_net), .B(GND_net), .Z(mult_24s_7s_0_pp_3_13_adj_6053)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t15_adj_55 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_14_adj_6054)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t14_adj_56 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_15_adj_6055)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t13_adj_57 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_16_adj_6056)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t12_adj_58 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_17_adj_6057)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t11_adj_59 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_18_adj_6058)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t10_adj_60 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_19_adj_6059)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t9_adj_61 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_20_adj_6060)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t8_adj_62 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_21_adj_6061)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t7_adj_63 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_22_adj_6062)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t6_adj_64 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_23_adj_6063)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t5_adj_65 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_24_adj_6064)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t4_adj_66 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_25_adj_6065)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t3_adj_67 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_26_adj_6066)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t2_adj_68 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_27_adj_6067)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t1_adj_69 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_28_adj_6068)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t0_adj_70 (.A(\rom4_w_i[12] ), .B(GND_net), .Z(mult_24s_7s_0_pp_3_29_adj_6069)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(361[10:66])
    CCU2C mult_24s_7s_0_Cadd_0_12_adj_71 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_adj_6071), .S0(mult_24s_7s_0_pp_0_25_adj_6070)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(375[11] 377[80])
    defparam mult_24s_7s_0_Cadd_0_12_adj_71.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_0_12_adj_71.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_0_12_adj_71.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_Cadd_0_12_adj_71.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_cin_lr_add_2_adj_72 (.A0(VCC_net), .B0(VCC_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(mult_24s_7s_0_cin_lr_2_adj_6072)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(383[11] 385[77])
    defparam mult_24s_7s_0_cin_lr_add_2_adj_72.INIT0 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_2_adj_72.INIT1 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_2_adj_72.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_cin_lr_add_2_adj_72.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_Cadd_2_12_adj_73 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_1_adj_6074), .S0(mult_24s_7s_0_pp_1_27_adj_6073)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(391[11] 394[17])
    defparam mult_24s_7s_0_Cadd_2_12_adj_73.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_2_12_adj_73.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_2_12_adj_73.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_Cadd_2_12_adj_73.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_cin_lr_add_4_adj_74 (.A0(VCC_net), .B0(VCC_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(mult_24s_7s_0_cin_lr_4_adj_6075)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(400[11] 402[77])
    defparam mult_24s_7s_0_cin_lr_add_4_adj_74.INIT0 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_4_adj_74.INIT1 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_4_adj_74.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_cin_lr_add_4_adj_74.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_Cadd_4_12_adj_75 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_2_adj_6077), .S0(mult_24s_7s_0_pp_2_29_adj_6076)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(408[11] 411[17])
    defparam mult_24s_7s_0_Cadd_4_12_adj_75.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_4_12_adj_75.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_Cadd_4_12_adj_75.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_Cadd_4_12_adj_75.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_0_1_adj_76 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(mult_24s_7s_0_pp_0_2_adj_6080), .B1(mult_24s_7s_0_pp_1_2_adj_6040), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_mult_24s_7s_0_0_1_adj_6079), 
          .S1(\op_i_23__N_1310[2]_adj_40 )) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(417[11] 420[37])
    defparam Cadd_mult_24s_7s_0_0_1_adj_76.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_1_adj_76.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_1_adj_76.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_0_1_adj_76.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_2_adj_77 (.A0(mult_24s_7s_0_pp_0_3_adj_6085), 
          .B0(mult_24s_7s_0_pp_1_3_adj_6087), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_4_adj_6084), .B1(mult_24s_7s_0_pp_1_4_adj_6086), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_1_adj_6079), 
          .COUT(co_mult_24s_7s_0_0_2_adj_6082), .S0(\op_i_23__N_1310[3]_adj_41 ), 
          .S1(s_mult_24s_7s_0_0_4_adj_6083)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(426[11] 429[89])
    defparam mult_24s_7s_0_add_0_2_adj_77.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_2_adj_77.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_2_adj_77.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_2_adj_77.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_3_adj_78 (.A0(mult_24s_7s_0_pp_0_5_adj_6092), 
          .B0(mult_24s_7s_0_pp_1_5_adj_6094), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_6_adj_6091), .B1(mult_24s_7s_0_pp_1_6_adj_6093), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_2_adj_6082), 
          .COUT(co_mult_24s_7s_0_0_3_adj_6088), .S0(s_mult_24s_7s_0_0_5_adj_6090), 
          .S1(s_mult_24s_7s_0_0_6_adj_6089)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(435[11] 438[89])
    defparam mult_24s_7s_0_add_0_3_adj_78.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_3_adj_78.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_3_adj_78.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_3_adj_78.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_4_adj_79 (.A0(mult_24s_7s_0_pp_0_7_adj_6099), 
          .B0(mult_24s_7s_0_pp_1_7_adj_6101), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_8_adj_6098), .B1(mult_24s_7s_0_pp_1_8_adj_6100), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_3_adj_6088), 
          .COUT(co_mult_24s_7s_0_0_4_adj_6095), .S0(s_mult_24s_7s_0_0_7_adj_6097), 
          .S1(s_mult_24s_7s_0_0_8_adj_6096)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(444[11] 447[89])
    defparam mult_24s_7s_0_add_0_4_adj_79.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_4_adj_79.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_4_adj_79.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_4_adj_79.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_5_adj_80 (.A0(mult_24s_7s_0_pp_0_9_adj_6106), 
          .B0(mult_24s_7s_0_pp_1_9_adj_6108), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_10_adj_6105), .B1(mult_24s_7s_0_pp_1_10_adj_6107), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_4_adj_6095), 
          .COUT(co_mult_24s_7s_0_0_5_adj_6102), .S0(s_mult_24s_7s_0_0_9_adj_6104), 
          .S1(s_mult_24s_7s_0_0_10_adj_6103)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(453[11] 456[90])
    defparam mult_24s_7s_0_add_0_5_adj_80.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_5_adj_80.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_5_adj_80.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_5_adj_80.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_6_adj_81 (.A0(mult_24s_7s_0_pp_0_11_adj_6113), 
          .B0(mult_24s_7s_0_pp_1_11_adj_6115), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_12_adj_6112), .B1(mult_24s_7s_0_pp_1_12_adj_6114), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_5_adj_6102), 
          .COUT(co_mult_24s_7s_0_0_6_adj_6109), .S0(s_mult_24s_7s_0_0_11_adj_6111), 
          .S1(s_mult_24s_7s_0_0_12_adj_6110)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(462[11] 465[91])
    defparam mult_24s_7s_0_add_0_6_adj_81.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_6_adj_81.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_6_adj_81.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_6_adj_81.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_7_adj_82 (.A0(mult_24s_7s_0_pp_0_13_adj_6120), 
          .B0(mult_24s_7s_0_pp_1_13_adj_6122), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_14_adj_6119), .B1(mult_24s_7s_0_pp_1_14_adj_6121), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_6_adj_6109), 
          .COUT(co_mult_24s_7s_0_0_7_adj_6116), .S0(s_mult_24s_7s_0_0_13_adj_6118), 
          .S1(s_mult_24s_7s_0_0_14_adj_6117)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(471[11] 474[91])
    defparam mult_24s_7s_0_add_0_7_adj_82.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_7_adj_82.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_7_adj_82.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_7_adj_82.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_8_adj_83 (.A0(mult_24s_7s_0_pp_0_15_adj_6127), 
          .B0(mult_24s_7s_0_pp_1_15_adj_6129), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_16_adj_6126), .B1(mult_24s_7s_0_pp_1_16_adj_6128), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_7_adj_6116), 
          .COUT(co_mult_24s_7s_0_0_8_adj_6123), .S0(s_mult_24s_7s_0_0_15_adj_6125), 
          .S1(s_mult_24s_7s_0_0_16_adj_6124)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(480[11] 483[91])
    defparam mult_24s_7s_0_add_0_8_adj_83.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_8_adj_83.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_8_adj_83.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_8_adj_83.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_9_adj_84 (.A0(mult_24s_7s_0_pp_0_17_adj_6134), 
          .B0(mult_24s_7s_0_pp_1_17_adj_6136), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_18_adj_6133), .B1(mult_24s_7s_0_pp_1_18_adj_6135), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_8_adj_6123), 
          .COUT(co_mult_24s_7s_0_0_9_adj_6130), .S0(s_mult_24s_7s_0_0_17_adj_6132), 
          .S1(s_mult_24s_7s_0_0_18_adj_6131)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(489[11] 492[91])
    defparam mult_24s_7s_0_add_0_9_adj_84.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_9_adj_84.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_9_adj_84.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_9_adj_84.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_10_adj_85 (.A0(mult_24s_7s_0_pp_0_19_adj_6141), 
          .B0(mult_24s_7s_0_pp_1_19_adj_6143), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_20_adj_6140), .B1(mult_24s_7s_0_pp_1_20_adj_6142), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_9_adj_6130), 
          .COUT(co_mult_24s_7s_0_0_10_adj_6137), .S0(s_mult_24s_7s_0_0_19_adj_6139), 
          .S1(s_mult_24s_7s_0_0_20_adj_6138)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(498[11] 501[92])
    defparam mult_24s_7s_0_add_0_10_adj_85.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_10_adj_85.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_10_adj_85.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_10_adj_85.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_11_adj_86 (.A0(mult_24s_7s_0_pp_0_21_adj_6148), 
          .B0(mult_24s_7s_0_pp_1_21_adj_6150), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_22_adj_6147), .B1(mult_24s_7s_0_pp_1_22_adj_6149), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_10_adj_6137), 
          .COUT(co_mult_24s_7s_0_0_11_adj_6144), .S0(s_mult_24s_7s_0_0_21_adj_6146), 
          .S1(s_mult_24s_7s_0_0_22_adj_6145)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(507[11] 510[92])
    defparam mult_24s_7s_0_add_0_11_adj_86.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_11_adj_86.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_11_adj_86.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_11_adj_86.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_12_adj_87 (.A0(mult_24s_7s_0_pp_0_23_adj_6155), 
          .B0(mult_24s_7s_0_pp_1_23_adj_6157), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_0_24_adj_6154), .B1(mult_24s_7s_0_pp_1_24_adj_6156), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_11_adj_6144), 
          .COUT(co_mult_24s_7s_0_0_12_adj_6151), .S0(s_mult_24s_7s_0_0_23_adj_6153), 
          .S1(s_mult_24s_7s_0_0_24_adj_6152)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(516[11] 519[92])
    defparam mult_24s_7s_0_add_0_12_adj_87.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_12_adj_87.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_12_adj_87.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_12_adj_87.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_13_adj_88 (.A0(mult_24s_7s_0_pp_0_25_adj_6070), 
          .B0(mult_24s_7s_0_pp_1_25_adj_6162), .C0(VCC_net), .D0(VCC_net), 
          .A1(GND_net), .B1(mult_24s_7s_0_pp_1_26_adj_6161), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_12_adj_6151), .COUT(co_mult_24s_7s_0_0_13_adj_6158), 
          .S0(s_mult_24s_7s_0_0_25_adj_6160), .S1(s_mult_24s_7s_0_0_26_adj_6159)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(525[11] 528[92])
    defparam mult_24s_7s_0_add_0_13_adj_88.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_13_adj_88.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_13_adj_88.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_13_adj_88.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_0_14_adj_89 (.A0(GND_net), .B0(mult_24s_7s_0_pp_1_27_adj_6073), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_mult_24s_7s_0_0_13_adj_6158), .COUT(co_mult_24s_7s_0_0_14_adj_6163), 
          .S0(s_mult_24s_7s_0_0_27_adj_6165), .S1(s_mult_24s_7s_0_0_28_adj_6164)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(534[11] 537[65])
    defparam mult_24s_7s_0_add_0_14_adj_89.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_14_adj_89.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_0_14_adj_89.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_0_14_adj_89.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_0_15_adj_90 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_mult_24s_7s_0_0_14_adj_6163), .S0(s_mult_24s_7s_0_0_29_adj_6166)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(543[11] 546[24])
    defparam Cadd_mult_24s_7s_0_0_15_adj_90.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_15_adj_90.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_0_15_adj_90.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_0_15_adj_90.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_1_1_adj_91 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(mult_24s_7s_0_pp_2_6_adj_6169), .B1(mult_24s_7s_0_pp_3_6_adj_6046), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_mult_24s_7s_0_1_1_adj_6167), 
          .S1(s_mult_24s_7s_0_1_6_adj_6168)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(552[11] 555[37])
    defparam Cadd_mult_24s_7s_0_1_1_adj_91.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_1_1_adj_91.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_1_1_adj_91.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_1_1_adj_91.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_2_adj_92 (.A0(mult_24s_7s_0_pp_2_7_adj_6174), 
          .B0(mult_24s_7s_0_pp_3_7_adj_6047), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_8_adj_6173), .B1(mult_24s_7s_0_pp_3_8_adj_6048), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_1_adj_6167), 
          .COUT(co_mult_24s_7s_0_1_2_adj_6170), .S0(s_mult_24s_7s_0_1_7_adj_6172), 
          .S1(s_mult_24s_7s_0_1_8_adj_6171)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(561[11] 564[89])
    defparam mult_24s_7s_0_add_1_2_adj_92.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_2_adj_92.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_2_adj_92.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_2_adj_92.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_3_adj_93 (.A0(mult_24s_7s_0_pp_2_9_adj_6179), 
          .B0(mult_24s_7s_0_pp_3_9_adj_6049), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_10_adj_6178), .B1(mult_24s_7s_0_pp_3_10_adj_6050), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_2_adj_6170), 
          .COUT(co_mult_24s_7s_0_1_3_adj_6175), .S0(s_mult_24s_7s_0_1_9_adj_6177), 
          .S1(s_mult_24s_7s_0_1_10_adj_6176)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(570[11] 573[90])
    defparam mult_24s_7s_0_add_1_3_adj_93.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_3_adj_93.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_3_adj_93.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_3_adj_93.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_4_adj_94 (.A0(mult_24s_7s_0_pp_2_11_adj_6184), 
          .B0(mult_24s_7s_0_pp_3_11_adj_6051), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_12_adj_6183), .B1(mult_24s_7s_0_pp_3_12_adj_6052), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_3_adj_6175), 
          .COUT(co_mult_24s_7s_0_1_4_adj_6180), .S0(s_mult_24s_7s_0_1_11_adj_6182), 
          .S1(s_mult_24s_7s_0_1_12_adj_6181)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(579[11] 582[91])
    defparam mult_24s_7s_0_add_1_4_adj_94.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_4_adj_94.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_4_adj_94.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_4_adj_94.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_5_adj_95 (.A0(mult_24s_7s_0_pp_2_13_adj_6189), 
          .B0(mult_24s_7s_0_pp_3_13_adj_6053), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_14_adj_6188), .B1(mult_24s_7s_0_pp_3_14_adj_6054), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_4_adj_6180), 
          .COUT(co_mult_24s_7s_0_1_5_adj_6185), .S0(s_mult_24s_7s_0_1_13_adj_6187), 
          .S1(s_mult_24s_7s_0_1_14_adj_6186)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(588[11] 591[91])
    defparam mult_24s_7s_0_add_1_5_adj_95.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_5_adj_95.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_5_adj_95.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_5_adj_95.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_6_adj_96 (.A0(mult_24s_7s_0_pp_2_15_adj_6194), 
          .B0(mult_24s_7s_0_pp_3_15_adj_6055), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_16_adj_6193), .B1(mult_24s_7s_0_pp_3_16_adj_6056), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_5_adj_6185), 
          .COUT(co_mult_24s_7s_0_1_6_adj_6190), .S0(s_mult_24s_7s_0_1_15_adj_6192), 
          .S1(s_mult_24s_7s_0_1_16_adj_6191)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(597[11] 600[91])
    defparam mult_24s_7s_0_add_1_6_adj_96.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_6_adj_96.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_6_adj_96.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_6_adj_96.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_7_adj_97 (.A0(mult_24s_7s_0_pp_2_17_adj_6199), 
          .B0(mult_24s_7s_0_pp_3_17_adj_6057), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_18_adj_6198), .B1(mult_24s_7s_0_pp_3_18_adj_6058), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_6_adj_6190), 
          .COUT(co_mult_24s_7s_0_1_7_adj_6195), .S0(s_mult_24s_7s_0_1_17_adj_6197), 
          .S1(s_mult_24s_7s_0_1_18_adj_6196)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(606[11] 609[91])
    defparam mult_24s_7s_0_add_1_7_adj_97.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_7_adj_97.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_7_adj_97.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_7_adj_97.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_8_adj_98 (.A0(mult_24s_7s_0_pp_2_19_adj_6204), 
          .B0(mult_24s_7s_0_pp_3_19_adj_6059), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_20_adj_6203), .B1(mult_24s_7s_0_pp_3_20_adj_6060), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_7_adj_6195), 
          .COUT(co_mult_24s_7s_0_1_8_adj_6200), .S0(s_mult_24s_7s_0_1_19_adj_6202), 
          .S1(s_mult_24s_7s_0_1_20_adj_6201)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(615[11] 618[91])
    defparam mult_24s_7s_0_add_1_8_adj_98.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_8_adj_98.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_8_adj_98.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_8_adj_98.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_9_adj_99 (.A0(mult_24s_7s_0_pp_2_21_adj_6209), 
          .B0(mult_24s_7s_0_pp_3_21_adj_6061), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_22_adj_6208), .B1(mult_24s_7s_0_pp_3_22_adj_6062), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_8_adj_6200), 
          .COUT(co_mult_24s_7s_0_1_9_adj_6205), .S0(s_mult_24s_7s_0_1_21_adj_6207), 
          .S1(s_mult_24s_7s_0_1_22_adj_6206)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(624[11] 627[91])
    defparam mult_24s_7s_0_add_1_9_adj_99.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_9_adj_99.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_9_adj_99.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_9_adj_99.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_10_adj_100 (.A0(mult_24s_7s_0_pp_2_23_adj_6214), 
          .B0(mult_24s_7s_0_pp_3_23_adj_6063), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_24_adj_6213), .B1(mult_24s_7s_0_pp_3_24_adj_6064), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_9_adj_6205), 
          .COUT(co_mult_24s_7s_0_1_10_adj_6210), .S0(s_mult_24s_7s_0_1_23_adj_6212), 
          .S1(s_mult_24s_7s_0_1_24_adj_6211)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(633[11] 636[92])
    defparam mult_24s_7s_0_add_1_10_adj_100.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_10_adj_100.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_10_adj_100.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_10_adj_100.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_11_adj_101 (.A0(mult_24s_7s_0_pp_2_25_adj_6219), 
          .B0(mult_24s_7s_0_pp_3_25_adj_6065), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_26_adj_6218), .B1(mult_24s_7s_0_pp_3_26_adj_6066), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_10_adj_6210), 
          .COUT(co_mult_24s_7s_0_1_11_adj_6215), .S0(s_mult_24s_7s_0_1_25_adj_6217), 
          .S1(s_mult_24s_7s_0_1_26_adj_6216)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(642[11] 645[92])
    defparam mult_24s_7s_0_add_1_11_adj_101.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_11_adj_101.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_11_adj_101.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_11_adj_101.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_12_adj_102 (.A0(mult_24s_7s_0_pp_2_27_adj_6224), 
          .B0(mult_24s_7s_0_pp_3_27_adj_6067), .C0(VCC_net), .D0(VCC_net), 
          .A1(mult_24s_7s_0_pp_2_28_adj_6223), .B1(mult_24s_7s_0_pp_3_28_adj_6068), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_11_adj_6215), 
          .COUT(co_mult_24s_7s_0_1_12_adj_6220), .S0(s_mult_24s_7s_0_1_27_adj_6222), 
          .S1(s_mult_24s_7s_0_1_28_adj_6221)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(651[11] 654[92])
    defparam mult_24s_7s_0_add_1_12_adj_102.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_12_adj_102.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_12_adj_102.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_12_adj_102.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_1_13_adj_103 (.A0(mult_24s_7s_0_pp_2_29_adj_6076), 
          .B0(mult_24s_7s_0_pp_3_29_adj_6069), .C0(VCC_net), .D0(VCC_net), 
          .A1(GND_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_1_12_adj_6220), 
          .S0(s_mult_24s_7s_0_1_29_adj_6226), .S1(s_mult_24s_7s_0_1_30_adj_6225)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(660[11] 663[65])
    defparam mult_24s_7s_0_add_1_13_adj_103.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_13_adj_103.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_1_13_adj_103.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_1_13_adj_103.INJECT1_1 = "NO";
    CCU2C Cadd_mult_24s_7s_0_2_1_adj_104 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(s_mult_24s_7s_0_0_4_adj_6083), .B1(mult_24s_7s_0_pp_2_4_adj_6043), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_mult_24s_7s_0_2_1_adj_6228), 
          .S1(\op_i_23__N_1310[4]_adj_42 )) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(669[11] 672[37])
    defparam Cadd_mult_24s_7s_0_2_1_adj_104.INIT0 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_2_1_adj_104.INIT1 = 16'b0110011010101010;
    defparam Cadd_mult_24s_7s_0_2_1_adj_104.INJECT1_0 = "NO";
    defparam Cadd_mult_24s_7s_0_2_1_adj_104.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_2_adj_105 (.A0(s_mult_24s_7s_0_0_5_adj_6090), 
          .B0(mult_24s_7s_0_pp_2_5_adj_6232), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_6_adj_6089), .B1(s_mult_24s_7s_0_1_6_adj_6168), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_1_adj_6228), 
          .COUT(co_mult_24s_7s_0_2_2_adj_6230), .S0(\op_i_23__N_1310[5]_adj_43 ), 
          .S1(s_mult_24s_7s_0_2_6_adj_6231)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(678[11] 681[89])
    defparam mult_24s_7s_0_add_2_2_adj_105.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_2_adj_105.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_2_adj_105.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_2_adj_105.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_3_adj_106 (.A0(s_mult_24s_7s_0_0_7_adj_6097), 
          .B0(s_mult_24s_7s_0_1_7_adj_6172), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_8_adj_6096), .B1(s_mult_24s_7s_0_1_8_adj_6171), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_2_adj_6230), 
          .COUT(co_mult_24s_7s_0_2_3_adj_6233), .S0(s_mult_24s_7s_0_2_7_adj_6235), 
          .S1(s_mult_24s_7s_0_2_8_adj_6234)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(687[11] 690[89])
    defparam mult_24s_7s_0_add_2_3_adj_106.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_3_adj_106.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_3_adj_106.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_3_adj_106.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_4_adj_107 (.A0(s_mult_24s_7s_0_0_9_adj_6104), 
          .B0(s_mult_24s_7s_0_1_9_adj_6177), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_10_adj_6103), .B1(s_mult_24s_7s_0_1_10_adj_6176), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_3_adj_6233), 
          .COUT(co_mult_24s_7s_0_2_4_adj_6236), .S0(s_mult_24s_7s_0_2_9_adj_6238), 
          .S1(s_mult_24s_7s_0_2_10_adj_6237)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(696[11] 699[90])
    defparam mult_24s_7s_0_add_2_4_adj_107.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_4_adj_107.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_4_adj_107.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_4_adj_107.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_5_adj_108 (.A0(s_mult_24s_7s_0_0_11_adj_6111), 
          .B0(s_mult_24s_7s_0_1_11_adj_6182), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_12_adj_6110), .B1(s_mult_24s_7s_0_1_12_adj_6181), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_4_adj_6236), 
          .COUT(co_mult_24s_7s_0_2_5_adj_6239), .S0(s_mult_24s_7s_0_2_11_adj_6241), 
          .S1(s_mult_24s_7s_0_2_12_adj_6240)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(705[11] 708[91])
    defparam mult_24s_7s_0_add_2_5_adj_108.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_5_adj_108.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_5_adj_108.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_5_adj_108.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_6_adj_109 (.A0(s_mult_24s_7s_0_0_13_adj_6118), 
          .B0(s_mult_24s_7s_0_1_13_adj_6187), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_14_adj_6117), .B1(s_mult_24s_7s_0_1_14_adj_6186), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_5_adj_6239), 
          .COUT(co_mult_24s_7s_0_2_6_adj_6242), .S0(s_mult_24s_7s_0_2_13_adj_6244), 
          .S1(s_mult_24s_7s_0_2_14_adj_6243)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(714[11] 717[91])
    defparam mult_24s_7s_0_add_2_6_adj_109.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_6_adj_109.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_6_adj_109.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_6_adj_109.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_7_adj_110 (.A0(s_mult_24s_7s_0_0_15_adj_6125), 
          .B0(s_mult_24s_7s_0_1_15_adj_6192), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_16_adj_6124), .B1(s_mult_24s_7s_0_1_16_adj_6191), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_6_adj_6242), 
          .COUT(co_mult_24s_7s_0_2_7_adj_6245), .S0(s_mult_24s_7s_0_2_15_adj_6247), 
          .S1(s_mult_24s_7s_0_2_16_adj_6246)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(723[11] 726[91])
    defparam mult_24s_7s_0_add_2_7_adj_110.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_7_adj_110.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_7_adj_110.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_7_adj_110.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_8_adj_111 (.A0(s_mult_24s_7s_0_0_17_adj_6132), 
          .B0(s_mult_24s_7s_0_1_17_adj_6197), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_18_adj_6131), .B1(s_mult_24s_7s_0_1_18_adj_6196), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_7_adj_6245), 
          .COUT(co_mult_24s_7s_0_2_8_adj_6248), .S0(s_mult_24s_7s_0_2_17_adj_6250), 
          .S1(s_mult_24s_7s_0_2_18_adj_6249)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(732[11] 735[91])
    defparam mult_24s_7s_0_add_2_8_adj_111.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_8_adj_111.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_8_adj_111.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_8_adj_111.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_9_adj_112 (.A0(s_mult_24s_7s_0_0_19_adj_6139), 
          .B0(s_mult_24s_7s_0_1_19_adj_6202), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_20_adj_6138), .B1(s_mult_24s_7s_0_1_20_adj_6201), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_8_adj_6248), 
          .COUT(co_mult_24s_7s_0_2_9_adj_6251), .S0(s_mult_24s_7s_0_2_19_adj_6253), 
          .S1(s_mult_24s_7s_0_2_20_adj_6252)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(741[11] 744[91])
    defparam mult_24s_7s_0_add_2_9_adj_112.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_9_adj_112.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_9_adj_112.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_9_adj_112.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_10_adj_113 (.A0(s_mult_24s_7s_0_0_21_adj_6146), 
          .B0(s_mult_24s_7s_0_1_21_adj_6207), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_22_adj_6145), .B1(s_mult_24s_7s_0_1_22_adj_6206), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_9_adj_6251), 
          .COUT(co_mult_24s_7s_0_2_10_adj_6254), .S0(s_mult_24s_7s_0_2_21_adj_6256), 
          .S1(s_mult_24s_7s_0_2_22_adj_6255)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(750[11] 753[92])
    defparam mult_24s_7s_0_add_2_10_adj_113.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_10_adj_113.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_10_adj_113.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_10_adj_113.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_11_adj_114 (.A0(s_mult_24s_7s_0_0_23_adj_6153), 
          .B0(s_mult_24s_7s_0_1_23_adj_6212), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_24_adj_6152), .B1(s_mult_24s_7s_0_1_24_adj_6211), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_10_adj_6254), 
          .COUT(co_mult_24s_7s_0_2_11_adj_6257), .S0(s_mult_24s_7s_0_2_23_adj_6259), 
          .S1(s_mult_24s_7s_0_2_24_adj_6258)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(759[11] 762[92])
    defparam mult_24s_7s_0_add_2_11_adj_114.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_11_adj_114.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_11_adj_114.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_11_adj_114.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_12_adj_115 (.A0(s_mult_24s_7s_0_0_25_adj_6160), 
          .B0(s_mult_24s_7s_0_1_25_adj_6217), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_26_adj_6159), .B1(s_mult_24s_7s_0_1_26_adj_6216), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_11_adj_6257), 
          .COUT(co_mult_24s_7s_0_2_12_adj_6260), .S0(s_mult_24s_7s_0_2_25_adj_6262), 
          .S1(s_mult_24s_7s_0_2_26_adj_6261)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(768[11] 771[92])
    defparam mult_24s_7s_0_add_2_12_adj_115.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_12_adj_115.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_12_adj_115.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_12_adj_115.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_13_adj_116 (.A0(s_mult_24s_7s_0_0_27_adj_6165), 
          .B0(s_mult_24s_7s_0_1_27_adj_6222), .C0(VCC_net), .D0(VCC_net), 
          .A1(s_mult_24s_7s_0_0_28_adj_6164), .B1(s_mult_24s_7s_0_1_28_adj_6221), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_12_adj_6260), 
          .COUT(co_mult_24s_7s_0_2_13_adj_6263), .S0(s_mult_24s_7s_0_2_27_adj_6265), 
          .S1(s_mult_24s_7s_0_2_28_adj_6264)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(777[11] 780[92])
    defparam mult_24s_7s_0_add_2_13_adj_116.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_13_adj_116.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_13_adj_116.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_13_adj_116.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_add_2_14_adj_117 (.A0(s_mult_24s_7s_0_0_29_adj_6166), 
          .B0(s_mult_24s_7s_0_1_29_adj_6226), .C0(VCC_net), .D0(VCC_net), 
          .A1(GND_net), .B1(s_mult_24s_7s_0_1_30_adj_6225), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_mult_24s_7s_0_2_13_adj_6263), .S0(s_mult_24s_7s_0_2_29_adj_6267), 
          .S1(s_mult_24s_7s_0_2_30_adj_6266)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(786[11] 789[92])
    defparam mult_24s_7s_0_add_2_14_adj_117.INIT0 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_14_adj_117.INIT1 = 16'b0110011010101010;
    defparam mult_24s_7s_0_add_2_14_adj_117.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_add_2_14_adj_117.INJECT1_1 = "NO";
    CCU2C Cadd_t_mult_24s_7s_0_3_1_adj_118 (.A0(GND_net), .B0(GND_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_6_adj_6231), 
          .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), .COUT(co_t_mult_24s_7s_0_3_1_adj_6269), 
          .S1(n89_adj_44)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(795[11] 797[97])
    defparam Cadd_t_mult_24s_7s_0_3_1_adj_118.INIT0 = 16'b0110011010101010;
    defparam Cadd_t_mult_24s_7s_0_3_1_adj_118.INIT1 = 16'b0110011010101010;
    defparam Cadd_t_mult_24s_7s_0_3_1_adj_118.INJECT1_0 = "NO";
    defparam Cadd_t_mult_24s_7s_0_3_1_adj_118.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_2_adj_119 (.A0(s_mult_24s_7s_0_2_7_adj_6235), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_8_adj_6234), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_1_adj_6269), 
          .COUT(co_t_mult_24s_7s_0_3_2_adj_6272), .S0(n88_adj_46), .S1(n87_adj_45)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(803[11] 806[50])
    defparam t_mult_24s_7s_0_add_3_2_adj_119.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_2_adj_119.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_2_adj_119.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_2_adj_119.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_3_adj_120 (.A0(s_mult_24s_7s_0_2_9_adj_6238), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_10_adj_6237), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_2_adj_6272), 
          .COUT(co_t_mult_24s_7s_0_3_3_adj_6275), .S0(n86_adj_48), .S1(n85_adj_47)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(812[11] 815[51])
    defparam t_mult_24s_7s_0_add_3_3_adj_120.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_3_adj_120.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_3_adj_120.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_3_adj_120.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_4_adj_121 (.A0(s_mult_24s_7s_0_2_11_adj_6241), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_12_adj_6240), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_3_adj_6275), 
          .COUT(co_t_mult_24s_7s_0_3_4_adj_6278), .S0(n84_adj_50), .S1(n83_adj_49)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(821[11] 824[51])
    defparam t_mult_24s_7s_0_add_3_4_adj_121.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_4_adj_121.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_4_adj_121.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_4_adj_121.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_5_adj_122 (.A0(s_mult_24s_7s_0_2_13_adj_6244), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_14_adj_6243), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_4_adj_6278), 
          .COUT(co_t_mult_24s_7s_0_3_5_adj_6281), .S0(n82_adj_52), .S1(n81_adj_51)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(830[11] 833[51])
    defparam t_mult_24s_7s_0_add_3_5_adj_122.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_5_adj_122.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_5_adj_122.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_5_adj_122.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_6_adj_123 (.A0(s_mult_24s_7s_0_2_15_adj_6247), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_16_adj_6246), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_5_adj_6281), 
          .COUT(co_t_mult_24s_7s_0_3_6_adj_6284), .S0(n80_adj_54), .S1(n79_adj_53)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(839[11] 842[51])
    defparam t_mult_24s_7s_0_add_3_6_adj_123.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_6_adj_123.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_6_adj_123.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_6_adj_123.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_7_adj_124 (.A0(s_mult_24s_7s_0_2_17_adj_6250), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_18_adj_6249), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_6_adj_6284), 
          .COUT(co_t_mult_24s_7s_0_3_7_adj_6287), .S0(n78_adj_56), .S1(n77_adj_55)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(848[11] 851[51])
    defparam t_mult_24s_7s_0_add_3_7_adj_124.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_7_adj_124.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_7_adj_124.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_7_adj_124.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_8_adj_125 (.A0(s_mult_24s_7s_0_2_19_adj_6253), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_20_adj_6252), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_7_adj_6287), 
          .COUT(co_t_mult_24s_7s_0_3_8_adj_6290), .S0(n76_adj_58), .S1(n75_adj_57)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(857[11] 860[51])
    defparam t_mult_24s_7s_0_add_3_8_adj_125.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_8_adj_125.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_8_adj_125.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_8_adj_125.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_9_adj_126 (.A0(s_mult_24s_7s_0_2_21_adj_6256), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_22_adj_6255), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_8_adj_6290), 
          .COUT(co_t_mult_24s_7s_0_3_9_adj_6293), .S0(n74_adj_60), .S1(n73_adj_59)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(866[11] 869[51])
    defparam t_mult_24s_7s_0_add_3_9_adj_126.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_9_adj_126.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_9_adj_126.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_9_adj_126.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_10_adj_127 (.A0(s_mult_24s_7s_0_2_23_adj_6259), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_24_adj_6258), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_9_adj_6293), 
          .COUT(co_t_mult_24s_7s_0_3_10_adj_6296), .S0(n72_adj_62), .S1(n71_adj_61)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(875[11] 878[52])
    defparam t_mult_24s_7s_0_add_3_10_adj_127.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_10_adj_127.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_10_adj_127.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_10_adj_127.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_11_adj_128 (.A0(s_mult_24s_7s_0_2_25_adj_6262), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_26_adj_6261), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_10_adj_6296), 
          .COUT(co_t_mult_24s_7s_0_3_11_adj_6299), .S0(n70_adj_64), .S1(n69_adj_63)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(884[11] 887[52])
    defparam t_mult_24s_7s_0_add_3_11_adj_128.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_11_adj_128.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_11_adj_128.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_11_adj_128.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_12_adj_129 (.A0(s_mult_24s_7s_0_2_27_adj_6265), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_28_adj_6264), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_11_adj_6299), 
          .COUT(co_t_mult_24s_7s_0_3_12_adj_6302), .S0(n68_adj_66), .S1(n67_adj_65)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(893[11] 896[52])
    defparam t_mult_24s_7s_0_add_3_12_adj_129.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_12_adj_129.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_12_adj_129.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_12_adj_129.INJECT1_1 = "NO";
    CCU2C t_mult_24s_7s_0_add_3_13_adj_130 (.A0(s_mult_24s_7s_0_2_29_adj_6267), 
          .B0(GND_net), .C0(VCC_net), .D0(VCC_net), .A1(s_mult_24s_7s_0_2_30_adj_6266), 
          .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co_t_mult_24s_7s_0_3_12_adj_6302), 
          .S0(n66_adj_68), .S1(n65_adj_67)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(902[11] 905[52])
    defparam t_mult_24s_7s_0_add_3_13_adj_130.INIT0 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_13_adj_130.INIT1 = 16'b0110011010101010;
    defparam t_mult_24s_7s_0_add_3_13_adj_130.INJECT1_0 = "NO";
    defparam t_mult_24s_7s_0_add_3_13_adj_130.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_0_adj_131 (.A0(n34777), .B0(n123_adj_37), 
          .C0(n34777), .D0(n126_adj_35), .A1(n34777), .B1(n123_adj_37), 
          .C1(GND_net), .D1(n126_adj_35), .CIN(mult_24s_7s_0_cin_lr_0_adj_6306), 
          .COUT(mco_adj_6307), .S0(\op_i_23__N_1310[1]_adj_69 ), .S1(mult_24s_7s_0_pp_0_2_adj_6080)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(911[11] 913[74])
    defparam mult_24s_7s_0_mult_0_0_adj_131.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_0_adj_131.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_0_adj_131.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_0_adj_131.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_1_adj_132 (.A0(GND_net), .B0(n123_adj_37), 
          .C0(n34777), .D0(n126_adj_35), .A1(n34777), .B1(n123_adj_37), 
          .C1(GND_net), .D1(n126_adj_35), .CIN(mco_adj_6307), .COUT(mco_1_adj_6308), 
          .S0(mult_24s_7s_0_pp_0_3_adj_6085), .S1(mult_24s_7s_0_pp_0_4_adj_6084)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(919[11] 921[49])
    defparam mult_24s_7s_0_mult_0_1_adj_132.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_1_adj_132.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_1_adj_132.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_1_adj_132.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_2_adj_133 (.A0(GND_net), .B0(n123_adj_37), 
          .C0(GND_net), .D0(n126_adj_35), .A1(GND_net), .B1(n123_adj_37), 
          .C1(n34777), .D1(n126_adj_35), .CIN(mco_1_adj_6308), .COUT(mco_2_adj_6309), 
          .S0(mult_24s_7s_0_pp_0_5_adj_6092), .S1(mult_24s_7s_0_pp_0_6_adj_6091)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(927[11] 929[49])
    defparam mult_24s_7s_0_mult_0_2_adj_133.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_2_adj_133.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_2_adj_133.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_2_adj_133.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_3_adj_134 (.A0(n34777), .B0(n123_adj_37), 
          .C0(GND_net), .D0(n126_adj_35), .A1(GND_net), .B1(n123_adj_37), 
          .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_2_adj_6309), 
          .COUT(mco_3_adj_6310), .S0(mult_24s_7s_0_pp_0_7_adj_6099), .S1(mult_24s_7s_0_pp_0_8_adj_6098)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(935[11] 937[49])
    defparam mult_24s_7s_0_mult_0_3_adj_134.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_3_adj_134.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_3_adj_134.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_3_adj_134.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_4_adj_135 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_3_adj_6310), 
          .COUT(mco_4_adj_6311), .S0(mult_24s_7s_0_pp_0_9_adj_6106), .S1(mult_24s_7s_0_pp_0_10_adj_6105)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(943[11] 945[50])
    defparam mult_24s_7s_0_mult_0_4_adj_135.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_4_adj_135.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_4_adj_135.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_4_adj_135.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_5_adj_136 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_4_adj_6311), 
          .COUT(mco_5_adj_6312), .S0(mult_24s_7s_0_pp_0_11_adj_6113), .S1(mult_24s_7s_0_pp_0_12_adj_6112)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(951[11] 953[50])
    defparam mult_24s_7s_0_mult_0_5_adj_136.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_5_adj_136.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_5_adj_136.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_5_adj_136.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_6_adj_137 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_5_adj_6312), 
          .COUT(mco_6_adj_6313), .S0(mult_24s_7s_0_pp_0_13_adj_6120), .S1(mult_24s_7s_0_pp_0_14_adj_6119)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(959[11] 961[50])
    defparam mult_24s_7s_0_mult_0_6_adj_137.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_6_adj_137.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_6_adj_137.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_6_adj_137.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_7_adj_138 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_6_adj_6313), 
          .COUT(mco_7_adj_6314), .S0(mult_24s_7s_0_pp_0_15_adj_6127), .S1(mult_24s_7s_0_pp_0_16_adj_6126)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(967[11] 969[50])
    defparam mult_24s_7s_0_mult_0_7_adj_138.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_7_adj_138.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_7_adj_138.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_7_adj_138.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_8_adj_139 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_7_adj_6314), 
          .COUT(mco_8_adj_6315), .S0(mult_24s_7s_0_pp_0_17_adj_6134), .S1(mult_24s_7s_0_pp_0_18_adj_6133)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(975[11] 977[50])
    defparam mult_24s_7s_0_mult_0_8_adj_139.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_8_adj_139.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_8_adj_139.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_8_adj_139.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_9_adj_140 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_8_adj_6315), 
          .COUT(mco_9_adj_6316), .S0(mult_24s_7s_0_pp_0_19_adj_6141), .S1(mult_24s_7s_0_pp_0_20_adj_6140)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(983[11] 985[50])
    defparam mult_24s_7s_0_mult_0_9_adj_140.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_9_adj_140.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_9_adj_140.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_9_adj_140.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_10_adj_141 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(\rom4_w_i[12] ), 
          .B1(n123_adj_37), .C1(\rom4_w_i[12] ), .D1(n126_adj_35), .CIN(mco_9_adj_6316), 
          .COUT(mco_10_adj_6317), .S0(mult_24s_7s_0_pp_0_21_adj_6148), .S1(mult_24s_7s_0_pp_0_22_adj_6147)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(991[11] 993[51])
    defparam mult_24s_7s_0_mult_0_10_adj_141.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_10_adj_141.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_10_adj_141.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_10_adj_141.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_0_11_adj_142 (.A0(\rom4_w_i[12] ), .B0(n123_adj_37), 
          .C0(\rom4_w_i[12] ), .D0(n126_adj_35), .A1(mult_24s_7s_0_mult_0_11_n1_adj_6039), 
          .B1(VCC_net), .C1(mult_24s_7s_0_mult_0_11_n3_adj_6036), .D1(VCC_net), 
          .CIN(mco_10_adj_6317), .COUT(mfco_adj_6071), .S0(mult_24s_7s_0_pp_0_23_adj_6155), 
          .S1(mult_24s_7s_0_pp_0_24_adj_6154)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(999[11] 1002[49])
    defparam mult_24s_7s_0_mult_0_11_adj_142.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_11_adj_142.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_0_11_adj_142.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_0_11_adj_142.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_0_adj_143 (.A0(n34777), .B0(n117_adj_38), 
          .C0(n34777), .D0(n120_adj_34), .A1(n34777), .B1(n117_adj_38), 
          .C1(GND_net), .D1(n120_adj_34), .CIN(mult_24s_7s_0_cin_lr_2_adj_6072), 
          .COUT(mco_11_adj_6318), .S0(mult_24s_7s_0_pp_1_3_adj_6087), .S1(mult_24s_7s_0_pp_1_4_adj_6086)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1008[11] 1010[77])
    defparam mult_24s_7s_0_mult_2_0_adj_143.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_0_adj_143.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_0_adj_143.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_0_adj_143.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_1_adj_144 (.A0(GND_net), .B0(n117_adj_38), 
          .C0(n34777), .D0(n120_adj_34), .A1(n34777), .B1(n117_adj_38), 
          .C1(GND_net), .D1(n120_adj_34), .CIN(mco_11_adj_6318), .COUT(mco_12_adj_6319), 
          .S0(mult_24s_7s_0_pp_1_5_adj_6094), .S1(mult_24s_7s_0_pp_1_6_adj_6093)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1016[11] 1018[50])
    defparam mult_24s_7s_0_mult_2_1_adj_144.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_1_adj_144.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_1_adj_144.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_1_adj_144.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_2_adj_145 (.A0(GND_net), .B0(n117_adj_38), 
          .C0(GND_net), .D0(n120_adj_34), .A1(GND_net), .B1(n117_adj_38), 
          .C1(n34777), .D1(n120_adj_34), .CIN(mco_12_adj_6319), .COUT(mco_13_adj_6320), 
          .S0(mult_24s_7s_0_pp_1_7_adj_6101), .S1(mult_24s_7s_0_pp_1_8_adj_6100)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1024[11] 1026[50])
    defparam mult_24s_7s_0_mult_2_2_adj_145.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_2_adj_145.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_2_adj_145.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_2_adj_145.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_3_adj_146 (.A0(n34777), .B0(n117_adj_38), 
          .C0(GND_net), .D0(n120_adj_34), .A1(GND_net), .B1(n117_adj_38), 
          .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_13_adj_6320), 
          .COUT(mco_14_adj_6321), .S0(mult_24s_7s_0_pp_1_9_adj_6108), .S1(mult_24s_7s_0_pp_1_10_adj_6107)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1032[11] 1034[51])
    defparam mult_24s_7s_0_mult_2_3_adj_146.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_3_adj_146.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_3_adj_146.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_3_adj_146.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_4_adj_147 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_14_adj_6321), 
          .COUT(mco_15_adj_6322), .S0(mult_24s_7s_0_pp_1_11_adj_6115), .S1(mult_24s_7s_0_pp_1_12_adj_6114)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1040[11] 1042[51])
    defparam mult_24s_7s_0_mult_2_4_adj_147.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_4_adj_147.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_4_adj_147.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_4_adj_147.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_5_adj_148 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_15_adj_6322), 
          .COUT(mco_16_adj_6323), .S0(mult_24s_7s_0_pp_1_13_adj_6122), .S1(mult_24s_7s_0_pp_1_14_adj_6121)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1048[11] 1050[51])
    defparam mult_24s_7s_0_mult_2_5_adj_148.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_5_adj_148.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_5_adj_148.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_5_adj_148.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_6_adj_149 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_16_adj_6323), 
          .COUT(mco_17_adj_6324), .S0(mult_24s_7s_0_pp_1_15_adj_6129), .S1(mult_24s_7s_0_pp_1_16_adj_6128)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1056[11] 1058[51])
    defparam mult_24s_7s_0_mult_2_6_adj_149.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_6_adj_149.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_6_adj_149.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_6_adj_149.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_7_adj_150 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_17_adj_6324), 
          .COUT(mco_18_adj_6325), .S0(mult_24s_7s_0_pp_1_17_adj_6136), .S1(mult_24s_7s_0_pp_1_18_adj_6135)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1064[11] 1066[51])
    defparam mult_24s_7s_0_mult_2_7_adj_150.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_7_adj_150.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_7_adj_150.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_7_adj_150.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_8_adj_151 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_18_adj_6325), 
          .COUT(mco_19_adj_6326), .S0(mult_24s_7s_0_pp_1_19_adj_6143), .S1(mult_24s_7s_0_pp_1_20_adj_6142)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1072[11] 1074[51])
    defparam mult_24s_7s_0_mult_2_8_adj_151.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_8_adj_151.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_8_adj_151.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_8_adj_151.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_9_adj_152 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_19_adj_6326), 
          .COUT(mco_20_adj_6327), .S0(mult_24s_7s_0_pp_1_21_adj_6150), .S1(mult_24s_7s_0_pp_1_22_adj_6149)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1080[11] 1082[51])
    defparam mult_24s_7s_0_mult_2_9_adj_152.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_9_adj_152.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_9_adj_152.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_9_adj_152.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_10_adj_153 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(\rom4_w_i[12] ), .D0(n120_adj_34), .A1(\rom4_w_i[12] ), 
          .B1(n117_adj_38), .C1(\rom4_w_i[12] ), .D1(n120_adj_34), .CIN(mco_20_adj_6327), 
          .COUT(mco_21_adj_6328), .S0(mult_24s_7s_0_pp_1_23_adj_6157), .S1(mult_24s_7s_0_pp_1_24_adj_6156)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1088[11] 1090[51])
    defparam mult_24s_7s_0_mult_2_10_adj_153.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_10_adj_153.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_10_adj_153.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_10_adj_153.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_2_11_adj_154 (.A0(\rom4_w_i[12] ), .B0(n117_adj_38), 
          .C0(mult_24s_7s_0_mult_2_11_n2_adj_6034), .D0(VCC_net), .A1(mult_24s_7s_0_mult_2_11_n1_adj_6042), 
          .B1(VCC_net), .C1(GND_net), .D1(n120_adj_34), .CIN(mco_21_adj_6328), 
          .COUT(mfco_1_adj_6074), .S0(mult_24s_7s_0_pp_1_25_adj_6162), .S1(mult_24s_7s_0_pp_1_26_adj_6161)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1096[11] 1099[51])
    defparam mult_24s_7s_0_mult_2_11_adj_154.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_11_adj_154.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_2_11_adj_154.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_2_11_adj_154.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_0_adj_155 (.A0(n34777), .B0(n111_adj_39), 
          .C0(n34777), .D0(n114_adj_33), .A1(n34777), .B1(n111_adj_39), 
          .C1(GND_net), .D1(n114_adj_33), .CIN(mult_24s_7s_0_cin_lr_4_adj_6075), 
          .COUT(mco_22_adj_6329), .S0(mult_24s_7s_0_pp_2_5_adj_6232), .S1(mult_24s_7s_0_pp_2_6_adj_6169)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1105[11] 1107[77])
    defparam mult_24s_7s_0_mult_4_0_adj_155.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_0_adj_155.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_0_adj_155.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_0_adj_155.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_1_adj_156 (.A0(GND_net), .B0(n111_adj_39), 
          .C0(n34777), .D0(n114_adj_33), .A1(n34777), .B1(n111_adj_39), 
          .C1(GND_net), .D1(n114_adj_33), .CIN(mco_22_adj_6329), .COUT(mco_23_adj_6330), 
          .S0(mult_24s_7s_0_pp_2_7_adj_6174), .S1(mult_24s_7s_0_pp_2_8_adj_6173)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1113[11] 1115[50])
    defparam mult_24s_7s_0_mult_4_1_adj_156.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_1_adj_156.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_1_adj_156.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_1_adj_156.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_2_adj_157 (.A0(GND_net), .B0(n111_adj_39), 
          .C0(GND_net), .D0(n114_adj_33), .A1(GND_net), .B1(n111_adj_39), 
          .C1(n34777), .D1(n114_adj_33), .CIN(mco_23_adj_6330), .COUT(mco_24_adj_6331), 
          .S0(mult_24s_7s_0_pp_2_9_adj_6179), .S1(mult_24s_7s_0_pp_2_10_adj_6178)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1121[11] 1123[51])
    defparam mult_24s_7s_0_mult_4_2_adj_157.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_2_adj_157.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_2_adj_157.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_2_adj_157.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_3_adj_158 (.A0(n34777), .B0(n111_adj_39), 
          .C0(GND_net), .D0(n114_adj_33), .A1(GND_net), .B1(n111_adj_39), 
          .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_24_adj_6331), 
          .COUT(mco_25_adj_6332), .S0(mult_24s_7s_0_pp_2_11_adj_6184), .S1(mult_24s_7s_0_pp_2_12_adj_6183)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1129[11] 1131[51])
    defparam mult_24s_7s_0_mult_4_3_adj_158.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_3_adj_158.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_3_adj_158.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_3_adj_158.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_4_adj_159 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_25_adj_6332), 
          .COUT(mco_26_adj_6333), .S0(mult_24s_7s_0_pp_2_13_adj_6189), .S1(mult_24s_7s_0_pp_2_14_adj_6188)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1137[11] 1139[51])
    defparam mult_24s_7s_0_mult_4_4_adj_159.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_4_adj_159.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_4_adj_159.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_4_adj_159.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_5_adj_160 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_26_adj_6333), 
          .COUT(mco_27_adj_6334), .S0(mult_24s_7s_0_pp_2_15_adj_6194), .S1(mult_24s_7s_0_pp_2_16_adj_6193)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1145[11] 1147[51])
    defparam mult_24s_7s_0_mult_4_5_adj_160.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_5_adj_160.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_5_adj_160.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_5_adj_160.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_6_adj_161 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_27_adj_6334), 
          .COUT(mco_28_adj_6335), .S0(mult_24s_7s_0_pp_2_17_adj_6199), .S1(mult_24s_7s_0_pp_2_18_adj_6198)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1153[11] 1155[51])
    defparam mult_24s_7s_0_mult_4_6_adj_161.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_6_adj_161.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_6_adj_161.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_6_adj_161.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_7_adj_162 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_28_adj_6335), 
          .COUT(mco_29_adj_6336), .S0(mult_24s_7s_0_pp_2_19_adj_6204), .S1(mult_24s_7s_0_pp_2_20_adj_6203)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1161[11] 1163[51])
    defparam mult_24s_7s_0_mult_4_7_adj_162.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_7_adj_162.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_7_adj_162.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_7_adj_162.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_8_adj_163 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_29_adj_6336), 
          .COUT(mco_30_adj_6337), .S0(mult_24s_7s_0_pp_2_21_adj_6209), .S1(mult_24s_7s_0_pp_2_22_adj_6208)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1169[11] 1171[51])
    defparam mult_24s_7s_0_mult_4_8_adj_163.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_8_adj_163.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_8_adj_163.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_8_adj_163.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_9_adj_164 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_30_adj_6337), 
          .COUT(mco_31_adj_6338), .S0(mult_24s_7s_0_pp_2_23_adj_6214), .S1(mult_24s_7s_0_pp_2_24_adj_6213)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1177[11] 1179[51])
    defparam mult_24s_7s_0_mult_4_9_adj_164.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_9_adj_164.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_9_adj_164.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_9_adj_164.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_10_adj_165 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(\rom4_w_i[12] ), .D0(n114_adj_33), .A1(\rom4_w_i[12] ), 
          .B1(n111_adj_39), .C1(\rom4_w_i[12] ), .D1(n114_adj_33), .CIN(mco_31_adj_6338), 
          .COUT(mco_32_adj_6339), .S0(mult_24s_7s_0_pp_2_25_adj_6219), .S1(mult_24s_7s_0_pp_2_26_adj_6218)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1185[11] 1187[51])
    defparam mult_24s_7s_0_mult_4_10_adj_165.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_10_adj_165.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_10_adj_165.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_10_adj_165.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_mult_4_11_adj_166 (.A0(\rom4_w_i[12] ), .B0(n111_adj_39), 
          .C0(mult_24s_7s_0_mult_4_11_n2_adj_6032), .D0(VCC_net), .A1(mult_24s_7s_0_mult_4_11_n1_adj_6045), 
          .B1(VCC_net), .C1(GND_net), .D1(n114_adj_33), .CIN(mco_32_adj_6339), 
          .COUT(mfco_2_adj_6077), .S0(mult_24s_7s_0_pp_2_27_adj_6224), .S1(mult_24s_7s_0_pp_2_28_adj_6223)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(1197[11] 1200[51])
    defparam mult_24s_7s_0_mult_4_11_adj_166.INIT0 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_11_adj_166.INIT1 = 16'b0111100010001000;
    defparam mult_24s_7s_0_mult_4_11_adj_166.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_mult_4_11_adj_166.INJECT1_1 = "NO";
    CCU2C mult_24s_7s_0_cin_lr_add_0_adj_167 (.A0(VCC_net), .B0(VCC_net), 
          .C0(VCC_net), .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(mult_24s_7s_0_cin_lr_0_adj_6306)) /* synthesis syn_instantiated=1 */ ;   // mult_24s_7s.v(367[11] 369[77])
    defparam mult_24s_7s_0_cin_lr_add_0_adj_167.INIT0 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_0_adj_167.INIT1 = 16'b0000000000000000;
    defparam mult_24s_7s_0_cin_lr_add_0_adj_167.INJECT1_0 = "NO";
    defparam mult_24s_7s_0_cin_lr_add_0_adj_167.INJECT1_1 = "NO";
    LUT4 i20_3_lut_4_lut_adj_168 (.A(\op_r_23__N_1106[19] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[19] ), .Z(\dout_r_23__N_5681[19] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_168.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_169 (.A(\op_r_23__N_1106[11] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[11] ), .Z(\dout_r_23__N_5681[11] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_169.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_170 (.A(\op_r_23__N_1106[10] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[10] ), .Z(\dout_r_23__N_5681[10] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_170.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_171 (.A(\op_i_23__N_1154[9] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[9] ), .Z(\dout_i_23__N_5777[9] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_171.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_172 (.A(\op_r_23__N_1106[18] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[18] ), .Z(\dout_r_23__N_5681[18] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_172.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_173 (.A(\op_i_23__N_1154[8] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[8] ), .Z(\dout_i_23__N_5777[8] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_173.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_174 (.A(\op_r_23__N_1106[9] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[9] ), .Z(\dout_r_23__N_5681[9] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_174.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_175 (.A(\op_r_23__N_1106[8] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[8] ), .Z(\dout_r_23__N_5681[8] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_175.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_176 (.A(\op_i_23__N_1154[7] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[7] ), .Z(\dout_i_23__N_5777[7] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_176.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_177 (.A(\op_i_23__N_1154[6] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[6] ), .Z(\dout_i_23__N_5777[6] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_177.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_178 (.A(\op_i_23__N_1154[17] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[17] ), .Z(\dout_i_23__N_5777[17] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_178.init = 16'h8f80;
    LUT4 i10783_3_lut_4_lut (.A(\op_i_23__N_1154[23] ), .B(n34841), .C(n30179), 
         .D(\delay_i_23__N_1202[23] ), .Z(\dout_i_23__N_5777[23] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i10783_3_lut_4_lut.init = 16'h8f80;
    LUT4 i10736_3_lut_4_lut (.A(\op_r_23__N_1106[23] ), .B(n34841), .C(n30179), 
         .D(\delay_r_23__N_1178[23] ), .Z(\dout_r_23__N_5681[23] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i10736_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_179 (.A(\op_r_23__N_1106[22] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[22] ), .Z(\dout_r_23__N_5681[22] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_179.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_180 (.A(\op_i_23__N_1154[21] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[21] ), .Z(\dout_i_23__N_5777[21] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_180.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_181 (.A(\op_i_23__N_1154[16] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[16] ), .Z(\dout_i_23__N_5777[16] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_181.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_182 (.A(\op_i_23__N_1154[20] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[20] ), .Z(\dout_i_23__N_5777[20] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_182.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_183 (.A(\op_i_23__N_1154[5] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[5] ), .Z(\dout_i_23__N_5777[5] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_183.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_184 (.A(\op_i_23__N_1154[4] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[4] ), .Z(\dout_i_23__N_5777[4] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_184.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_185 (.A(\op_i_23__N_1154[3] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[3] ), .Z(\dout_i_23__N_5777[3] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_185.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_186 (.A(\op_i_23__N_1154[22] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[22] ), .Z(\dout_i_23__N_5777[22] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_186.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_187 (.A(\op_r_23__N_1106[7] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[7] ), .Z(\dout_r_23__N_5681[7] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_187.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_188 (.A(\op_r_23__N_1106[6] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[6] ), .Z(\dout_r_23__N_5681[6] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_188.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_189 (.A(\op_r_23__N_1106[5] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[5] ), .Z(\dout_r_23__N_5681[5] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_189.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_190 (.A(\op_r_23__N_1106[4] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[4] ), .Z(\dout_r_23__N_5681[4] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_190.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_191 (.A(\op_r_23__N_1106[17] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[17] ), .Z(\dout_r_23__N_5681[17] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_191.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_192 (.A(\op_r_23__N_1106[3] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[3] ), .Z(\dout_r_23__N_5681[3] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_192.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_193 (.A(\op_r_23__N_1106[2] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[2] ), .Z(\dout_r_23__N_5681[2] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_193.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_194 (.A(\op_r_23__N_1106[16] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[16] ), .Z(\dout_r_23__N_5681[16] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_194.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_195 (.A(\op_r_23__N_1106[1] ), .B(n34841), 
         .C(n30179), .D(\delay_r_23__N_1178[1] ), .Z(\dout_r_23__N_5681[1] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_195.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_196 (.A(\op_i_23__N_1154[15] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[15] ), .Z(\dout_i_23__N_5777[15] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_196.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut_adj_197 (.A(\op_i_23__N_1154[14] ), .B(n34841), 
         .C(n30179), .D(\delay_i_23__N_1202[14] ), .Z(\dout_i_23__N_5777[14] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i20_3_lut_4_lut_adj_197.init = 16'h8f80;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module shift_8
//

module shift_8 (clk_c, clk_c_enable_1419, \dout_i_23__N_4670[0] , \dout_r_23__N_4286[0] , 
            valid, clk_c_enable_2310, VCC_net, \dout_i_23__N_4670[1] , 
            \dout_i_23__N_4670[2] , \dout_i_23__N_4670[3] , \dout_i_23__N_4670[4] , 
            \dout_i_23__N_4670[5] , \dout_i_23__N_4670[6] , \dout_i_23__N_4670[7] , 
            \dout_i_23__N_4670[8] , \dout_i_23__N_4670[9] , \dout_i_23__N_4670[10] , 
            \dout_i_23__N_4670[11] , \dout_i_23__N_4670[12] , \dout_i_23__N_4670[13] , 
            \dout_i_23__N_4670[14] , \dout_i_23__N_4670[15] , \dout_i_23__N_4670[16] , 
            \dout_i_23__N_4670[17] , \dout_i_23__N_4670[18] , \dout_i_23__N_4670[19] , 
            \dout_i_23__N_4670[20] , \dout_i_23__N_4670[21] , \dout_i_23__N_4670[22] , 
            \dout_i_23__N_4670[23] , \dout_r_23__N_4286[1] , \dout_r_23__N_4286[2] , 
            \dout_r_23__N_4286[3] , \dout_r_23__N_4286[4] , \dout_r_23__N_4286[5] , 
            \dout_r_23__N_4286[6] , \dout_r_23__N_4286[7] , \dout_r_23__N_4286[8] , 
            \dout_r_23__N_4286[9] , \dout_r_23__N_4286[10] , \dout_r_23__N_4286[11] , 
            \dout_r_23__N_4286[12] , \dout_r_23__N_4286[13] , \dout_r_23__N_4286[14] , 
            \dout_r_23__N_4286[15] , \dout_r_23__N_4286[16] , \dout_r_23__N_4286[17] , 
            \dout_r_23__N_4286[18] , \dout_r_23__N_4286[19] , \dout_r_23__N_4286[20] , 
            \dout_r_23__N_4286[21] , \dout_r_23__N_4286[22] , \dout_r_23__N_4286[23] , 
            shift_8_dout_i, shift_8_dout_r) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input clk_c_enable_1419;
    input \dout_i_23__N_4670[0] ;
    input \dout_r_23__N_4286[0] ;
    output valid;
    input clk_c_enable_2310;
    input VCC_net;
    input \dout_i_23__N_4670[1] ;
    input \dout_i_23__N_4670[2] ;
    input \dout_i_23__N_4670[3] ;
    input \dout_i_23__N_4670[4] ;
    input \dout_i_23__N_4670[5] ;
    input \dout_i_23__N_4670[6] ;
    input \dout_i_23__N_4670[7] ;
    input \dout_i_23__N_4670[8] ;
    input \dout_i_23__N_4670[9] ;
    input \dout_i_23__N_4670[10] ;
    input \dout_i_23__N_4670[11] ;
    input \dout_i_23__N_4670[12] ;
    input \dout_i_23__N_4670[13] ;
    input \dout_i_23__N_4670[14] ;
    input \dout_i_23__N_4670[15] ;
    input \dout_i_23__N_4670[16] ;
    input \dout_i_23__N_4670[17] ;
    input \dout_i_23__N_4670[18] ;
    input \dout_i_23__N_4670[19] ;
    input \dout_i_23__N_4670[20] ;
    input \dout_i_23__N_4670[21] ;
    input \dout_i_23__N_4670[22] ;
    input \dout_i_23__N_4670[23] ;
    input \dout_r_23__N_4286[1] ;
    input \dout_r_23__N_4286[2] ;
    input \dout_r_23__N_4286[3] ;
    input \dout_r_23__N_4286[4] ;
    input \dout_r_23__N_4286[5] ;
    input \dout_r_23__N_4286[6] ;
    input \dout_r_23__N_4286[7] ;
    input \dout_r_23__N_4286[8] ;
    input \dout_r_23__N_4286[9] ;
    input \dout_r_23__N_4286[10] ;
    input \dout_r_23__N_4286[11] ;
    input \dout_r_23__N_4286[12] ;
    input \dout_r_23__N_4286[13] ;
    input \dout_r_23__N_4286[14] ;
    input \dout_r_23__N_4286[15] ;
    input \dout_r_23__N_4286[16] ;
    input \dout_r_23__N_4286[17] ;
    input \dout_r_23__N_4286[18] ;
    input \dout_r_23__N_4286[19] ;
    input \dout_r_23__N_4286[20] ;
    input \dout_r_23__N_4286[21] ;
    input \dout_r_23__N_4286[22] ;
    input \dout_r_23__N_4286[23] ;
    output [23:0]shift_8_dout_i;
    output [23:0]shift_8_dout_r;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    wire [191:0]dout_i_23__N_4670;
    wire [191:0]dout_r_23__N_4286;
    
    wire n29967, n29968, n29969, n29970, n29971, n29972, n29973, 
        n29974, n29975, n29976, n29977, n29978, n29979, n29980, 
        n29981, n29982, n29983, n29984, n29985, n29986, n29987, 
        n29988, n29989, n29990, n29991, n29992, n29993, n29994, 
        n29995, n29996, n29997, n29998, n29999, n30000, n30001, 
        n30002, n30003, n30004, n30005, n30006, n30007, n30008, 
        n30009, n30010, n30011, n30012, n30013, n30014;
    
    FD1P3AX shift_reg_i__i1 (.D(dout_i_23__N_4670[24]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i1.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i1 (.D(\dout_i_23__N_4670[0] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[24]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i1.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i1 (.D(dout_r_23__N_4286[24]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i1.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i1 (.D(\dout_r_23__N_4286[0] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[24]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i1.GSR = "ENABLED";
    FD1P3AX valid_26 (.D(VCC_net), .SP(clk_c_enable_2310), .CK(clk_c), 
            .Q(valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam valid_26.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i2 (.D(dout_i_23__N_4670[25]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i3 (.D(dout_i_23__N_4670[26]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i4 (.D(dout_i_23__N_4670[27]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i5 (.D(dout_i_23__N_4670[28]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i6 (.D(dout_i_23__N_4670[29]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i7 (.D(dout_i_23__N_4670[30]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i8 (.D(dout_i_23__N_4670[31]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i9 (.D(dout_i_23__N_4670[32]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i10 (.D(dout_i_23__N_4670[33]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i11 (.D(dout_i_23__N_4670[34]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i12 (.D(dout_i_23__N_4670[35]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i13 (.D(dout_i_23__N_4670[36]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i14 (.D(dout_i_23__N_4670[37]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i15 (.D(dout_i_23__N_4670[38]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i16 (.D(dout_i_23__N_4670[39]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i17 (.D(dout_i_23__N_4670[40]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i18 (.D(dout_i_23__N_4670[41]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i19 (.D(dout_i_23__N_4670[42]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i20 (.D(dout_i_23__N_4670[43]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i21 (.D(dout_i_23__N_4670[44]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i22 (.D(dout_i_23__N_4670[45]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i23 (.D(dout_i_23__N_4670[46]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i24 (.D(dout_i_23__N_4670[47]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i24.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i25 (.D(dout_i_23__N_4670[48]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i25.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i26 (.D(dout_i_23__N_4670[49]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i26.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i27 (.D(dout_i_23__N_4670[50]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i27.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i28 (.D(dout_i_23__N_4670[51]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i28.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i29 (.D(dout_i_23__N_4670[52]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i29.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i30 (.D(dout_i_23__N_4670[53]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[77])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i30.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i31 (.D(dout_i_23__N_4670[54]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[78])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i31.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i32 (.D(dout_i_23__N_4670[55]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[79])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i32.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i33 (.D(dout_i_23__N_4670[56]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i33.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i34 (.D(dout_i_23__N_4670[57]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i34.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i35 (.D(dout_i_23__N_4670[58]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i35.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i36 (.D(dout_i_23__N_4670[59]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i36.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i37 (.D(dout_i_23__N_4670[60]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i37.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i38 (.D(dout_i_23__N_4670[61]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[85])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i38.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i39 (.D(dout_i_23__N_4670[62]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[86])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i39.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i40 (.D(dout_i_23__N_4670[63]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[87])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i40.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i41 (.D(dout_i_23__N_4670[64]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i41.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i42 (.D(dout_i_23__N_4670[65]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i42.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i43 (.D(dout_i_23__N_4670[66]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i43.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i44 (.D(dout_i_23__N_4670[67]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i44.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i45 (.D(dout_i_23__N_4670[68]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i45.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i46 (.D(dout_i_23__N_4670[69]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[93])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i46.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i47 (.D(dout_i_23__N_4670[70]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[94])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i47.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i48 (.D(dout_i_23__N_4670[71]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[95])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i48.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i49 (.D(dout_i_23__N_4670[72]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[96])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i49.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i50 (.D(dout_i_23__N_4670[73]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[97])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i50.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i51 (.D(dout_i_23__N_4670[74]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[98])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i51.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i52 (.D(dout_i_23__N_4670[75]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[99])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i52.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i53 (.D(dout_i_23__N_4670[76]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[100])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i53.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i54 (.D(dout_i_23__N_4670[77]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[101])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i54.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i55 (.D(dout_i_23__N_4670[78]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[102])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i55.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i56 (.D(dout_i_23__N_4670[79]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[103])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i56.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i57 (.D(dout_i_23__N_4670[80]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[104])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i57.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i58 (.D(dout_i_23__N_4670[81]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[105])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i58.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i59 (.D(dout_i_23__N_4670[82]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[106])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i59.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i60 (.D(dout_i_23__N_4670[83]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[107])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i60.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i61 (.D(dout_i_23__N_4670[84]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[108])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i61.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i62 (.D(dout_i_23__N_4670[85]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[109])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i62.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i63 (.D(dout_i_23__N_4670[86]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[110])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i63.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i64 (.D(dout_i_23__N_4670[87]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[111])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i64.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i65 (.D(dout_i_23__N_4670[88]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[112])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i65.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i66 (.D(dout_i_23__N_4670[89]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[113])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i66.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i67 (.D(dout_i_23__N_4670[90]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[114])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i67.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i68 (.D(dout_i_23__N_4670[91]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[115])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i68.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i69 (.D(dout_i_23__N_4670[92]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[116])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i69.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i70 (.D(dout_i_23__N_4670[93]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[117])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i70.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i71 (.D(dout_i_23__N_4670[94]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[118])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i71.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i72 (.D(dout_i_23__N_4670[95]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[119])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i72.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i73 (.D(dout_i_23__N_4670[96]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[120])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i73.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i74 (.D(dout_i_23__N_4670[97]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[121])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i74.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i75 (.D(dout_i_23__N_4670[98]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[122])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i75.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i76 (.D(dout_i_23__N_4670[99]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[123])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i76.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i77 (.D(dout_i_23__N_4670[100]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[124])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i77.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i78 (.D(dout_i_23__N_4670[101]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[125])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i78.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i79 (.D(dout_i_23__N_4670[102]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[126])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i79.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i80 (.D(dout_i_23__N_4670[103]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[127])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i80.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i81 (.D(dout_i_23__N_4670[104]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[128])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i81.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i82 (.D(dout_i_23__N_4670[105]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[129])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i82.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i83 (.D(dout_i_23__N_4670[106]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[130])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i83.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i84 (.D(dout_i_23__N_4670[107]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[131])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i84.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i85 (.D(dout_i_23__N_4670[108]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[132])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i85.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i86 (.D(dout_i_23__N_4670[109]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[133])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i86.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i87 (.D(dout_i_23__N_4670[110]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[134])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i87.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i88 (.D(dout_i_23__N_4670[111]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[135])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i88.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i89 (.D(dout_i_23__N_4670[112]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[136])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i89.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i90 (.D(dout_i_23__N_4670[113]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[137])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i90.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i91 (.D(dout_i_23__N_4670[114]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[138])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i91.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i92 (.D(dout_i_23__N_4670[115]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[139])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i92.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i93 (.D(dout_i_23__N_4670[116]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[140])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i93.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i94 (.D(dout_i_23__N_4670[117]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[141])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i94.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i95 (.D(dout_i_23__N_4670[118]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[142])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i95.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i96 (.D(dout_i_23__N_4670[119]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[143])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i96.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i97 (.D(dout_i_23__N_4670[120]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[144])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i97.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i98 (.D(dout_i_23__N_4670[121]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[145])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i98.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i99 (.D(dout_i_23__N_4670[122]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[146])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i99.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i100 (.D(dout_i_23__N_4670[123]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[147])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i100.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i101 (.D(dout_i_23__N_4670[124]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[148])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i101.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i102 (.D(dout_i_23__N_4670[125]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[149])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i102.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i103 (.D(dout_i_23__N_4670[126]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[150])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i103.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i104 (.D(dout_i_23__N_4670[127]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[151])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i104.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i105 (.D(dout_i_23__N_4670[128]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[152])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i105.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i106 (.D(dout_i_23__N_4670[129]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[153])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i106.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i107 (.D(dout_i_23__N_4670[130]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[154])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i107.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i108 (.D(dout_i_23__N_4670[131]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[155])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i108.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i109 (.D(dout_i_23__N_4670[132]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[156])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i109.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i110 (.D(dout_i_23__N_4670[133]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[157])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i110.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i111 (.D(dout_i_23__N_4670[134]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[158])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i111.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i112 (.D(dout_i_23__N_4670[135]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[159])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i112.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i113 (.D(dout_i_23__N_4670[136]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[160])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i113.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i114 (.D(dout_i_23__N_4670[137]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[161])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i114.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i115 (.D(dout_i_23__N_4670[138]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[162])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i115.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i116 (.D(dout_i_23__N_4670[139]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[163])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i116.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i117 (.D(dout_i_23__N_4670[140]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[164])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i117.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i118 (.D(dout_i_23__N_4670[141]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[165])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i118.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i119 (.D(dout_i_23__N_4670[142]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[166])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i119.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i120 (.D(dout_i_23__N_4670[143]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[167])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i120.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i121 (.D(dout_i_23__N_4670[144]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[168])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i121.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i122 (.D(dout_i_23__N_4670[145]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[169])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i122.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i123 (.D(dout_i_23__N_4670[146]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[170])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i123.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i124 (.D(dout_i_23__N_4670[147]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[171])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i124.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i125 (.D(dout_i_23__N_4670[148]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[172])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i125.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i126 (.D(dout_i_23__N_4670[149]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[173])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i126.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i127 (.D(dout_i_23__N_4670[150]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[174])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i127.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i128 (.D(dout_i_23__N_4670[151]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[175])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i128.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i129 (.D(dout_i_23__N_4670[152]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[176])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i129.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i130 (.D(dout_i_23__N_4670[153]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[177])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i130.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i131 (.D(dout_i_23__N_4670[154]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[178])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i131.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i132 (.D(dout_i_23__N_4670[155]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[179])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i132.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i133 (.D(dout_i_23__N_4670[156]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[180])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i133.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i134 (.D(dout_i_23__N_4670[157]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[181])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i134.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i135 (.D(dout_i_23__N_4670[158]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[182])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i135.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i136 (.D(dout_i_23__N_4670[159]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[183])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i136.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i137 (.D(dout_i_23__N_4670[160]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[184])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i137.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i138 (.D(dout_i_23__N_4670[161]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[185])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i138.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i139 (.D(dout_i_23__N_4670[162]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[186])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i139.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i140 (.D(dout_i_23__N_4670[163]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[187])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i140.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i141 (.D(dout_i_23__N_4670[164]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[188])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i141.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i142 (.D(dout_i_23__N_4670[165]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[189])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i142.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i143 (.D(dout_i_23__N_4670[166]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[190])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i143.GSR = "ENABLED";
    FD1P3AX shift_reg_i__i144 (.D(dout_i_23__N_4670[167]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[191])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i144.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i2 (.D(\dout_i_23__N_4670[1] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i3 (.D(\dout_i_23__N_4670[2] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[26]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i4 (.D(\dout_i_23__N_4670[3] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i5 (.D(\dout_i_23__N_4670[4] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[28]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i6 (.D(\dout_i_23__N_4670[5] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i7 (.D(\dout_i_23__N_4670[6] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[30]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i8 (.D(\dout_i_23__N_4670[7] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i9 (.D(\dout_i_23__N_4670[8] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[32]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i10 (.D(\dout_i_23__N_4670[9] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[33]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i11 (.D(\dout_i_23__N_4670[10] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[34]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i12 (.D(\dout_i_23__N_4670[11] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[35]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i13 (.D(\dout_i_23__N_4670[12] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[36]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i14 (.D(\dout_i_23__N_4670[13] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[37]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i15 (.D(\dout_i_23__N_4670[14] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[38]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i16 (.D(\dout_i_23__N_4670[15] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[39]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i17 (.D(\dout_i_23__N_4670[16] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[40]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i18 (.D(\dout_i_23__N_4670[17] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[41]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i19 (.D(\dout_i_23__N_4670[18] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[42]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i20 (.D(\dout_i_23__N_4670[19] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[43]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i21 (.D(\dout_i_23__N_4670[20] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[44]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i22 (.D(\dout_i_23__N_4670[21] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[45]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i23 (.D(\dout_i_23__N_4670[22] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[46]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_i_res4__i24 (.D(\dout_i_23__N_4670[23] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_i_23__N_4670[47]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i_res4__i24.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i2 (.D(dout_r_23__N_4286[25]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i3 (.D(dout_r_23__N_4286[26]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i4 (.D(dout_r_23__N_4286[27]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i5 (.D(dout_r_23__N_4286[28]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i6 (.D(dout_r_23__N_4286[29]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i7 (.D(dout_r_23__N_4286[30]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i8 (.D(dout_r_23__N_4286[31]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i9 (.D(dout_r_23__N_4286[32]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i10 (.D(dout_r_23__N_4286[33]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i11 (.D(dout_r_23__N_4286[34]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i12 (.D(dout_r_23__N_4286[35]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i13 (.D(dout_r_23__N_4286[36]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i14 (.D(dout_r_23__N_4286[37]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i15 (.D(dout_r_23__N_4286[38]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i16 (.D(dout_r_23__N_4286[39]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i17 (.D(dout_r_23__N_4286[40]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i18 (.D(dout_r_23__N_4286[41]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i19 (.D(dout_r_23__N_4286[42]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i20 (.D(dout_r_23__N_4286[43]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i21 (.D(dout_r_23__N_4286[44]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i22 (.D(dout_r_23__N_4286[45]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i23 (.D(dout_r_23__N_4286[46]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i24 (.D(dout_r_23__N_4286[47]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i24.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i25 (.D(dout_r_23__N_4286[48]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i25.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i26 (.D(dout_r_23__N_4286[49]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i26.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i27 (.D(dout_r_23__N_4286[50]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i27.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i28 (.D(dout_r_23__N_4286[51]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i28.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i29 (.D(dout_r_23__N_4286[52]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i29.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i30 (.D(dout_r_23__N_4286[53]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[77])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i30.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i31 (.D(dout_r_23__N_4286[54]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[78])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i31.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i32 (.D(dout_r_23__N_4286[55]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[79])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i32.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i33 (.D(dout_r_23__N_4286[56]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i33.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i34 (.D(dout_r_23__N_4286[57]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i34.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i35 (.D(dout_r_23__N_4286[58]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i35.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i36 (.D(dout_r_23__N_4286[59]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i36.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i37 (.D(dout_r_23__N_4286[60]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i37.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i38 (.D(dout_r_23__N_4286[61]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[85])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i38.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i39 (.D(dout_r_23__N_4286[62]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[86])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i39.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i40 (.D(dout_r_23__N_4286[63]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[87])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i40.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i41 (.D(dout_r_23__N_4286[64]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i41.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i42 (.D(dout_r_23__N_4286[65]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i42.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i43 (.D(dout_r_23__N_4286[66]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i43.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i44 (.D(dout_r_23__N_4286[67]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i44.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i45 (.D(dout_r_23__N_4286[68]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i45.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i46 (.D(dout_r_23__N_4286[69]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[93])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i46.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i47 (.D(dout_r_23__N_4286[70]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[94])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i47.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i48 (.D(dout_r_23__N_4286[71]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[95])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i48.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i49 (.D(dout_r_23__N_4286[72]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[96])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i49.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i50 (.D(dout_r_23__N_4286[73]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[97])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i50.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i51 (.D(dout_r_23__N_4286[74]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[98])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i51.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i52 (.D(dout_r_23__N_4286[75]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[99])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i52.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i53 (.D(dout_r_23__N_4286[76]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[100])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i53.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i54 (.D(dout_r_23__N_4286[77]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[101])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i54.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i55 (.D(dout_r_23__N_4286[78]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[102])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i55.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i56 (.D(dout_r_23__N_4286[79]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[103])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i56.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i57 (.D(dout_r_23__N_4286[80]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[104])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i57.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i58 (.D(dout_r_23__N_4286[81]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[105])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i58.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i59 (.D(dout_r_23__N_4286[82]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[106])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i59.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i60 (.D(dout_r_23__N_4286[83]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[107])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i60.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i61 (.D(dout_r_23__N_4286[84]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[108])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i61.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i62 (.D(dout_r_23__N_4286[85]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[109])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i62.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i63 (.D(dout_r_23__N_4286[86]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[110])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i63.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i64 (.D(dout_r_23__N_4286[87]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[111])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i64.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i65 (.D(dout_r_23__N_4286[88]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[112])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i65.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i66 (.D(dout_r_23__N_4286[89]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[113])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i66.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i67 (.D(dout_r_23__N_4286[90]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[114])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i67.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i68 (.D(dout_r_23__N_4286[91]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[115])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i68.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i69 (.D(dout_r_23__N_4286[92]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[116])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i69.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i70 (.D(dout_r_23__N_4286[93]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[117])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i70.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i71 (.D(dout_r_23__N_4286[94]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[118])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i71.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i72 (.D(dout_r_23__N_4286[95]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[119])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i72.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i73 (.D(dout_r_23__N_4286[96]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[120])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i73.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i74 (.D(dout_r_23__N_4286[97]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[121])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i74.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i75 (.D(dout_r_23__N_4286[98]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[122])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i75.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i76 (.D(dout_r_23__N_4286[99]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[123])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i76.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i77 (.D(dout_r_23__N_4286[100]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[124])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i77.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i78 (.D(dout_r_23__N_4286[101]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[125])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i78.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i79 (.D(dout_r_23__N_4286[102]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[126])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i79.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i80 (.D(dout_r_23__N_4286[103]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[127])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i80.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i81 (.D(dout_r_23__N_4286[104]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[128])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i81.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i82 (.D(dout_r_23__N_4286[105]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[129])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i82.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i83 (.D(dout_r_23__N_4286[106]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[130])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i83.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i84 (.D(dout_r_23__N_4286[107]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[131])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i84.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i85 (.D(dout_r_23__N_4286[108]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[132])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i85.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i86 (.D(dout_r_23__N_4286[109]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[133])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i86.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i87 (.D(dout_r_23__N_4286[110]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[134])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i87.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i88 (.D(dout_r_23__N_4286[111]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[135])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i88.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i89 (.D(dout_r_23__N_4286[112]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[136])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i89.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i90 (.D(dout_r_23__N_4286[113]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[137])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i90.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i91 (.D(dout_r_23__N_4286[114]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[138])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i91.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i92 (.D(dout_r_23__N_4286[115]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[139])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i92.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i93 (.D(dout_r_23__N_4286[116]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[140])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i93.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i94 (.D(dout_r_23__N_4286[117]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[141])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i94.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i95 (.D(dout_r_23__N_4286[118]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[142])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i95.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i96 (.D(dout_r_23__N_4286[119]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[143])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i96.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i97 (.D(dout_r_23__N_4286[120]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[144])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i97.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i98 (.D(dout_r_23__N_4286[121]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[145])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i98.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i99 (.D(dout_r_23__N_4286[122]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[146])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i99.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i100 (.D(dout_r_23__N_4286[123]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[147])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i100.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i101 (.D(dout_r_23__N_4286[124]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[148])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i101.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i102 (.D(dout_r_23__N_4286[125]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[149])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i102.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i103 (.D(dout_r_23__N_4286[126]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[150])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i103.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i104 (.D(dout_r_23__N_4286[127]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[151])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i104.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i105 (.D(dout_r_23__N_4286[128]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[152])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i105.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i106 (.D(dout_r_23__N_4286[129]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[153])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i106.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i107 (.D(dout_r_23__N_4286[130]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[154])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i107.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i108 (.D(dout_r_23__N_4286[131]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[155])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i108.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i109 (.D(dout_r_23__N_4286[132]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[156])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i109.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i110 (.D(dout_r_23__N_4286[133]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[157])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i110.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i111 (.D(dout_r_23__N_4286[134]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[158])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i111.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i112 (.D(dout_r_23__N_4286[135]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[159])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i112.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i113 (.D(dout_r_23__N_4286[136]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[160])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i113.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i114 (.D(dout_r_23__N_4286[137]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[161])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i114.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i115 (.D(dout_r_23__N_4286[138]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[162])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i115.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i116 (.D(dout_r_23__N_4286[139]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[163])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i116.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i117 (.D(dout_r_23__N_4286[140]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[164])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i117.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i118 (.D(dout_r_23__N_4286[141]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[165])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i118.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i119 (.D(dout_r_23__N_4286[142]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[166])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i119.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i120 (.D(dout_r_23__N_4286[143]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[167])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i120.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i121 (.D(dout_r_23__N_4286[144]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[168])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i121.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i122 (.D(dout_r_23__N_4286[145]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[169])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i122.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i123 (.D(dout_r_23__N_4286[146]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[170])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i123.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i124 (.D(dout_r_23__N_4286[147]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[171])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i124.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i125 (.D(dout_r_23__N_4286[148]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[172])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i125.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i126 (.D(dout_r_23__N_4286[149]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[173])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i126.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i127 (.D(dout_r_23__N_4286[150]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[174])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i127.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i128 (.D(dout_r_23__N_4286[151]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[175])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i128.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i129 (.D(dout_r_23__N_4286[152]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[176])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i129.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i130 (.D(dout_r_23__N_4286[153]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[177])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i130.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i131 (.D(dout_r_23__N_4286[154]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[178])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i131.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i132 (.D(dout_r_23__N_4286[155]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[179])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i132.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i133 (.D(dout_r_23__N_4286[156]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[180])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i133.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i134 (.D(dout_r_23__N_4286[157]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[181])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i134.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i135 (.D(dout_r_23__N_4286[158]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[182])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i135.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i136 (.D(dout_r_23__N_4286[159]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[183])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i136.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i137 (.D(dout_r_23__N_4286[160]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[184])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i137.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i138 (.D(dout_r_23__N_4286[161]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[185])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i138.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i139 (.D(dout_r_23__N_4286[162]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[186])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i139.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i140 (.D(dout_r_23__N_4286[163]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[187])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i140.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i141 (.D(dout_r_23__N_4286[164]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[188])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i141.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i142 (.D(dout_r_23__N_4286[165]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[189])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i142.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i143 (.D(dout_r_23__N_4286[166]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[190])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i143.GSR = "ENABLED";
    FD1P3AX shift_reg_r__i144 (.D(dout_r_23__N_4286[167]), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[191])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i144.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i2 (.D(\dout_r_23__N_4286[1] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[25]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i2.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i3 (.D(\dout_r_23__N_4286[2] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[26]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i3.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i4 (.D(\dout_r_23__N_4286[3] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[27]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i4.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i5 (.D(\dout_r_23__N_4286[4] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[28]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i5.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i6 (.D(\dout_r_23__N_4286[5] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[29]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i6.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i7 (.D(\dout_r_23__N_4286[6] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[30]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i7.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i8 (.D(\dout_r_23__N_4286[7] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[31]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i8.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i9 (.D(\dout_r_23__N_4286[8] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[32]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i9.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i10 (.D(\dout_r_23__N_4286[9] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[33]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i10.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i11 (.D(\dout_r_23__N_4286[10] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[34]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i11.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i12 (.D(\dout_r_23__N_4286[11] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[35]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i12.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i13 (.D(\dout_r_23__N_4286[12] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[36]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i13.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i14 (.D(\dout_r_23__N_4286[13] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[37]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i14.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i15 (.D(\dout_r_23__N_4286[14] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[38]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i15.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i16 (.D(\dout_r_23__N_4286[15] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[39]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i16.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i17 (.D(\dout_r_23__N_4286[16] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[40]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i17.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i18 (.D(\dout_r_23__N_4286[17] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[41]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i18.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i19 (.D(\dout_r_23__N_4286[18] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[42]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i19.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i20 (.D(\dout_r_23__N_4286[19] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[43]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i20.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i21 (.D(\dout_r_23__N_4286[20] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[44]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i21.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i22 (.D(\dout_r_23__N_4286[21] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[45]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i22.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i23 (.D(\dout_r_23__N_4286[22] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[46]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i23.GSR = "ENABLED";
    FD1P3AX shift_reg_r_res1__i24 (.D(\dout_r_23__N_4286[23] ), .SP(clk_c_enable_1419), 
            .CK(clk_c), .Q(dout_r_23__N_4286[47]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r_res1__i24.GSR = "ENABLED";
    LUT4 i12257_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[191]), 
         .D(shift_8_dout_i[23]), .Z(n29967)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12257_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12258_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[190]), 
         .D(shift_8_dout_i[22]), .Z(n29968)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12258_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12259_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[189]), 
         .D(shift_8_dout_i[21]), .Z(n29969)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12259_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12260_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[188]), 
         .D(shift_8_dout_i[20]), .Z(n29970)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12260_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12261_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[187]), 
         .D(shift_8_dout_i[19]), .Z(n29971)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12261_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12262_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[186]), 
         .D(shift_8_dout_i[18]), .Z(n29972)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12262_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12263_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[185]), 
         .D(shift_8_dout_i[17]), .Z(n29973)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12263_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12264_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[184]), 
         .D(shift_8_dout_i[16]), .Z(n29974)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12264_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12265_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[183]), 
         .D(shift_8_dout_i[15]), .Z(n29975)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12265_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12266_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[182]), 
         .D(shift_8_dout_i[14]), .Z(n29976)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12266_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12267_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[181]), 
         .D(shift_8_dout_i[13]), .Z(n29977)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12267_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12268_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[180]), 
         .D(shift_8_dout_i[12]), .Z(n29978)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12268_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12269_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[179]), 
         .D(shift_8_dout_i[11]), .Z(n29979)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12269_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12270_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[178]), 
         .D(shift_8_dout_i[10]), .Z(n29980)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12270_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12271_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[177]), 
         .D(shift_8_dout_i[9]), .Z(n29981)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12271_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12272_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[176]), 
         .D(shift_8_dout_i[8]), .Z(n29982)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12272_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12273_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[175]), 
         .D(shift_8_dout_i[7]), .Z(n29983)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12273_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12274_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[174]), 
         .D(shift_8_dout_i[6]), .Z(n29984)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12274_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12275_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[173]), 
         .D(shift_8_dout_i[5]), .Z(n29985)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12275_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12276_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[172]), 
         .D(shift_8_dout_i[4]), .Z(n29986)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12276_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12277_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[171]), 
         .D(shift_8_dout_i[3]), .Z(n29987)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12277_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12278_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[170]), 
         .D(shift_8_dout_i[2]), .Z(n29988)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12278_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12279_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[169]), 
         .D(shift_8_dout_i[1]), .Z(n29989)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12279_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12280_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_i_23__N_4670[168]), 
         .D(shift_8_dout_i[0]), .Z(n29990)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12280_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12281_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[191]), 
         .D(shift_8_dout_r[23]), .Z(n29991)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12281_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12282_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[190]), 
         .D(shift_8_dout_r[22]), .Z(n29992)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12282_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12283_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[189]), 
         .D(shift_8_dout_r[21]), .Z(n29993)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12283_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12284_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[188]), 
         .D(shift_8_dout_r[20]), .Z(n29994)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12284_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12285_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[187]), 
         .D(shift_8_dout_r[19]), .Z(n29995)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12285_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12286_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[186]), 
         .D(shift_8_dout_r[18]), .Z(n29996)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12286_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12287_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[185]), 
         .D(shift_8_dout_r[17]), .Z(n29997)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12287_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12288_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[184]), 
         .D(shift_8_dout_r[16]), .Z(n29998)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12288_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12289_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[183]), 
         .D(shift_8_dout_r[15]), .Z(n29999)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12289_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12290_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[182]), 
         .D(shift_8_dout_r[14]), .Z(n30000)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12290_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12291_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[181]), 
         .D(shift_8_dout_r[13]), .Z(n30001)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12291_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12292_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[180]), 
         .D(shift_8_dout_r[12]), .Z(n30002)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12292_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12293_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[179]), 
         .D(shift_8_dout_r[11]), .Z(n30003)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12293_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12294_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[178]), 
         .D(shift_8_dout_r[10]), .Z(n30004)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12294_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12295_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[177]), 
         .D(shift_8_dout_r[9]), .Z(n30005)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12295_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12296_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[176]), 
         .D(shift_8_dout_r[8]), .Z(n30006)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12296_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12297_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[175]), 
         .D(shift_8_dout_r[7]), .Z(n30007)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12297_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12298_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[174]), 
         .D(shift_8_dout_r[6]), .Z(n30008)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12298_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12299_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[173]), 
         .D(shift_8_dout_r[5]), .Z(n30009)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12299_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12300_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[172]), 
         .D(shift_8_dout_r[4]), .Z(n30010)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12300_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12301_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[171]), 
         .D(shift_8_dout_r[3]), .Z(n30011)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12301_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12302_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[170]), 
         .D(shift_8_dout_r[2]), .Z(n30012)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12302_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12303_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[169]), 
         .D(shift_8_dout_r[1]), .Z(n30013)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12303_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12304_3_lut_4_lut (.A(valid), .B(clk_c_enable_2310), .C(dout_r_23__N_4286[168]), 
         .D(shift_8_dout_r[0]), .Z(n30014)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(41[14] 46[8])
    defparam i12304_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX shift_reg_r__i145 (.D(n30014), .CK(clk_c), .Q(shift_8_dout_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i145.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i146 (.D(n30013), .CK(clk_c), .Q(shift_8_dout_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i146.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i147 (.D(n30012), .CK(clk_c), .Q(shift_8_dout_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i147.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i148 (.D(n30011), .CK(clk_c), .Q(shift_8_dout_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i148.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i149 (.D(n30010), .CK(clk_c), .Q(shift_8_dout_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i149.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i150 (.D(n30009), .CK(clk_c), .Q(shift_8_dout_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i150.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i151 (.D(n30008), .CK(clk_c), .Q(shift_8_dout_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i151.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i152 (.D(n30007), .CK(clk_c), .Q(shift_8_dout_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i152.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i153 (.D(n30006), .CK(clk_c), .Q(shift_8_dout_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i153.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i154 (.D(n30005), .CK(clk_c), .Q(shift_8_dout_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i154.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i155 (.D(n30004), .CK(clk_c), .Q(shift_8_dout_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i155.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i156 (.D(n30003), .CK(clk_c), .Q(shift_8_dout_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i156.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i157 (.D(n30002), .CK(clk_c), .Q(shift_8_dout_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i157.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i158 (.D(n30001), .CK(clk_c), .Q(shift_8_dout_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i158.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i159 (.D(n30000), .CK(clk_c), .Q(shift_8_dout_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i159.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i160 (.D(n29999), .CK(clk_c), .Q(shift_8_dout_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i160.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i161 (.D(n29998), .CK(clk_c), .Q(shift_8_dout_r[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i161.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i162 (.D(n29997), .CK(clk_c), .Q(shift_8_dout_r[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i162.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i163 (.D(n29996), .CK(clk_c), .Q(shift_8_dout_r[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i163.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i164 (.D(n29995), .CK(clk_c), .Q(shift_8_dout_r[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i164.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i165 (.D(n29994), .CK(clk_c), .Q(shift_8_dout_r[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i165.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i166 (.D(n29993), .CK(clk_c), .Q(shift_8_dout_r[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i166.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i167 (.D(n29992), .CK(clk_c), .Q(shift_8_dout_r[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i167.GSR = "ENABLED";
    FD1S3AX shift_reg_r__i168 (.D(n29991), .CK(clk_c), .Q(shift_8_dout_r[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_r__i168.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i145 (.D(n29990), .CK(clk_c), .Q(shift_8_dout_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i145.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i146 (.D(n29989), .CK(clk_c), .Q(shift_8_dout_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i146.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i147 (.D(n29988), .CK(clk_c), .Q(shift_8_dout_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i147.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i148 (.D(n29987), .CK(clk_c), .Q(shift_8_dout_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i148.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i149 (.D(n29986), .CK(clk_c), .Q(shift_8_dout_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i149.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i150 (.D(n29985), .CK(clk_c), .Q(shift_8_dout_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i150.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i151 (.D(n29984), .CK(clk_c), .Q(shift_8_dout_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i151.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i152 (.D(n29983), .CK(clk_c), .Q(shift_8_dout_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i152.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i153 (.D(n29982), .CK(clk_c), .Q(shift_8_dout_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i153.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i154 (.D(n29981), .CK(clk_c), .Q(shift_8_dout_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i154.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i155 (.D(n29980), .CK(clk_c), .Q(shift_8_dout_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i155.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i156 (.D(n29979), .CK(clk_c), .Q(shift_8_dout_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i156.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i157 (.D(n29978), .CK(clk_c), .Q(shift_8_dout_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i157.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i158 (.D(n29977), .CK(clk_c), .Q(shift_8_dout_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i158.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i159 (.D(n29976), .CK(clk_c), .Q(shift_8_dout_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i159.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i160 (.D(n29975), .CK(clk_c), .Q(shift_8_dout_i[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i160.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i161 (.D(n29974), .CK(clk_c), .Q(shift_8_dout_i[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i161.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i162 (.D(n29973), .CK(clk_c), .Q(shift_8_dout_i[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i162.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i163 (.D(n29972), .CK(clk_c), .Q(shift_8_dout_i[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i163.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i164 (.D(n29971), .CK(clk_c), .Q(shift_8_dout_i[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i164.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i165 (.D(n29970), .CK(clk_c), .Q(shift_8_dout_i[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i165.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i166 (.D(n29969), .CK(clk_c), .Q(shift_8_dout_i[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i166.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i167 (.D(n29968), .CK(clk_c), .Q(shift_8_dout_i[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i167.GSR = "ENABLED";
    FD1S3AX shift_reg_i__i168 (.D(n29967), .CK(clk_c), .Q(shift_8_dout_i[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=130, LSE_RLINE=137 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_8.v(36[5] 46[8])
    defparam shift_reg_i__i168.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module radix2
//

module radix2 (dout_i_23__N_5974, GND_net, VCC_net, clk_c, n34738, 
            rst_n_N_2, \op_r_23__N_1226[0] , \op_r_23__N_1226[1] , \op_r_23__N_1226[2] , 
            \op_r_23__N_1226[3] , \op_r_23__N_1226[4] , \op_r_23__N_1226[5] , 
            \op_r_23__N_1226[6] , \op_r_23__N_1226[7] , \op_r_23__N_1226[8] , 
            \op_r_23__N_1226[9] , \op_r_23__N_1226[10] , \op_r_23__N_1226[11] , 
            \op_r_23__N_1226[12] , \op_r_23__N_1226[13] , \op_r_23__N_1226[14] , 
            \op_r_23__N_1226[15] , \op_r_23__N_1226[16] , \op_r_23__N_1226[17] , 
            \op_r_23__N_1226[18] , \op_r_23__N_1226[19] , \op_r_23__N_1226[20] , 
            \op_r_23__N_1226[21] , \op_r_23__N_1226[22] , \op_r_23__N_1226[23] , 
            \op_r_23__N_1226[24] , \op_r_23__N_1226[25] , \op_r_23__N_1226[26] , 
            \op_r_23__N_1226[27] , \op_r_23__N_1226[28] , \op_r_23__N_1226[29] , 
            \op_r_23__N_1226[30] , \op_r_23__N_1226[31] , \op_i_23__N_1310[0] , 
            \op_i_23__N_1310[1] , \op_i_23__N_1310[2] , \op_i_23__N_1310[3] , 
            \op_i_23__N_1310[4] , \op_i_23__N_1310[5] , n89, n88, n87, 
            n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, 
            n76, n75, n74, n73, n72, n71, n70, n69, n68, n67, 
            n66, n65, n11556, n11557, n11558, n11559, n11560, 
            n11561, n12083, n12084, n12085, n12086, n12087, n12088, 
            n12089, n12065, n12066, n12067, n12068, n12069, n12070, 
            n12071, n12072, n12073, n12074, n12075, n12076, n12077, 
            n12078, n12079, n12080, n12081, n12082, \op_r_23__N_1268[0] , 
            \op_r_23__N_1268[1] , \op_r_23__N_1268[2] , \op_r_23__N_1268[3] , 
            \op_r_23__N_1268[4] , \op_r_23__N_1268[5] , \op_r_23__N_1268[6] , 
            \op_r_23__N_1268[7] , \op_r_23__N_1268[8] , \op_r_23__N_1268[9] , 
            \op_r_23__N_1268[10] , \op_r_23__N_1268[11] , \op_r_23__N_1268[12] , 
            \op_r_23__N_1268[13] , \op_r_23__N_1268[14] , \op_r_23__N_1268[15] , 
            \op_r_23__N_1268[16] , \op_r_23__N_1268[17] , \op_r_23__N_1268[18] , 
            \op_r_23__N_1268[19] , \op_r_23__N_1268[20] , \op_r_23__N_1268[21] , 
            \op_r_23__N_1268[22] , \op_r_23__N_1268[23] , \op_r_23__N_1268[24] , 
            \op_r_23__N_1268[25] , \op_r_23__N_1268[26] , \op_r_23__N_1268[27] , 
            \op_r_23__N_1268[28] , \op_r_23__N_1268[29] , \op_r_23__N_1268[30] , 
            \op_r_23__N_1268[31] , n9105, n9104, n9103, n9102, n9101, 
            n9100, n9099, n9098, n9097, n9096, n9095, n9094, n9093, 
            n9092, n9091, n9090, n9089, n9088, n9087, n9086, n9085, 
            n9084, n9083, n9082, n9081, n9080, n319, n11562, n11563, 
            n11564, n11565, n11566, n11567, n11568, n11569, n11570, 
            n11571, n11572, n11573, n11574, n11575, n11576, n11577, 
            n11578, n11579, n34843, delay_i_23__N_1202, \no5_state[0] , 
            op_i_23__N_1154, delay_r_23__N_1178, op_r_23__N_1106, dout_r_23__N_5926, 
            s5_count, r4_valid, \op_i_23__N_1130[16] , \op_i_23__N_1154[8]_adj_1 , 
            \out_i[8] , \op_i_23__N_1130[21] , \op_i_23__N_1154[13]_adj_2 , 
            \out_i[13] , \op_i_23__N_1130[20] , \op_i_23__N_1154[12]_adj_3 , 
            \out_i[12] , \op_i_23__N_1130[19] , \op_i_23__N_1154[11]_adj_4 , 
            \out_i[11] , \op_i_23__N_1130[18] , \op_i_23__N_1154[10]_adj_5 , 
            \out_i[10] , \op_i_23__N_1130[17] , \op_i_23__N_1154[9]_adj_6 , 
            \out_i[9] , \op_i_23__N_1130[31] , \op_i_23__N_1154[23]_adj_7 , 
            \out_i[23] , \op_i_23__N_1130[30] , \op_i_23__N_1154[22]_adj_8 , 
            \out_i[22] , \op_i_23__N_1130[29] , \op_i_23__N_1154[21]_adj_9 , 
            \out_i[21] , \op_i_23__N_1130[28] , \op_i_23__N_1154[20]_adj_10 , 
            \out_i[20] , \op_i_23__N_1130[27] , \op_i_23__N_1154[19]_adj_11 , 
            \out_i[19] , \op_i_23__N_1130[26] , \op_i_23__N_1154[18]_adj_12 , 
            \out_i[18] , \op_i_23__N_1130[25] , \op_i_23__N_1154[17]_adj_13 , 
            \out_i[17] , \op_i_23__N_1130[24] , \op_i_23__N_1154[16]_adj_14 , 
            \out_i[16] , \op_i_23__N_1130[23] , \op_i_23__N_1154[15]_adj_15 , 
            \out_i[15] , \op_i_23__N_1130[22] , \op_i_23__N_1154[14]_adj_16 , 
            \out_i[14] , \op_r_23__N_1082[16] , \op_r_23__N_1106[8]_adj_17 , 
            \out_r[8] , \op_r_23__N_1082[17] , \op_r_23__N_1106[9]_adj_18 , 
            \out_r[9] , \op_r_23__N_1082[18] , \op_r_23__N_1106[10]_adj_19 , 
            \out_r[10] , \op_r_23__N_1082[19] , \op_r_23__N_1106[11]_adj_20 , 
            \out_r[11] , \op_r_23__N_1082[20] , \op_r_23__N_1106[12]_adj_21 , 
            \out_r[12] , \op_r_23__N_1082[21] , \op_r_23__N_1106[13]_adj_22 , 
            \out_r[13] , \op_r_23__N_1082[22] , \op_r_23__N_1106[14]_adj_23 , 
            \out_r[14] , \op_r_23__N_1082[23] , \op_r_23__N_1106[15]_adj_24 , 
            \out_r[15] , \op_r_23__N_1082[24] , \op_r_23__N_1106[16]_adj_25 , 
            \out_r[16] , \op_r_23__N_1082[25] , \op_r_23__N_1106[17]_adj_26 , 
            \out_r[17] , \op_r_23__N_1082[26] , \op_r_23__N_1106[18]_adj_27 , 
            \out_r[18] , \op_r_23__N_1082[27] , \op_r_23__N_1106[19]_adj_28 , 
            \out_r[19] , \op_r_23__N_1082[28] , \op_r_23__N_1106[20]_adj_29 , 
            \out_r[20] , \op_r_23__N_1082[29] , \op_r_23__N_1106[21]_adj_30 , 
            \out_r[21] , \op_r_23__N_1082[30] , \op_r_23__N_1106[22]_adj_31 , 
            \out_r[22] , \op_r_23__N_1082[31] , \op_r_23__N_1106[23]_adj_32 , 
            \out_r[23] ) /* synthesis syn_module_defined=1 */ ;
    output [23:0]dout_i_23__N_5974;
    input GND_net;
    input VCC_net;
    input clk_c;
    input n34738;
    input rst_n_N_2;
    output \op_r_23__N_1226[0] ;
    output \op_r_23__N_1226[1] ;
    output \op_r_23__N_1226[2] ;
    output \op_r_23__N_1226[3] ;
    output \op_r_23__N_1226[4] ;
    output \op_r_23__N_1226[5] ;
    output \op_r_23__N_1226[6] ;
    output \op_r_23__N_1226[7] ;
    output \op_r_23__N_1226[8] ;
    output \op_r_23__N_1226[9] ;
    output \op_r_23__N_1226[10] ;
    output \op_r_23__N_1226[11] ;
    output \op_r_23__N_1226[12] ;
    output \op_r_23__N_1226[13] ;
    output \op_r_23__N_1226[14] ;
    output \op_r_23__N_1226[15] ;
    output \op_r_23__N_1226[16] ;
    output \op_r_23__N_1226[17] ;
    output \op_r_23__N_1226[18] ;
    output \op_r_23__N_1226[19] ;
    output \op_r_23__N_1226[20] ;
    output \op_r_23__N_1226[21] ;
    output \op_r_23__N_1226[22] ;
    output \op_r_23__N_1226[23] ;
    output \op_r_23__N_1226[24] ;
    output \op_r_23__N_1226[25] ;
    output \op_r_23__N_1226[26] ;
    output \op_r_23__N_1226[27] ;
    output \op_r_23__N_1226[28] ;
    output \op_r_23__N_1226[29] ;
    output \op_r_23__N_1226[30] ;
    output \op_r_23__N_1226[31] ;
    output \op_i_23__N_1310[0] ;
    output \op_i_23__N_1310[1] ;
    output \op_i_23__N_1310[2] ;
    output \op_i_23__N_1310[3] ;
    output \op_i_23__N_1310[4] ;
    output \op_i_23__N_1310[5] ;
    output n89;
    output n88;
    output n87;
    output n86;
    output n85;
    output n84;
    output n83;
    output n82;
    output n81;
    output n80;
    output n79;
    output n78;
    output n77;
    output n76;
    output n75;
    output n74;
    output n73;
    output n72;
    output n71;
    output n70;
    output n69;
    output n68;
    output n67;
    output n66;
    output n65;
    input n11556;
    input n11557;
    input n11558;
    input n11559;
    input n11560;
    input n11561;
    input n12083;
    input n12084;
    input n12085;
    input n12086;
    input n12087;
    input n12088;
    input n12089;
    input n12065;
    input n12066;
    input n12067;
    input n12068;
    input n12069;
    input n12070;
    input n12071;
    input n12072;
    input n12073;
    input n12074;
    input n12075;
    input n12076;
    input n12077;
    input n12078;
    input n12079;
    input n12080;
    input n12081;
    input n12082;
    output \op_r_23__N_1268[0] ;
    output \op_r_23__N_1268[1] ;
    output \op_r_23__N_1268[2] ;
    output \op_r_23__N_1268[3] ;
    output \op_r_23__N_1268[4] ;
    output \op_r_23__N_1268[5] ;
    output \op_r_23__N_1268[6] ;
    output \op_r_23__N_1268[7] ;
    output \op_r_23__N_1268[8] ;
    output \op_r_23__N_1268[9] ;
    output \op_r_23__N_1268[10] ;
    output \op_r_23__N_1268[11] ;
    output \op_r_23__N_1268[12] ;
    output \op_r_23__N_1268[13] ;
    output \op_r_23__N_1268[14] ;
    output \op_r_23__N_1268[15] ;
    output \op_r_23__N_1268[16] ;
    output \op_r_23__N_1268[17] ;
    output \op_r_23__N_1268[18] ;
    output \op_r_23__N_1268[19] ;
    output \op_r_23__N_1268[20] ;
    output \op_r_23__N_1268[21] ;
    output \op_r_23__N_1268[22] ;
    output \op_r_23__N_1268[23] ;
    output \op_r_23__N_1268[24] ;
    output \op_r_23__N_1268[25] ;
    output \op_r_23__N_1268[26] ;
    output \op_r_23__N_1268[27] ;
    output \op_r_23__N_1268[28] ;
    output \op_r_23__N_1268[29] ;
    output \op_r_23__N_1268[30] ;
    output \op_r_23__N_1268[31] ;
    output n9105;
    output n9104;
    output n9103;
    output n9102;
    output n9101;
    output n9100;
    output n9099;
    output n9098;
    output n9097;
    output n9096;
    output n9095;
    output n9094;
    output n9093;
    output n9092;
    output n9091;
    output n9090;
    output n9089;
    output n9088;
    output n9087;
    output n9086;
    output n9085;
    output n9084;
    output n9083;
    output n9082;
    output n9081;
    output n9080;
    input n319;
    input n11562;
    input n11563;
    input n11564;
    input n11565;
    input n11566;
    input n11567;
    input n11568;
    input n11569;
    input n11570;
    input n11571;
    input n11572;
    input n11573;
    input n11574;
    input n11575;
    input n11576;
    input n11577;
    input n11578;
    input n11579;
    input n34843;
    input [23:0]delay_i_23__N_1202;
    input \no5_state[0] ;
    input [23:0]op_i_23__N_1154;
    input [23:0]delay_r_23__N_1178;
    input [23:0]op_r_23__N_1106;
    output [23:0]dout_r_23__N_5926;
    input s5_count;
    input r4_valid;
    input \op_i_23__N_1130[16] ;
    input \op_i_23__N_1154[8]_adj_1 ;
    output \out_i[8] ;
    input \op_i_23__N_1130[21] ;
    input \op_i_23__N_1154[13]_adj_2 ;
    output \out_i[13] ;
    input \op_i_23__N_1130[20] ;
    input \op_i_23__N_1154[12]_adj_3 ;
    output \out_i[12] ;
    input \op_i_23__N_1130[19] ;
    input \op_i_23__N_1154[11]_adj_4 ;
    output \out_i[11] ;
    input \op_i_23__N_1130[18] ;
    input \op_i_23__N_1154[10]_adj_5 ;
    output \out_i[10] ;
    input \op_i_23__N_1130[17] ;
    input \op_i_23__N_1154[9]_adj_6 ;
    output \out_i[9] ;
    input \op_i_23__N_1130[31] ;
    input \op_i_23__N_1154[23]_adj_7 ;
    output \out_i[23] ;
    input \op_i_23__N_1130[30] ;
    input \op_i_23__N_1154[22]_adj_8 ;
    output \out_i[22] ;
    input \op_i_23__N_1130[29] ;
    input \op_i_23__N_1154[21]_adj_9 ;
    output \out_i[21] ;
    input \op_i_23__N_1130[28] ;
    input \op_i_23__N_1154[20]_adj_10 ;
    output \out_i[20] ;
    input \op_i_23__N_1130[27] ;
    input \op_i_23__N_1154[19]_adj_11 ;
    output \out_i[19] ;
    input \op_i_23__N_1130[26] ;
    input \op_i_23__N_1154[18]_adj_12 ;
    output \out_i[18] ;
    input \op_i_23__N_1130[25] ;
    input \op_i_23__N_1154[17]_adj_13 ;
    output \out_i[17] ;
    input \op_i_23__N_1130[24] ;
    input \op_i_23__N_1154[16]_adj_14 ;
    output \out_i[16] ;
    input \op_i_23__N_1130[23] ;
    input \op_i_23__N_1154[15]_adj_15 ;
    output \out_i[15] ;
    input \op_i_23__N_1130[22] ;
    input \op_i_23__N_1154[14]_adj_16 ;
    output \out_i[14] ;
    input \op_r_23__N_1082[16] ;
    input \op_r_23__N_1106[8]_adj_17 ;
    output \out_r[8] ;
    input \op_r_23__N_1082[17] ;
    input \op_r_23__N_1106[9]_adj_18 ;
    output \out_r[9] ;
    input \op_r_23__N_1082[18] ;
    input \op_r_23__N_1106[10]_adj_19 ;
    output \out_r[10] ;
    input \op_r_23__N_1082[19] ;
    input \op_r_23__N_1106[11]_adj_20 ;
    output \out_r[11] ;
    input \op_r_23__N_1082[20] ;
    input \op_r_23__N_1106[12]_adj_21 ;
    output \out_r[12] ;
    input \op_r_23__N_1082[21] ;
    input \op_r_23__N_1106[13]_adj_22 ;
    output \out_r[13] ;
    input \op_r_23__N_1082[22] ;
    input \op_r_23__N_1106[14]_adj_23 ;
    output \out_r[14] ;
    input \op_r_23__N_1082[23] ;
    input \op_r_23__N_1106[15]_adj_24 ;
    output \out_r[15] ;
    input \op_r_23__N_1082[24] ;
    input \op_r_23__N_1106[16]_adj_25 ;
    output \out_r[16] ;
    input \op_r_23__N_1082[25] ;
    input \op_r_23__N_1106[17]_adj_26 ;
    output \out_r[17] ;
    input \op_r_23__N_1082[26] ;
    input \op_r_23__N_1106[18]_adj_27 ;
    output \out_r[18] ;
    input \op_r_23__N_1082[27] ;
    input \op_r_23__N_1106[19]_adj_28 ;
    output \out_r[19] ;
    input \op_r_23__N_1082[28] ;
    input \op_r_23__N_1106[20]_adj_29 ;
    output \out_r[20] ;
    input \op_r_23__N_1082[29] ;
    input \op_r_23__N_1106[21]_adj_30 ;
    output \out_r[21] ;
    input \op_r_23__N_1082[30] ;
    input \op_r_23__N_1106[22]_adj_31 ;
    output \out_r[22] ;
    input \op_r_23__N_1082[31] ;
    input \op_r_23__N_1106[23]_adj_32 ;
    output \out_r[23] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire n16014, n16015, n16016, n16017, n16018, n16019, n16020, 
        n16021, n16022, n16023, n16024, n16025, n16026, n16027, 
        n16028, n16029, n16030, n16031, n16032, n16033, n16034, 
        n16035, n16036, n16037, n16038, n16039, n16040, n16041, 
        n16042, n16043, n16044, n16045, n16046, n16047, n16048, 
        n16049, n16050, n16051, n16052, n16053, n16054, n16055, 
        n16056, n16057, n16058, n16059, n16060, n16061, n16062, 
        n16063, n16064, n16065, n16066, n16067, n16068, n16069, 
        n16070, n16071, n16072, n16073, n16074, n16075, n16076, 
        n16077, n16078, n16079, n16080, n16081, n16082, n16083, 
        n16084, n16085, n16086, n15468, n15469, n15470, n15471, 
        n15472, n15473, n15474, n15475, n15476, n15477, n15478, 
        n15479, n15480, n15481, n15482, n15483, n15484, n15485, 
        n15486, n15487, n15488, n15489, n15490, n15491, n15492, 
        n15493, n15494, n15495, n15496, n15497, n15498, n15499, 
        n15500, n15501, n15502, n15503, n15504, n15505, n15506, 
        n15507, n15508, n15509, n15510, n15511, n15512, n15513, 
        n15514, n15515, n15516, n15517, n15518, n15519, n15520, 
        n15521, n15522, n15523, n15524, n15525, n15526, n15527, 
        n15528, n15529, n15530, n15531, n15532, n15533, n15534, 
        n15535, n15536, n15537, n15538, n15539, n15540, n15541, 
        n15542, n15543, n15544, n15545, n15546, n15547, n15548, 
        n15549, n15550, n15551, n15552, n15553, n15554, n15555, 
        n15556, n15557, n15558, n15559, n15560, n15561, n15562, 
        n15563, n15564, n15565, n15566, n15567, n15568, n15569, 
        n15570, n15571, n15572, n15573, n15574, n15575, n15576, 
        n15577, n15578, n15579, n15580, n15581, n15582, n15583, 
        n15584, n15585, n15586, n15587, n15588, n15589, n15590, 
        n15591, n15592, n15593, n15594, n15595, n15596, n15597, 
        n15598, n15599, n15600, n15601, n15602, n15603, n15604, 
        n15605, n15606, n15607, n15608, n15609, n15610, n15611, 
        n15612, n15613, n15614, n15615, n15616, n15617, n15618, 
        n15619, n15620, n15621, n15622, n15623, n15624, n15625, 
        n15626, n15627, n15628, n15629, n15630, n15631, n15632, 
        n15633, n15634, n15635, n15636, n15637, n15638, n15639, 
        n15640, n15641, n15642, n15643, n15644, n15645, n15646, 
        n15647, n15648, n15649, n15650, n18711, n18712, n18713, 
        n18714, n18715, n18716, n18717, n18718, n18719, n18720, 
        n18721, n18722, n18723, n18724, n18725, n18726, n18727, 
        n18728, n18729, n18730, n18731, n18732, n18733, n18734, 
        n18735, n18736, n18737, n18738, n18739, n18740, n18741, 
        n18742, n18743, n18744, n18745, n18746, n18747, n18748, 
        n18749, n18750, n18751, n18752, n18753, n18754, n18755, 
        n18756, n18757, n18758, n18759, n18760, n18761, n18762, 
        n18763, n18764, n18765, n18766, n18767, n18768, n18769, 
        n18770, n18771, n18772, n18773, n18774, n18775, n18776, 
        n18777, n18778, n18779, n18780, n18781, n18782, n18783, 
        n18784, n18785, n18786, n18787, n18788, n18789, n18790, 
        n18791, n18792, n18793, n18794, n18795, n18796, n18797, 
        n18798, n18799, n18800, n18801, n18802, n18803, n18804, 
        n18805, n18806, n18807, n18808, n18809, n18810, n18811, 
        n18812, n18813, n18814, n18815, n18816, n18817, n18818, 
        n18819, n18820, n18821, n18822, n18823, n18824, n18825, 
        n18826, n18827, n18828, n18829, n18830, n18831, n18832, 
        n18833, n18834, n18835, n18836, n18837, n18838, n18839, 
        n18840, n18841, n18842, n18843, n18844, n18845, n18846, 
        n18847, n18848, n18849, n18850, n18851, n18852, n18853, 
        n18854, n18855, n18856, n15322, n15323, n15324, n15325, 
        n15326, n15327, n15328, n15329, n15330, n15331, n15332, 
        n15333, n15334, n15335, n15336, n15337, n15338, n15339, 
        n15340, n15341, n15342, n15343, n15344, n15345, n15346, 
        n15347, n15348, n15349, n15350, n15351, n15352, n15353, 
        n15354, n15355, n15356, n15357, n15358, n15359, n15360, 
        n15361, n15362, n15363, n15364, n15365, n15366, n15367, 
        n15368, n15369, n15370, n15371, n15372, n15373, n15374, 
        n15375, n15376, n15377, n15378, n15379, n15380, n15381, 
        n15382, n15383, n15384, n15385, n15386, n15387, n15388, 
        n15389, n15390, n15391, n15392, n15393, n15394, n15395, 
        n15396, n15397, n15398, n15399, n15400, n15401, n15402, 
        n15403, n15404, n15405, n15406, n15407, n15408, n15409, 
        n15410, n15411, n15412, n15413, n15414, n15415, n15416, 
        n15417, n15418, n15419, n15420, n15421, n15422, n15423, 
        n15424, n15425, n15426, n15427, n15428, n15429, n15430, 
        n15431, n15432, n15433, n15434, n15435, n15436, n15437, 
        n15438, n15439, n15440, n15441, n15442, n15443, n15444, 
        n15445, n15446, n15447, n15448, n15449, n15450, n15451, 
        n15452, n15453, n15454, n15455, n15456, n15457, n15458, 
        n15459, n15460, n15461, n15462, n15463, n15464, n15465, 
        n15466, n15467, n16233, n16234, n16235, n16236, n16237, 
        n16238, n16239, n16240, n16241, n16242, n16243, n16244, 
        n16245, n16246, n16247, n16248, n16249, n16250, n16251, 
        n16252, n16253, n16254, n16255, n16256, n16257, n16258, 
        n16259, n16260, n16261, n16262, n16263, n16264, n16265, 
        n16266, n16267, n16268, n16269, n16270, n16271, n16272, 
        n16273, n16274, n16275, n16276, n16277, n16278, n16279, 
        n16280, n16281, n16282, n16283, n16284, n16285, n16286, 
        n16287, n16288, n16289, n16290, n16291, n16292, n16293, 
        n16294, n16295, n16296, n16297, n16298, n16299, n16300, 
        n16301, n16302, n16303, n16304, n16305, n16160, n16161, 
        n16162, n16163, n16164, n16165, n16166, n16167, n16168, 
        n16169, n16170, n16171, n16172, n16173, n16174, n16175, 
        n16176, n16177, n16178, n16179, n16180, n16181, n16182, 
        n16183, n16184, n16185, n16186, n16187, n16188, n16189, 
        n16190, n16191, n16192, n16193, n16194, n16195, n16196, 
        n16197, n16198, n16199, n16200, n16201, n16202, n16203, 
        n16204, n16205, n16206, n16207, n16208, n16209, n16210, 
        n16211, n16212, n16213, n16214, n16215, n16216, n16217, 
        n16218, n16219, n16220, n16221, n16222, n16223, n16224, 
        n16225, n16226, n16227, n16228, n16229, n16230, n16231, 
        n16232, n16087, n16088, n16089, n16090, n16091, n16092, 
        n16093, n16094, n16095, n16096, n16097, n16098, n16099, 
        n16100, n16101, n16102, n16103, n16104, n16105, n16106, 
        n16107, n16108, n16109, n16110, n16111, n16112, n16113, 
        n16114, n16115, n16116, n16117, n16118, n16119, n16120, 
        n16121, n16122, n16123, n16124, n16125, n16126, n16127, 
        n16128, n16129, n16130, n16131, n16132, n16133, n16134, 
        n16135, n16136, n16137, n16138, n16139, n16140, n16141, 
        n16142, n16143, n16144, n16145, n16146, n16147, n16148, 
        n16149, n16150, n16151, n16152, n16153, n16154, n16155, 
        n16156, n16157, n16158, n16159, n16306, n16307, n16308, 
        n16309, n16310, n16311, n16312, n16313, n16314, n16315, 
        n16316, n16317, n16318, n16319, n16320, n16321, n16322, 
        n16323, n16324, n16325, n16326, n16327, n16328, n16329, 
        n16330, n16331, n16332, n16333, n16334, n16335, n16336, 
        n16337, n16338, n16339, n16340, n16341, n16342, n14776, 
        n14777, n14778, n14779, n14780, n14781, n14782, n14783, 
        n14784, n14785, n14786, n14787, n14788, n14789, n14790, 
        n14791, n14792, n14793, n14794, n14795, n14796, n14797, 
        n14798, n14799, n14800, n14801, n14802, n14803, n14804, 
        n14805, n14806, n14807, n14808, n14809, n14810, n14811, 
        n14812, n14813, n14814, n14815, n14816, n14817, n14818, 
        n14819, n14820, n14821, n14822, n14823, n14824, n14825, 
        n14826, n14827, n14828, n14829, n14830, n14831, n14832, 
        n14833, n14834, n14835, n14836, n14837, n14838, n14839, 
        n14840, n14841, n14842, n14843, n14844, n14845, n14846, 
        n14847, n14848, n14849, n14850, n14851, n14852, n14853, 
        n14854, n14855, n14856, n14857, n14858, n14859, n14860, 
        n14861, n14862, n14863, n14864, n14865, n14866, n14867, 
        n14868, n14869, n14870, n14871, n14872, n14873, n14874, 
        n14875, n14876, n14877, n14878, n14879, n14880, n14881, 
        n14882, n14883, n14884, n14885, n14886, n14887, n14888, 
        n14889, n14890, n14891, n14892, n14893, n14894, n14895, 
        n14896, n14897, n14898, n14899, n14900, n14901, n14902, 
        n14903, n14904, n14905, n14906, n14907, n14908, n14909, 
        n14910, n14911, n14912, n14913, n14914, n14915, n14916, 
        n14917, n14918, n14919, n14920, n14921, n14922, n14923, 
        n14924, n14925, n14926, n14927, n14928, n14929, n14930, 
        n14931, n14932, n14933, n14934, n14935, n14936, n14937, 
        n14938, n14939, n14940, n14941, n14942, n14943, n14944, 
        n14945, n14946, n14947, n14948, n14949, n14950, n14951, 
        n14952, n14953, n14954, n14955, n14956, n14957, n14958, 
        n14630, n14631, n14632, n14633, n14634, n14635, n14636, 
        n14637, n14638, n14639, n14640, n14641, n14642, n14643, 
        n14644, n14645, n14646, n14647, n14648, n14649, n14650, 
        n14651, n14652, n14653, n14654, n14655, n14656, n14657, 
        n14658, n14659, n14660, n14661, n14662, n14663, n14664, 
        n14665, n14666, n14667, n14668, n14669, n14670, n14671, 
        n14672, n14673, n14674, n14675, n14676, n14677, n14678, 
        n14679, n14680, n14681, n14682, n14683, n14684, n14685, 
        n14686, n14687, n14688, n14689, n14690, n14691, n14692, 
        n14693, n14694, n14695, n14696, n14697, n14698, n14699, 
        n14700, n14701, n14702, n14703, n14704, n14705, n14706, 
        n14707, n14708, n14709, n14710, n14711, n14712, n14713, 
        n14714, n14715, n14716, n14717, n14718, n14719, n14720, 
        n14721, n14722, n14723, n14724, n14725, n14726, n14727, 
        n14728, n14729, n14730, n14731, n14732, n14733, n14734, 
        n14735, n14736, n14737, n14738, n14739, n14740, n14741, 
        n14742, n14743, n14744, n14745, n14746, n14747, n14748, 
        n14749, n14750, n14751, n14752, n14753, n14754, n14755, 
        n14756, n14757, n14758, n14759, n14760, n14761, n14762, 
        n14763, n14764, n14765, n14766, n14767, n14768, n14769, 
        n14770, n14771, n14772, n14773, n14774, n14775;
    
    MULT18X18D mult_8 (.A17(dout_i_23__N_5974[17]), .A16(dout_i_23__N_5974[16]), 
            .A15(dout_i_23__N_5974[15]), .A14(dout_i_23__N_5974[14]), .A13(dout_i_23__N_5974[13]), 
            .A12(dout_i_23__N_5974[12]), .A11(dout_i_23__N_5974[11]), .A10(dout_i_23__N_5974[10]), 
            .A9(dout_i_23__N_5974[9]), .A8(dout_i_23__N_5974[8]), .A7(dout_i_23__N_5974[7]), 
            .A6(dout_i_23__N_5974[6]), .A5(dout_i_23__N_5974[5]), .A4(dout_i_23__N_5974[4]), 
            .A3(dout_i_23__N_5974[3]), .A2(dout_i_23__N_5974[2]), .A1(dout_i_23__N_5974[1]), 
            .A0(dout_i_23__N_5974[0]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(VCC_net), .B7(GND_net), 
            .B6(GND_net), .B5(GND_net), .B4(GND_net), .B3(GND_net), 
            .B2(GND_net), .B1(GND_net), .B0(GND_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(n34738), .CE2(GND_net), .CE1(GND_net), 
            .CE0(GND_net), .RST3(rst_n_N_2), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n16031), .ROA16(n16030), .ROA15(n16029), 
            .ROA14(n16028), .ROA13(n16027), .ROA12(n16026), .ROA11(n16025), 
            .ROA10(n16024), .ROA9(n16023), .ROA8(n16022), .ROA7(n16021), 
            .ROA6(n16020), .ROA5(n16019), .ROA4(n16018), .ROA3(n16017), 
            .ROA2(n16016), .ROA1(n16015), .ROA0(n16014), .ROB17(n16049), 
            .ROB16(n16048), .ROB15(n16047), .ROB14(n16046), .ROB13(n16045), 
            .ROB12(n16044), .ROB11(n16043), .ROB10(n16042), .ROB9(n16041), 
            .ROB8(n16040), .ROB7(n16039), .ROB6(n16038), .ROB5(n16037), 
            .ROB4(n16036), .ROB3(n16035), .ROB2(n16034), .ROB1(n16033), 
            .ROB0(n16032), .P35(n16086), .P34(n16085), .P33(n16084), 
            .P32(n16083), .P31(n16082), .P30(n16081), .P29(n16080), 
            .P28(n16079), .P27(n16078), .P26(n16077), .P25(n16076), 
            .P24(n16075), .P23(n16074), .P22(n16073), .P21(n16072), 
            .P20(n16071), .P19(n16070), .P18(n16069), .P17(n16068), 
            .P16(n16067), .P15(n16066), .P14(n16065), .P13(n16064), 
            .P12(n16063), .P11(n16062), .P10(n16061), .P9(n16060), .P8(n16059), 
            .P7(n16058), .P6(n16057), .P5(n16056), .P4(n16055), .P3(n16054), 
            .P2(n16053), .P1(n16052), .P0(n16051), .SIGNEDP(n16050));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam mult_8.REG_INPUTA_CLK = "CLK3";
    defparam mult_8.REG_INPUTA_CE = "CE3";
    defparam mult_8.REG_INPUTA_RST = "RST3";
    defparam mult_8.REG_INPUTB_CLK = "NONE";
    defparam mult_8.REG_INPUTB_CE = "CE0";
    defparam mult_8.REG_INPUTB_RST = "RST0";
    defparam mult_8.REG_INPUTC_CLK = "NONE";
    defparam mult_8.REG_INPUTC_CE = "CE0";
    defparam mult_8.REG_INPUTC_RST = "RST0";
    defparam mult_8.REG_PIPELINE_CLK = "NONE";
    defparam mult_8.REG_PIPELINE_CE = "CE0";
    defparam mult_8.REG_PIPELINE_RST = "RST0";
    defparam mult_8.REG_OUTPUT_CLK = "NONE";
    defparam mult_8.REG_OUTPUT_CE = "CE0";
    defparam mult_8.REG_OUTPUT_RST = "RST0";
    defparam mult_8.CLK0_DIV = "ENABLED";
    defparam mult_8.CLK1_DIV = "ENABLED";
    defparam mult_8.CLK2_DIV = "ENABLED";
    defparam mult_8.CLK3_DIV = "ENABLED";
    defparam mult_8.HIGHSPEED_CLK = "NONE";
    defparam mult_8.GSR = "DISABLED";
    defparam mult_8.CAS_MATCH_REG = "FALSE";
    defparam mult_8.SOURCEB_MODE = "B_SHIFT";
    defparam mult_8.MULT_BYPASS = "DISABLED";
    defparam mult_8.RESETMODE = "ASYNC";
    ALU54B lat_alu_34 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n15504), .SIGNEDIB(n15577), .SIGNEDCIN(n15650), .A35(n15503), 
           .A34(n15502), .A33(n15501), .A32(n15500), .A31(n15499), .A30(n15498), 
           .A29(n15497), .A28(n15496), .A27(n15495), .A26(n15494), .A25(n15493), 
           .A24(n15492), .A23(n15491), .A22(n15490), .A21(n15489), .A20(n15488), 
           .A19(n15487), .A18(n15486), .A17(n15485), .A16(n15484), .A15(n15483), 
           .A14(n15482), .A13(n15481), .A12(n15480), .A11(n15479), .A10(n15478), 
           .A9(n15477), .A8(n15476), .A7(n15475), .A6(n15474), .A5(n15473), 
           .A4(n15472), .A3(n15471), .A2(n15470), .A1(n15469), .A0(n15468), 
           .B35(n15576), .B34(n15575), .B33(n15574), .B32(n15573), .B31(n15572), 
           .B30(n15571), .B29(n15570), .B28(n15569), .B27(n15568), .B26(n15567), 
           .B25(n15566), .B24(n15565), .B23(n15564), .B22(n15563), .B21(n15562), 
           .B20(n15561), .B19(n15560), .B18(n15559), .B17(n15558), .B16(n15557), 
           .B15(n15556), .B14(n15555), .B13(n15554), .B12(n15553), .B11(n15552), 
           .B10(n15551), .B9(n15550), .B8(n15549), .B7(n15548), .B6(n15547), 
           .B5(n15546), .B4(n15545), .B3(n15544), .B2(n15543), .B1(n15542), 
           .B0(n15541), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n15540), .MA34(n15539), .MA33(n15538), .MA32(n15537), 
           .MA31(n15536), .MA30(n15535), .MA29(n15534), .MA28(n15533), 
           .MA27(n15532), .MA26(n15531), .MA25(n15530), .MA24(n15529), 
           .MA23(n15528), .MA22(n15527), .MA21(n15526), .MA20(n15525), 
           .MA19(n15524), .MA18(n15523), .MA17(n15522), .MA16(n15521), 
           .MA15(n15520), .MA14(n15519), .MA13(n15518), .MA12(n15517), 
           .MA11(n15516), .MA10(n15515), .MA9(n15514), .MA8(n15513), 
           .MA7(n15512), .MA6(n15511), .MA5(n15510), .MA4(n15509), .MA3(n15508), 
           .MA2(n15507), .MA1(n15506), .MA0(n15505), .MB35(n15613), 
           .MB34(n15612), .MB33(n15611), .MB32(n15610), .MB31(n15609), 
           .MB30(n15608), .MB29(n15607), .MB28(n15606), .MB27(n15605), 
           .MB26(n15604), .MB25(n15603), .MB24(n15602), .MB23(n15601), 
           .MB22(n15600), .MB21(n15599), .MB20(n15598), .MB19(n15597), 
           .MB18(n15596), .MB17(n15595), .MB16(n15594), .MB15(n15593), 
           .MB14(n15592), .MB13(n15591), .MB12(n15590), .MB11(n15589), 
           .MB10(n15588), .MB9(n15587), .MB8(n15586), .MB7(n15585), 
           .MB6(n15584), .MB5(n15583), .MB4(n15582), .MB3(n15581), .MB2(n15580), 
           .MB1(n15579), .MB0(n15578), .CIN53(n15649), .CIN52(n15648), 
           .CIN51(n15647), .CIN50(n15646), .CIN49(n15645), .CIN48(n15644), 
           .CIN47(n15643), .CIN46(n15642), .CIN45(n15641), .CIN44(n15640), 
           .CIN43(n15639), .CIN42(n15638), .CIN41(n15637), .CIN40(n15636), 
           .CIN39(n15635), .CIN38(n15634), .CIN37(n15633), .CIN36(n15632), 
           .CIN35(n15631), .CIN34(n15630), .CIN33(n15629), .CIN32(n15628), 
           .CIN31(n15627), .CIN30(n15626), .CIN29(n15625), .CIN28(n15624), 
           .CIN27(n15623), .CIN26(n15622), .CIN25(n15621), .CIN24(n15620), 
           .CIN23(n15619), .CIN22(n15618), .CIN21(n15617), .CIN20(n15616), 
           .CIN19(n15615), .CIN18(n15614), .CIN17(\op_r_23__N_1226[17] ), 
           .CIN16(\op_r_23__N_1226[16] ), .CIN15(\op_r_23__N_1226[15] ), 
           .CIN14(\op_r_23__N_1226[14] ), .CIN13(\op_r_23__N_1226[13] ), 
           .CIN12(\op_r_23__N_1226[12] ), .CIN11(\op_r_23__N_1226[11] ), 
           .CIN10(\op_r_23__N_1226[10] ), .CIN9(\op_r_23__N_1226[9] ), .CIN8(\op_r_23__N_1226[8] ), 
           .CIN7(\op_r_23__N_1226[7] ), .CIN6(\op_r_23__N_1226[6] ), .CIN5(\op_r_23__N_1226[5] ), 
           .CIN4(\op_r_23__N_1226[4] ), .CIN3(\op_r_23__N_1226[3] ), .CIN2(\op_r_23__N_1226[2] ), 
           .CIN1(\op_r_23__N_1226[1] ), .CIN0(\op_r_23__N_1226[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1226[31] ), 
           .R12(\op_r_23__N_1226[30] ), .R11(\op_r_23__N_1226[29] ), .R10(\op_r_23__N_1226[28] ), 
           .R9(\op_r_23__N_1226[27] ), .R8(\op_r_23__N_1226[26] ), .R7(\op_r_23__N_1226[25] ), 
           .R6(\op_r_23__N_1226[24] ), .R5(\op_r_23__N_1226[23] ), .R4(\op_r_23__N_1226[22] ), 
           .R3(\op_r_23__N_1226[21] ), .R2(\op_r_23__N_1226[20] ), .R1(\op_r_23__N_1226[19] ), 
           .R0(\op_r_23__N_1226[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_34.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_34.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_34.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_34.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_34.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_34.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_34.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_34.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_34.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_34.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_34.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_34.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_34.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_34.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_34.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_34.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_34.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_34.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_34.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_34.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_34.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_34.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_34.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_34.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_34.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_34.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_34.REG_FLAG_CLK = "NONE";
    defparam lat_alu_34.REG_FLAG_CE = "CE0";
    defparam lat_alu_34.REG_FLAG_RST = "RST0";
    defparam lat_alu_34.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_34.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_34.MASK01 = "0x00000000000000";
    defparam lat_alu_34.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_34.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_34.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_34.CLK0_DIV = "ENABLED";
    defparam lat_alu_34.CLK1_DIV = "ENABLED";
    defparam lat_alu_34.CLK2_DIV = "ENABLED";
    defparam lat_alu_34.CLK3_DIV = "ENABLED";
    defparam lat_alu_34.MCPAT = "0x00000000000000";
    defparam lat_alu_34.MASKPAT = "0x00000000000000";
    defparam lat_alu_34.RNDPAT = "0x00000000000000";
    defparam lat_alu_34.GSR = "DISABLED";
    defparam lat_alu_34.RESETMODE = "SYNC";
    defparam lat_alu_34.MULT9_MODE = "DISABLED";
    defparam lat_alu_34.LEGACY = "DISABLED";
    ALU54B lat_alu_80 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n18747), .SIGNEDIB(n18820), .SIGNEDCIN(GND_net), 
           .A35(n18746), .A34(n18745), .A33(n18744), .A32(n18743), .A31(n18742), 
           .A30(n18741), .A29(n18740), .A28(n18739), .A27(n18738), .A26(n18737), 
           .A25(n18736), .A24(n18735), .A23(n18734), .A22(n18733), .A21(n18732), 
           .A20(n18731), .A19(n18730), .A18(n18729), .A17(n18728), .A16(n18727), 
           .A15(n18726), .A14(n18725), .A13(n18724), .A12(n18723), .A11(n18722), 
           .A10(n18721), .A9(n18720), .A8(n18719), .A7(n18718), .A6(n18717), 
           .A5(n18716), .A4(n18715), .A3(n18714), .A2(n18713), .A1(n18712), 
           .A0(n18711), .B35(n18819), .B34(n18818), .B33(n18817), .B32(n18816), 
           .B31(n18815), .B30(n18814), .B29(n18813), .B28(n18812), .B27(n18811), 
           .B26(n18810), .B25(n18809), .B24(n18808), .B23(n18807), .B22(n18806), 
           .B21(n18805), .B20(n18804), .B19(n18803), .B18(n18802), .B17(n18801), 
           .B16(n18800), .B15(n18799), .B14(n18798), .B13(n18797), .B12(n18796), 
           .B11(n18795), .B10(n18794), .B9(n18793), .B8(n18792), .B7(n18791), 
           .B6(n18790), .B5(n18789), .B4(n18788), .B3(n18787), .B2(n18786), 
           .B1(n18785), .B0(n18784), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n18783), .MA34(n18782), .MA33(n18781), .MA32(n18780), 
           .MA31(n18779), .MA30(n18778), .MA29(n18777), .MA28(n18776), 
           .MA27(n18775), .MA26(n18774), .MA25(n18773), .MA24(n18772), 
           .MA23(n18771), .MA22(n18770), .MA21(n18769), .MA20(n18768), 
           .MA19(n18767), .MA18(n18766), .MA17(n18765), .MA16(n18764), 
           .MA15(n18763), .MA14(n18762), .MA13(n18761), .MA12(n18760), 
           .MA11(n18759), .MA10(n18758), .MA9(n18757), .MA8(n18756), 
           .MA7(n18755), .MA6(n18754), .MA5(n18753), .MA4(n18752), .MA3(n18751), 
           .MA2(n18750), .MA1(n18749), .MA0(n18748), .MB35(n18856), 
           .MB34(n18855), .MB33(n18854), .MB32(n18853), .MB31(n18852), 
           .MB30(n18851), .MB29(n18850), .MB28(n18849), .MB27(n18848), 
           .MB26(n18847), .MB25(n18846), .MB24(n18845), .MB23(n18844), 
           .MB22(n18843), .MB21(n18842), .MB20(n18841), .MB19(n18840), 
           .MB18(n18839), .MB17(n18838), .MB16(n18837), .MB15(n18836), 
           .MB14(n18835), .MB13(n18834), .MB12(n18833), .MB11(n18832), 
           .MB10(n18831), .MB9(n18830), .MB8(n18829), .MB7(n18828), 
           .MB6(n18827), .MB5(n18826), .MB4(n18825), .MB3(n18824), .MB2(n18823), 
           .MB1(n18822), .MB0(n18821), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R30(n65), .R29(n66), 
           .R28(n67), .R27(n68), .R26(n69), .R25(n70), .R24(n71), 
           .R23(n72), .R22(n73), .R21(n74), .R20(n75), .R19(n76), 
           .R18(n77), .R17(n78), .R16(n79), .R15(n80), .R14(n81), 
           .R13(n82), .R12(n83), .R11(n84), .R10(n85), .R9(n86), .R8(n87), 
           .R7(n88), .R6(n89), .R5(\op_i_23__N_1310[5] ), .R4(\op_i_23__N_1310[4] ), 
           .R3(\op_i_23__N_1310[3] ), .R2(\op_i_23__N_1310[2] ), .R1(\op_i_23__N_1310[1] ), 
           .R0(\op_i_23__N_1310[0] ));
    defparam lat_alu_80.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_80.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_80.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_80.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_80.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_80.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_80.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_80.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_80.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_80.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_80.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_80.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_80.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_80.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_80.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_80.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_80.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_80.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_80.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_80.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_80.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_80.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_80.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_80.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_80.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_80.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_80.REG_FLAG_CLK = "NONE";
    defparam lat_alu_80.REG_FLAG_CE = "CE0";
    defparam lat_alu_80.REG_FLAG_RST = "RST0";
    defparam lat_alu_80.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_80.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_80.MASK01 = "0x00000000000000";
    defparam lat_alu_80.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_80.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_80.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_80.CLK0_DIV = "ENABLED";
    defparam lat_alu_80.CLK1_DIV = "ENABLED";
    defparam lat_alu_80.CLK2_DIV = "ENABLED";
    defparam lat_alu_80.CLK3_DIV = "ENABLED";
    defparam lat_alu_80.MCPAT = "0x00000000000000";
    defparam lat_alu_80.MASKPAT = "0x00000000000000";
    defparam lat_alu_80.RNDPAT = "0x00000000000000";
    defparam lat_alu_80.GSR = "DISABLED";
    defparam lat_alu_80.RESETMODE = "SYNC";
    defparam lat_alu_80.MULT9_MODE = "DISABLED";
    defparam lat_alu_80.LEGACY = "DISABLED";
    MULT18X18D lat_mult_79 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(GND_net), 
            .B16(GND_net), .B15(GND_net), .B14(GND_net), .B13(GND_net), 
            .B12(GND_net), .B11(GND_net), .B10(GND_net), .B9(GND_net), 
            .B8(GND_net), .B7(GND_net), .B6(GND_net), .B5(n11561), .B4(n11560), 
            .B3(n11559), .B2(n11558), .B1(n11557), .B0(n11556), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n18801), .ROA16(n18800), .ROA15(n18799), 
            .ROA14(n18798), .ROA13(n18797), .ROA12(n18796), .ROA11(n18795), 
            .ROA10(n18794), .ROA9(n18793), .ROA8(n18792), .ROA7(n18791), 
            .ROA6(n18790), .ROA5(n18789), .ROA4(n18788), .ROA3(n18787), 
            .ROA2(n18786), .ROA1(n18785), .ROA0(n18784), .ROB17(n18819), 
            .ROB16(n18818), .ROB15(n18817), .ROB14(n18816), .ROB13(n18815), 
            .ROB12(n18814), .ROB11(n18813), .ROB10(n18812), .ROB9(n18811), 
            .ROB8(n18810), .ROB7(n18809), .ROB6(n18808), .ROB5(n18807), 
            .ROB4(n18806), .ROB3(n18805), .ROB2(n18804), .ROB1(n18803), 
            .ROB0(n18802), .P35(n18856), .P34(n18855), .P33(n18854), 
            .P32(n18853), .P31(n18852), .P30(n18851), .P29(n18850), 
            .P28(n18849), .P27(n18848), .P26(n18847), .P25(n18846), 
            .P24(n18845), .P23(n18844), .P22(n18843), .P21(n18842), 
            .P20(n18841), .P19(n18840), .P18(n18839), .P17(n18838), 
            .P16(n18837), .P15(n18836), .P14(n18835), .P13(n18834), 
            .P12(n18833), .P11(n18832), .P10(n18831), .P9(n18830), .P8(n18829), 
            .P7(n18828), .P6(n18827), .P5(n18826), .P4(n18825), .P3(n18824), 
            .P2(n18823), .P1(n18822), .P0(n18821), .SIGNEDP(n18820));
    defparam lat_mult_79.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_79.REG_INPUTA_CE = "CE0";
    defparam lat_mult_79.REG_INPUTA_RST = "RST0";
    defparam lat_mult_79.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_79.REG_INPUTB_CE = "CE0";
    defparam lat_mult_79.REG_INPUTB_RST = "RST0";
    defparam lat_mult_79.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_79.REG_INPUTC_CE = "CE0";
    defparam lat_mult_79.REG_INPUTC_RST = "RST0";
    defparam lat_mult_79.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_79.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_79.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_79.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_79.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_79.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_79.CLK0_DIV = "ENABLED";
    defparam lat_mult_79.CLK1_DIV = "ENABLED";
    defparam lat_mult_79.CLK2_DIV = "ENABLED";
    defparam lat_mult_79.CLK3_DIV = "ENABLED";
    defparam lat_mult_79.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_79.GSR = "DISABLED";
    defparam lat_mult_79.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_79.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_79.MULT_BYPASS = "DISABLED";
    defparam lat_mult_79.RESETMODE = "SYNC";
    ALU54B lat_alu_33 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n15358), .SIGNEDIB(n15431), .SIGNEDCIN(GND_net), 
           .A35(n15357), .A34(n15356), .A33(n15355), .A32(n15354), .A31(n15353), 
           .A30(n15352), .A29(n15351), .A28(n15350), .A27(n15349), .A26(n15348), 
           .A25(n15347), .A24(n15346), .A23(n15345), .A22(n15344), .A21(n15343), 
           .A20(n15342), .A19(n15341), .A18(n15340), .A17(n15339), .A16(n15338), 
           .A15(n15337), .A14(n15336), .A13(n15335), .A12(n15334), .A11(n15333), 
           .A10(n15332), .A9(n15331), .A8(n15330), .A7(n15329), .A6(n15328), 
           .A5(n15327), .A4(n15326), .A3(n15325), .A2(n15324), .A1(n15323), 
           .A0(n15322), .B35(n15430), .B34(n15429), .B33(n15428), .B32(n15427), 
           .B31(n15426), .B30(n15425), .B29(n15424), .B28(n15423), .B27(n15422), 
           .B26(n15421), .B25(n15420), .B24(n15419), .B23(n15418), .B22(n15417), 
           .B21(n15416), .B20(n15415), .B19(n15414), .B18(n15413), .B17(n15412), 
           .B16(n15411), .B15(n15410), .B14(n15409), .B13(n15408), .B12(n15407), 
           .B11(n15406), .B10(n15405), .B9(n15404), .B8(n15403), .B7(n15402), 
           .B6(n15401), .B5(n15400), .B4(n15399), .B3(n15398), .B2(n15397), 
           .B1(n15396), .B0(n15395), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n15394), .MA34(n15393), .MA33(n15392), .MA32(n15391), 
           .MA31(n15390), .MA30(n15389), .MA29(n15388), .MA28(n15387), 
           .MA27(n15386), .MA26(n15385), .MA25(n15384), .MA24(n15383), 
           .MA23(n15382), .MA22(n15381), .MA21(n15380), .MA20(n15379), 
           .MA19(n15378), .MA18(n15377), .MA17(n15376), .MA16(n15375), 
           .MA15(n15374), .MA14(n15373), .MA13(n15372), .MA12(n15371), 
           .MA11(n15370), .MA10(n15369), .MA9(n15368), .MA8(n15367), 
           .MA7(n15366), .MA6(n15365), .MA5(n15364), .MA4(n15363), .MA3(n15362), 
           .MA2(n15361), .MA1(n15360), .MA0(n15359), .MB35(n15467), 
           .MB34(n15466), .MB33(n15465), .MB32(n15464), .MB31(n15463), 
           .MB30(n15462), .MB29(n15461), .MB28(n15460), .MB27(n15459), 
           .MB26(n15458), .MB25(n15457), .MB24(n15456), .MB23(n15455), 
           .MB22(n15454), .MB21(n15453), .MB20(n15452), .MB19(n15451), 
           .MB18(n15450), .MB17(n15449), .MB16(n15448), .MB15(n15447), 
           .MB14(n15446), .MB13(n15445), .MB12(n15444), .MB11(n15443), 
           .MB10(n15442), .MB9(n15441), .MB8(n15440), .MB7(n15439), 
           .MB6(n15438), .MB5(n15437), .MB4(n15436), .MB3(n15435), .MB2(n15434), 
           .MB1(n15433), .MB0(n15432), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n15649), 
           .R52(n15648), .R51(n15647), .R50(n15646), .R49(n15645), .R48(n15644), 
           .R47(n15643), .R46(n15642), .R45(n15641), .R44(n15640), .R43(n15639), 
           .R42(n15638), .R41(n15637), .R40(n15636), .R39(n15635), .R38(n15634), 
           .R37(n15633), .R36(n15632), .R35(n15631), .R34(n15630), .R33(n15629), 
           .R32(n15628), .R31(n15627), .R30(n15626), .R29(n15625), .R28(n15624), 
           .R27(n15623), .R26(n15622), .R25(n15621), .R24(n15620), .R23(n15619), 
           .R22(n15618), .R21(n15617), .R20(n15616), .R19(n15615), .R18(n15614), 
           .R17(\op_r_23__N_1226[17] ), .R16(\op_r_23__N_1226[16] ), .R15(\op_r_23__N_1226[15] ), 
           .R14(\op_r_23__N_1226[14] ), .R13(\op_r_23__N_1226[13] ), .R12(\op_r_23__N_1226[12] ), 
           .R11(\op_r_23__N_1226[11] ), .R10(\op_r_23__N_1226[10] ), .R9(\op_r_23__N_1226[9] ), 
           .R8(\op_r_23__N_1226[8] ), .R7(\op_r_23__N_1226[7] ), .R6(\op_r_23__N_1226[6] ), 
           .R5(\op_r_23__N_1226[5] ), .R4(\op_r_23__N_1226[4] ), .R3(\op_r_23__N_1226[3] ), 
           .R2(\op_r_23__N_1226[2] ), .R1(\op_r_23__N_1226[1] ), .R0(\op_r_23__N_1226[0] ), 
           .SIGNEDR(n15650));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_alu_33.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_33.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_33.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_33.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_33.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_33.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_33.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_33.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_33.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_33.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_33.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_33.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_33.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_33.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_33.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_33.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_33.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_33.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_33.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_33.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_33.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_33.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_33.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_33.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_33.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_33.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_33.REG_FLAG_CLK = "NONE";
    defparam lat_alu_33.REG_FLAG_CE = "CE0";
    defparam lat_alu_33.REG_FLAG_RST = "RST0";
    defparam lat_alu_33.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_33.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_33.MASK01 = "0x00000000000000";
    defparam lat_alu_33.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_33.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_33.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_33.CLK0_DIV = "ENABLED";
    defparam lat_alu_33.CLK1_DIV = "ENABLED";
    defparam lat_alu_33.CLK2_DIV = "ENABLED";
    defparam lat_alu_33.CLK3_DIV = "ENABLED";
    defparam lat_alu_33.MCPAT = "0x00000000000000";
    defparam lat_alu_33.MASKPAT = "0x00000000000000";
    defparam lat_alu_33.RNDPAT = "0x00000000000000";
    defparam lat_alu_33.GSR = "DISABLED";
    defparam lat_alu_33.RESETMODE = "SYNC";
    defparam lat_alu_33.MULT9_MODE = "DISABLED";
    defparam lat_alu_33.LEGACY = "DISABLED";
    MULT18X18D lat_mult_32 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12089), 
            .B16(n12089), .B15(n12089), .B14(n12089), .B13(n12089), 
            .B12(n12089), .B11(n12089), .B10(n12089), .B9(n12089), .B8(n12089), 
            .B7(n12089), .B6(n12089), .B5(n12088), .B4(n12087), .B3(n12086), 
            .B2(n12085), .B1(n12084), .B0(n12083), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15558), .ROA16(n15557), .ROA15(n15556), .ROA14(n15555), 
            .ROA13(n15554), .ROA12(n15553), .ROA11(n15552), .ROA10(n15551), 
            .ROA9(n15550), .ROA8(n15549), .ROA7(n15548), .ROA6(n15547), 
            .ROA5(n15546), .ROA4(n15545), .ROA3(n15544), .ROA2(n15543), 
            .ROA1(n15542), .ROA0(n15541), .ROB17(n15576), .ROB16(n15575), 
            .ROB15(n15574), .ROB14(n15573), .ROB13(n15572), .ROB12(n15571), 
            .ROB11(n15570), .ROB10(n15569), .ROB9(n15568), .ROB8(n15567), 
            .ROB7(n15566), .ROB6(n15565), .ROB5(n15564), .ROB4(n15563), 
            .ROB3(n15562), .ROB2(n15561), .ROB1(n15560), .ROB0(n15559), 
            .P35(n15613), .P34(n15612), .P33(n15611), .P32(n15610), 
            .P31(n15609), .P30(n15608), .P29(n15607), .P28(n15606), 
            .P27(n15605), .P26(n15604), .P25(n15603), .P24(n15602), 
            .P23(n15601), .P22(n15600), .P21(n15599), .P20(n15598), 
            .P19(n15597), .P18(n15596), .P17(n15595), .P16(n15594), 
            .P15(n15593), .P14(n15592), .P13(n15591), .P12(n15590), 
            .P11(n15589), .P10(n15588), .P9(n15587), .P8(n15586), .P7(n15585), 
            .P6(n15584), .P5(n15583), .P4(n15582), .P3(n15581), .P2(n15580), 
            .P1(n15579), .P0(n15578), .SIGNEDP(n15577));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_32.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_32.REG_INPUTA_CE = "CE0";
    defparam lat_mult_32.REG_INPUTA_RST = "RST0";
    defparam lat_mult_32.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_32.REG_INPUTB_CE = "CE0";
    defparam lat_mult_32.REG_INPUTB_RST = "RST0";
    defparam lat_mult_32.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_32.REG_INPUTC_CE = "CE0";
    defparam lat_mult_32.REG_INPUTC_RST = "RST0";
    defparam lat_mult_32.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_32.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_32.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_32.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_32.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_32.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_32.CLK0_DIV = "ENABLED";
    defparam lat_mult_32.CLK1_DIV = "ENABLED";
    defparam lat_mult_32.CLK2_DIV = "ENABLED";
    defparam lat_mult_32.CLK3_DIV = "ENABLED";
    defparam lat_mult_32.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_32.GSR = "DISABLED";
    defparam lat_mult_32.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_32.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_32.MULT_BYPASS = "DISABLED";
    defparam lat_mult_32.RESETMODE = "SYNC";
    MULT18X18D lat_mult_31 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(VCC_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12089), 
            .B16(n12089), .B15(n12089), .B14(n12089), .B13(n12089), 
            .B12(n12089), .B11(n12089), .B10(n12089), .B9(n12089), .B8(n12089), 
            .B7(n12089), .B6(n12089), .B5(n12088), .B4(n12087), .B3(n12086), 
            .B2(n12085), .B1(n12084), .B0(n12083), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15485), .ROA16(n15484), .ROA15(n15483), .ROA14(n15482), 
            .ROA13(n15481), .ROA12(n15480), .ROA11(n15479), .ROA10(n15478), 
            .ROA9(n15477), .ROA8(n15476), .ROA7(n15475), .ROA6(n15474), 
            .ROA5(n15473), .ROA4(n15472), .ROA3(n15471), .ROA2(n15470), 
            .ROA1(n15469), .ROA0(n15468), .ROB17(n15503), .ROB16(n15502), 
            .ROB15(n15501), .ROB14(n15500), .ROB13(n15499), .ROB12(n15498), 
            .ROB11(n15497), .ROB10(n15496), .ROB9(n15495), .ROB8(n15494), 
            .ROB7(n15493), .ROB6(n15492), .ROB5(n15491), .ROB4(n15490), 
            .ROB3(n15489), .ROB2(n15488), .ROB1(n15487), .ROB0(n15486), 
            .P35(n15540), .P34(n15539), .P33(n15538), .P32(n15537), 
            .P31(n15536), .P30(n15535), .P29(n15534), .P28(n15533), 
            .P27(n15532), .P26(n15531), .P25(n15530), .P24(n15529), 
            .P23(n15528), .P22(n15527), .P21(n15526), .P20(n15525), 
            .P19(n15524), .P18(n15523), .P17(n15522), .P16(n15521), 
            .P15(n15520), .P14(n15519), .P13(n15518), .P12(n15517), 
            .P11(n15516), .P10(n15515), .P9(n15514), .P8(n15513), .P7(n15512), 
            .P6(n15511), .P5(n15510), .P4(n15509), .P3(n15508), .P2(n15507), 
            .P1(n15506), .P0(n15505), .SIGNEDP(n15504));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_31.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_31.REG_INPUTA_CE = "CE0";
    defparam lat_mult_31.REG_INPUTA_RST = "RST0";
    defparam lat_mult_31.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_31.REG_INPUTB_CE = "CE0";
    defparam lat_mult_31.REG_INPUTB_RST = "RST0";
    defparam lat_mult_31.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_31.REG_INPUTC_CE = "CE0";
    defparam lat_mult_31.REG_INPUTC_RST = "RST0";
    defparam lat_mult_31.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_31.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_31.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_31.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_31.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_31.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_31.CLK0_DIV = "ENABLED";
    defparam lat_mult_31.CLK1_DIV = "ENABLED";
    defparam lat_mult_31.CLK2_DIV = "ENABLED";
    defparam lat_mult_31.CLK3_DIV = "ENABLED";
    defparam lat_mult_31.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_31.GSR = "DISABLED";
    defparam lat_mult_31.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_31.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_31.MULT_BYPASS = "DISABLED";
    defparam lat_mult_31.RESETMODE = "SYNC";
    MULT18X18D lat_mult_42 (.A17(dout_i_23__N_5974[23]), .A16(dout_i_23__N_5974[23]), 
            .A15(dout_i_23__N_5974[23]), .A14(dout_i_23__N_5974[23]), .A13(dout_i_23__N_5974[23]), 
            .A12(dout_i_23__N_5974[23]), .A11(dout_i_23__N_5974[23]), .A10(dout_i_23__N_5974[23]), 
            .A9(dout_i_23__N_5974[23]), .A8(dout_i_23__N_5974[23]), .A7(dout_i_23__N_5974[23]), 
            .A6(dout_i_23__N_5974[23]), .A5(dout_i_23__N_5974[23]), .A4(dout_i_23__N_5974[22]), 
            .A3(dout_i_23__N_5974[21]), .A2(dout_i_23__N_5974[20]), .A1(dout_i_23__N_5974[19]), 
            .A0(dout_i_23__N_5974[18]), .B17(GND_net), .B16(GND_net), 
            .B15(GND_net), .B14(GND_net), .B13(GND_net), .B12(GND_net), 
            .B11(GND_net), .B10(GND_net), .B9(GND_net), .B8(GND_net), 
            .B7(GND_net), .B6(GND_net), .B5(GND_net), .B4(GND_net), 
            .B3(GND_net), .B2(GND_net), .B1(GND_net), .B0(GND_net), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(n34738), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(rst_n_N_2), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n16250), .ROA16(n16249), 
            .ROA15(n16248), .ROA14(n16247), .ROA13(n16246), .ROA12(n16245), 
            .ROA11(n16244), .ROA10(n16243), .ROA9(n16242), .ROA8(n16241), 
            .ROA7(n16240), .ROA6(n16239), .ROA5(n16238), .ROA4(n16237), 
            .ROA3(n16236), .ROA2(n16235), .ROA1(n16234), .ROA0(n16233), 
            .ROB17(n16268), .ROB16(n16267), .ROB15(n16266), .ROB14(n16265), 
            .ROB13(n16264), .ROB12(n16263), .ROB11(n16262), .ROB10(n16261), 
            .ROB9(n16260), .ROB8(n16259), .ROB7(n16258), .ROB6(n16257), 
            .ROB5(n16256), .ROB4(n16255), .ROB3(n16254), .ROB2(n16253), 
            .ROB1(n16252), .ROB0(n16251), .P35(n16305), .P34(n16304), 
            .P33(n16303), .P32(n16302), .P31(n16301), .P30(n16300), 
            .P29(n16299), .P28(n16298), .P27(n16297), .P26(n16296), 
            .P25(n16295), .P24(n16294), .P23(n16293), .P22(n16292), 
            .P21(n16291), .P20(n16290), .P19(n16289), .P18(n16288), 
            .P17(n16287), .P16(n16286), .P15(n16285), .P14(n16284), 
            .P13(n16283), .P12(n16282), .P11(n16281), .P10(n16280), 
            .P9(n16279), .P8(n16278), .P7(n16277), .P6(n16276), .P5(n16275), 
            .P4(n16274), .P3(n16273), .P2(n16272), .P1(n16271), .P0(n16270), 
            .SIGNEDP(n16269));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_42.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_42.REG_INPUTA_CE = "CE3";
    defparam lat_mult_42.REG_INPUTA_RST = "RST3";
    defparam lat_mult_42.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_42.REG_INPUTB_CE = "CE0";
    defparam lat_mult_42.REG_INPUTB_RST = "RST0";
    defparam lat_mult_42.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_42.REG_INPUTC_CE = "CE0";
    defparam lat_mult_42.REG_INPUTC_RST = "RST0";
    defparam lat_mult_42.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_42.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_42.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_42.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_42.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_42.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_42.CLK0_DIV = "ENABLED";
    defparam lat_mult_42.CLK1_DIV = "ENABLED";
    defparam lat_mult_42.CLK2_DIV = "ENABLED";
    defparam lat_mult_42.CLK3_DIV = "ENABLED";
    defparam lat_mult_42.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_42.GSR = "DISABLED";
    defparam lat_mult_42.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_42.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_42.MULT_BYPASS = "DISABLED";
    defparam lat_mult_42.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_30 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12082), 
            .B16(n12081), .B15(n12080), .B14(n12079), .B13(n12078), 
            .B12(n12077), .B11(n12076), .B10(n12075), .B9(n12074), .B8(n12073), 
            .B7(n12072), .B6(n12071), .B5(n12070), .B4(n12069), .B3(n12068), 
            .B2(n12067), .B1(n12066), .B0(n12065), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15412), .ROA16(n15411), .ROA15(n15410), .ROA14(n15409), 
            .ROA13(n15408), .ROA12(n15407), .ROA11(n15406), .ROA10(n15405), 
            .ROA9(n15404), .ROA8(n15403), .ROA7(n15402), .ROA6(n15401), 
            .ROA5(n15400), .ROA4(n15399), .ROA3(n15398), .ROA2(n15397), 
            .ROA1(n15396), .ROA0(n15395), .ROB17(n15430), .ROB16(n15429), 
            .ROB15(n15428), .ROB14(n15427), .ROB13(n15426), .ROB12(n15425), 
            .ROB11(n15424), .ROB10(n15423), .ROB9(n15422), .ROB8(n15421), 
            .ROB7(n15420), .ROB6(n15419), .ROB5(n15418), .ROB4(n15417), 
            .ROB3(n15416), .ROB2(n15415), .ROB1(n15414), .ROB0(n15413), 
            .P35(n15467), .P34(n15466), .P33(n15465), .P32(n15464), 
            .P31(n15463), .P30(n15462), .P29(n15461), .P28(n15460), 
            .P27(n15459), .P26(n15458), .P25(n15457), .P24(n15456), 
            .P23(n15455), .P22(n15454), .P21(n15453), .P20(n15452), 
            .P19(n15451), .P18(n15450), .P17(n15449), .P16(n15448), 
            .P15(n15447), .P14(n15446), .P13(n15445), .P12(n15444), 
            .P11(n15443), .P10(n15442), .P9(n15441), .P8(n15440), .P7(n15439), 
            .P6(n15438), .P5(n15437), .P4(n15436), .P3(n15435), .P2(n15434), 
            .P1(n15433), .P0(n15432), .SIGNEDP(n15431));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam lat_mult_30.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_30.REG_INPUTA_CE = "CE0";
    defparam lat_mult_30.REG_INPUTA_RST = "RST0";
    defparam lat_mult_30.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_30.REG_INPUTB_CE = "CE0";
    defparam lat_mult_30.REG_INPUTB_RST = "RST0";
    defparam lat_mult_30.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_30.REG_INPUTC_CE = "CE0";
    defparam lat_mult_30.REG_INPUTC_RST = "RST0";
    defparam lat_mult_30.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_30.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_30.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_30.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_30.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_30.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_30.CLK0_DIV = "ENABLED";
    defparam lat_mult_30.CLK1_DIV = "ENABLED";
    defparam lat_mult_30.CLK2_DIV = "ENABLED";
    defparam lat_mult_30.CLK3_DIV = "ENABLED";
    defparam lat_mult_30.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_30.GSR = "DISABLED";
    defparam lat_mult_30.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_30.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_30.MULT_BYPASS = "DISABLED";
    defparam lat_mult_30.RESETMODE = "SYNC";
    MULT18X18D mult_979_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(GND_net), 
            .B16(GND_net), .B15(GND_net), .B14(GND_net), .B13(GND_net), 
            .B12(GND_net), .B11(GND_net), .B10(GND_net), .B9(GND_net), 
            .B8(GND_net), .B7(GND_net), .B6(GND_net), .B5(n11561), .B4(n11560), 
            .B3(n11559), .B2(n11558), .B1(n11557), .B0(n11556), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n18728), .ROA16(n18727), .ROA15(n18726), 
            .ROA14(n18725), .ROA13(n18724), .ROA12(n18723), .ROA11(n18722), 
            .ROA10(n18721), .ROA9(n18720), .ROA8(n18719), .ROA7(n18718), 
            .ROA6(n18717), .ROA5(n18716), .ROA4(n18715), .ROA3(n18714), 
            .ROA2(n18713), .ROA1(n18712), .ROA0(n18711), .ROB17(n18746), 
            .ROB16(n18745), .ROB15(n18744), .ROB14(n18743), .ROB13(n18742), 
            .ROB12(n18741), .ROB11(n18740), .ROB10(n18739), .ROB9(n18738), 
            .ROB8(n18737), .ROB7(n18736), .ROB6(n18735), .ROB5(n18734), 
            .ROB4(n18733), .ROB3(n18732), .ROB2(n18731), .ROB1(n18730), 
            .ROB0(n18729), .P35(n18783), .P34(n18782), .P33(n18781), 
            .P32(n18780), .P31(n18779), .P30(n18778), .P29(n18777), 
            .P28(n18776), .P27(n18775), .P26(n18774), .P25(n18773), 
            .P24(n18772), .P23(n18771), .P22(n18770), .P21(n18769), 
            .P20(n18768), .P19(n18767), .P18(n18766), .P17(n18765), 
            .P16(n18764), .P15(n18763), .P14(n18762), .P13(n18761), 
            .P12(n18760), .P11(n18759), .P10(n18758), .P9(n18757), .P8(n18756), 
            .P7(n18755), .P6(n18754), .P5(n18753), .P4(n18752), .P3(n18751), 
            .P2(n18750), .P1(n18749), .P0(n18748), .SIGNEDP(n18747));
    defparam mult_979_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_979_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_979_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_979_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_979_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_979_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_979_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_979_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_979_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_979_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_979_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_979_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_979_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_979_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_979_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_979_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_979_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_979_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_979_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_979_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_979_mult_2.GSR = "DISABLED";
    defparam mult_979_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_979_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_979_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_979_mult_2.RESETMODE = "SYNC";
    MULT18X18D mult_10_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(VCC_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n12082), 
            .B16(n12081), .B15(n12080), .B14(n12079), .B13(n12078), 
            .B12(n12077), .B11(n12076), .B10(n12075), .B9(n12074), .B8(n12073), 
            .B7(n12072), .B6(n12071), .B5(n12070), .B4(n12069), .B3(n12068), 
            .B2(n12067), .B1(n12066), .B0(n12065), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n15339), .ROA16(n15338), .ROA15(n15337), .ROA14(n15336), 
            .ROA13(n15335), .ROA12(n15334), .ROA11(n15333), .ROA10(n15332), 
            .ROA9(n15331), .ROA8(n15330), .ROA7(n15329), .ROA6(n15328), 
            .ROA5(n15327), .ROA4(n15326), .ROA3(n15325), .ROA2(n15324), 
            .ROA1(n15323), .ROA0(n15322), .ROB17(n15357), .ROB16(n15356), 
            .ROB15(n15355), .ROB14(n15354), .ROB13(n15353), .ROB12(n15352), 
            .ROB11(n15351), .ROB10(n15350), .ROB9(n15349), .ROB8(n15348), 
            .ROB7(n15347), .ROB6(n15346), .ROB5(n15345), .ROB4(n15344), 
            .ROB3(n15343), .ROB2(n15342), .ROB1(n15341), .ROB0(n15340), 
            .P35(n15394), .P34(n15393), .P33(n15392), .P32(n15391), 
            .P31(n15390), .P30(n15389), .P29(n15388), .P28(n15387), 
            .P27(n15386), .P26(n15385), .P25(n15384), .P24(n15383), 
            .P23(n15382), .P22(n15381), .P21(n15380), .P20(n15379), 
            .P19(n15378), .P18(n15377), .P17(n15376), .P16(n15375), 
            .P15(n15374), .P14(n15373), .P13(n15372), .P12(n15371), 
            .P11(n15370), .P10(n15369), .P9(n15368), .P8(n15367), .P7(n15366), 
            .P6(n15365), .P5(n15364), .P4(n15363), .P3(n15362), .P2(n15361), 
            .P1(n15360), .P0(n15359), .SIGNEDP(n15358));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(53[14:27])
    defparam mult_10_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_10_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_10_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_10_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_10_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_10_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_10_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_10_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_10_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_10_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_10_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_10_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_10_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_10_mult_2.GSR = "DISABLED";
    defparam mult_10_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_10_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_10_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_10_mult_2.RESETMODE = "SYNC";
    MULT18X18D lat_mult_41 (.A17(dout_i_23__N_5974[17]), .A16(dout_i_23__N_5974[16]), 
            .A15(dout_i_23__N_5974[15]), .A14(dout_i_23__N_5974[14]), .A13(dout_i_23__N_5974[13]), 
            .A12(dout_i_23__N_5974[12]), .A11(dout_i_23__N_5974[11]), .A10(dout_i_23__N_5974[10]), 
            .A9(dout_i_23__N_5974[9]), .A8(dout_i_23__N_5974[8]), .A7(dout_i_23__N_5974[7]), 
            .A6(dout_i_23__N_5974[6]), .A5(dout_i_23__N_5974[5]), .A4(dout_i_23__N_5974[4]), 
            .A3(dout_i_23__N_5974[3]), .A2(dout_i_23__N_5974[2]), .A1(dout_i_23__N_5974[1]), 
            .A0(dout_i_23__N_5974[0]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(GND_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(GND_net), .B7(GND_net), 
            .B6(GND_net), .B5(GND_net), .B4(GND_net), .B3(GND_net), 
            .B2(GND_net), .B1(GND_net), .B0(GND_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(n34738), .CE2(GND_net), .CE1(GND_net), 
            .CE0(GND_net), .RST3(rst_n_N_2), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n16177), .ROA16(n16176), .ROA15(n16175), 
            .ROA14(n16174), .ROA13(n16173), .ROA12(n16172), .ROA11(n16171), 
            .ROA10(n16170), .ROA9(n16169), .ROA8(n16168), .ROA7(n16167), 
            .ROA6(n16166), .ROA5(n16165), .ROA4(n16164), .ROA3(n16163), 
            .ROA2(n16162), .ROA1(n16161), .ROA0(n16160), .ROB17(n16195), 
            .ROB16(n16194), .ROB15(n16193), .ROB14(n16192), .ROB13(n16191), 
            .ROB12(n16190), .ROB11(n16189), .ROB10(n16188), .ROB9(n16187), 
            .ROB8(n16186), .ROB7(n16185), .ROB6(n16184), .ROB5(n16183), 
            .ROB4(n16182), .ROB3(n16181), .ROB2(n16180), .ROB1(n16179), 
            .ROB0(n16178), .P35(n16232), .P34(n16231), .P33(n16230), 
            .P32(n16229), .P31(n16228), .P30(n16227), .P29(n16226), 
            .P28(n16225), .P27(n16224), .P26(n16223), .P25(n16222), 
            .P24(n16221), .P23(n16220), .P22(n16219), .P21(n16218), 
            .P20(n16217), .P19(n16216), .P18(n16215), .P17(n16214), 
            .P16(n16213), .P15(n16212), .P14(n16211), .P13(n16210), 
            .P12(n16209), .P11(n16208), .P10(n16207), .P9(n16206), .P8(n16205), 
            .P7(n16204), .P6(n16203), .P5(n16202), .P4(n16201), .P3(n16200), 
            .P2(n16199), .P1(n16198), .P0(n16197), .SIGNEDP(n16196));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_41.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_41.REG_INPUTA_CE = "CE3";
    defparam lat_mult_41.REG_INPUTA_RST = "RST3";
    defparam lat_mult_41.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_41.REG_INPUTB_CE = "CE0";
    defparam lat_mult_41.REG_INPUTB_RST = "RST0";
    defparam lat_mult_41.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_41.REG_INPUTC_CE = "CE0";
    defparam lat_mult_41.REG_INPUTC_RST = "RST0";
    defparam lat_mult_41.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_41.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_41.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_41.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_41.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_41.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_41.CLK0_DIV = "ENABLED";
    defparam lat_mult_41.CLK1_DIV = "ENABLED";
    defparam lat_mult_41.CLK2_DIV = "ENABLED";
    defparam lat_mult_41.CLK3_DIV = "ENABLED";
    defparam lat_mult_41.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_41.GSR = "DISABLED";
    defparam lat_mult_41.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_41.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_41.MULT_BYPASS = "DISABLED";
    defparam lat_mult_41.RESETMODE = "ASYNC";
    ALU54B lat_alu_43 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n16050), .SIGNEDIB(n16123), .SIGNEDCIN(GND_net), 
           .A35(n16049), .A34(n16048), .A33(n16047), .A32(n16046), .A31(n16045), 
           .A30(n16044), .A29(n16043), .A28(n16042), .A27(n16041), .A26(n16040), 
           .A25(n16039), .A24(n16038), .A23(n16037), .A22(n16036), .A21(n16035), 
           .A20(n16034), .A19(n16033), .A18(n16032), .A17(n16031), .A16(n16030), 
           .A15(n16029), .A14(n16028), .A13(n16027), .A12(n16026), .A11(n16025), 
           .A10(n16024), .A9(n16023), .A8(n16022), .A7(n16021), .A6(n16020), 
           .A5(n16019), .A4(n16018), .A3(n16017), .A2(n16016), .A1(n16015), 
           .A0(n16014), .B35(n16122), .B34(n16121), .B33(n16120), .B32(n16119), 
           .B31(n16118), .B30(n16117), .B29(n16116), .B28(n16115), .B27(n16114), 
           .B26(n16113), .B25(n16112), .B24(n16111), .B23(n16110), .B22(n16109), 
           .B21(n16108), .B20(n16107), .B19(n16106), .B18(n16105), .B17(n16104), 
           .B16(n16103), .B15(n16102), .B14(n16101), .B13(n16100), .B12(n16099), 
           .B11(n16098), .B10(n16097), .B9(n16096), .B8(n16095), .B7(n16094), 
           .B6(n16093), .B5(n16092), .B4(n16091), .B3(n16090), .B2(n16089), 
           .B1(n16088), .B0(n16087), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n16086), .MA34(n16085), .MA33(n16084), .MA32(n16083), 
           .MA31(n16082), .MA30(n16081), .MA29(n16080), .MA28(n16079), 
           .MA27(n16078), .MA26(n16077), .MA25(n16076), .MA24(n16075), 
           .MA23(n16074), .MA22(n16073), .MA21(n16072), .MA20(n16071), 
           .MA19(n16070), .MA18(n16069), .MA17(n16068), .MA16(n16067), 
           .MA15(n16066), .MA14(n16065), .MA13(n16064), .MA12(n16063), 
           .MA11(n16062), .MA10(n16061), .MA9(n16060), .MA8(n16059), 
           .MA7(n16058), .MA6(n16057), .MA5(n16056), .MA4(n16055), .MA3(n16054), 
           .MA2(n16053), .MA1(n16052), .MA0(n16051), .MB35(n16159), 
           .MB34(n16158), .MB33(n16157), .MB32(n16156), .MB31(n16155), 
           .MB30(n16154), .MB29(n16153), .MB28(n16152), .MB27(n16151), 
           .MB26(n16150), .MB25(n16149), .MB24(n16148), .MB23(n16147), 
           .MB22(n16146), .MB21(n16145), .MB20(n16144), .MB19(n16143), 
           .MB18(n16142), .MB17(n16141), .MB16(n16140), .MB15(n16139), 
           .MB14(n16138), .MB13(n16137), .MB12(n16136), .MB11(n16135), 
           .MB10(n16134), .MB9(n16133), .MB8(n16132), .MB7(n16131), 
           .MB6(n16130), .MB5(n16129), .MB4(n16128), .MB3(n16127), .MB2(n16126), 
           .MB1(n16125), .MB0(n16124), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n16341), 
           .R52(n16340), .R51(n16339), .R50(n16338), .R49(n16337), .R48(n16336), 
           .R47(n16335), .R46(n16334), .R45(n16333), .R44(n16332), .R43(n16331), 
           .R42(n16330), .R41(n16329), .R40(n16328), .R39(n16327), .R38(n16326), 
           .R37(n16325), .R36(n16324), .R35(n16323), .R34(n16322), .R33(n16321), 
           .R32(n16320), .R31(n16319), .R30(n16318), .R29(n16317), .R28(n16316), 
           .R27(n16315), .R26(n16314), .R25(n16313), .R24(n16312), .R23(n16311), 
           .R22(n16310), .R21(n16309), .R20(n16308), .R19(n16307), .R18(n16306), 
           .R17(\op_r_23__N_1268[17] ), .R16(\op_r_23__N_1268[16] ), .R15(\op_r_23__N_1268[15] ), 
           .R14(\op_r_23__N_1268[14] ), .R13(\op_r_23__N_1268[13] ), .R12(\op_r_23__N_1268[12] ), 
           .R11(\op_r_23__N_1268[11] ), .R10(\op_r_23__N_1268[10] ), .R9(\op_r_23__N_1268[9] ), 
           .R8(\op_r_23__N_1268[8] ), .R7(\op_r_23__N_1268[7] ), .R6(\op_r_23__N_1268[6] ), 
           .R5(\op_r_23__N_1268[5] ), .R4(\op_r_23__N_1268[4] ), .R3(\op_r_23__N_1268[3] ), 
           .R2(\op_r_23__N_1268[2] ), .R1(\op_r_23__N_1268[1] ), .R0(\op_r_23__N_1268[0] ), 
           .SIGNEDR(n16342));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_43.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_43.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_43.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_43.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_43.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_43.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_43.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_43.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_43.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_43.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_43.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_43.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_43.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_43.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_43.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_43.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_43.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_43.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_43.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_43.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_43.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_43.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_43.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_43.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_43.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_43.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_43.REG_FLAG_CLK = "NONE";
    defparam lat_alu_43.REG_FLAG_CE = "CE0";
    defparam lat_alu_43.REG_FLAG_RST = "RST0";
    defparam lat_alu_43.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_43.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_43.MASK01 = "0x00000000000000";
    defparam lat_alu_43.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_43.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_43.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_43.CLK0_DIV = "ENABLED";
    defparam lat_alu_43.CLK1_DIV = "ENABLED";
    defparam lat_alu_43.CLK2_DIV = "ENABLED";
    defparam lat_alu_43.CLK3_DIV = "ENABLED";
    defparam lat_alu_43.MCPAT = "0x00000000000000";
    defparam lat_alu_43.MASKPAT = "0x00000000000000";
    defparam lat_alu_43.RNDPAT = "0x00000000000000";
    defparam lat_alu_43.GSR = "DISABLED";
    defparam lat_alu_43.RESETMODE = "SYNC";
    defparam lat_alu_43.MULT9_MODE = "DISABLED";
    defparam lat_alu_43.LEGACY = "DISABLED";
    ALU54B lat_alu_44 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n16196), .SIGNEDIB(n16269), .SIGNEDCIN(n16342), .A35(n16195), 
           .A34(n16194), .A33(n16193), .A32(n16192), .A31(n16191), .A30(n16190), 
           .A29(n16189), .A28(n16188), .A27(n16187), .A26(n16186), .A25(n16185), 
           .A24(n16184), .A23(n16183), .A22(n16182), .A21(n16181), .A20(n16180), 
           .A19(n16179), .A18(n16178), .A17(n16177), .A16(n16176), .A15(n16175), 
           .A14(n16174), .A13(n16173), .A12(n16172), .A11(n16171), .A10(n16170), 
           .A9(n16169), .A8(n16168), .A7(n16167), .A6(n16166), .A5(n16165), 
           .A4(n16164), .A3(n16163), .A2(n16162), .A1(n16161), .A0(n16160), 
           .B35(n16268), .B34(n16267), .B33(n16266), .B32(n16265), .B31(n16264), 
           .B30(n16263), .B29(n16262), .B28(n16261), .B27(n16260), .B26(n16259), 
           .B25(n16258), .B24(n16257), .B23(n16256), .B22(n16255), .B21(n16254), 
           .B20(n16253), .B19(n16252), .B18(n16251), .B17(n16250), .B16(n16249), 
           .B15(n16248), .B14(n16247), .B13(n16246), .B12(n16245), .B11(n16244), 
           .B10(n16243), .B9(n16242), .B8(n16241), .B7(n16240), .B6(n16239), 
           .B5(n16238), .B4(n16237), .B3(n16236), .B2(n16235), .B1(n16234), 
           .B0(n16233), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n16232), .MA34(n16231), .MA33(n16230), .MA32(n16229), 
           .MA31(n16228), .MA30(n16227), .MA29(n16226), .MA28(n16225), 
           .MA27(n16224), .MA26(n16223), .MA25(n16222), .MA24(n16221), 
           .MA23(n16220), .MA22(n16219), .MA21(n16218), .MA20(n16217), 
           .MA19(n16216), .MA18(n16215), .MA17(n16214), .MA16(n16213), 
           .MA15(n16212), .MA14(n16211), .MA13(n16210), .MA12(n16209), 
           .MA11(n16208), .MA10(n16207), .MA9(n16206), .MA8(n16205), 
           .MA7(n16204), .MA6(n16203), .MA5(n16202), .MA4(n16201), .MA3(n16200), 
           .MA2(n16199), .MA1(n16198), .MA0(n16197), .MB35(n16305), 
           .MB34(n16304), .MB33(n16303), .MB32(n16302), .MB31(n16301), 
           .MB30(n16300), .MB29(n16299), .MB28(n16298), .MB27(n16297), 
           .MB26(n16296), .MB25(n16295), .MB24(n16294), .MB23(n16293), 
           .MB22(n16292), .MB21(n16291), .MB20(n16290), .MB19(n16289), 
           .MB18(n16288), .MB17(n16287), .MB16(n16286), .MB15(n16285), 
           .MB14(n16284), .MB13(n16283), .MB12(n16282), .MB11(n16281), 
           .MB10(n16280), .MB9(n16279), .MB8(n16278), .MB7(n16277), 
           .MB6(n16276), .MB5(n16275), .MB4(n16274), .MB3(n16273), .MB2(n16272), 
           .MB1(n16271), .MB0(n16270), .CIN53(n16341), .CIN52(n16340), 
           .CIN51(n16339), .CIN50(n16338), .CIN49(n16337), .CIN48(n16336), 
           .CIN47(n16335), .CIN46(n16334), .CIN45(n16333), .CIN44(n16332), 
           .CIN43(n16331), .CIN42(n16330), .CIN41(n16329), .CIN40(n16328), 
           .CIN39(n16327), .CIN38(n16326), .CIN37(n16325), .CIN36(n16324), 
           .CIN35(n16323), .CIN34(n16322), .CIN33(n16321), .CIN32(n16320), 
           .CIN31(n16319), .CIN30(n16318), .CIN29(n16317), .CIN28(n16316), 
           .CIN27(n16315), .CIN26(n16314), .CIN25(n16313), .CIN24(n16312), 
           .CIN23(n16311), .CIN22(n16310), .CIN21(n16309), .CIN20(n16308), 
           .CIN19(n16307), .CIN18(n16306), .CIN17(\op_r_23__N_1268[17] ), 
           .CIN16(\op_r_23__N_1268[16] ), .CIN15(\op_r_23__N_1268[15] ), 
           .CIN14(\op_r_23__N_1268[14] ), .CIN13(\op_r_23__N_1268[13] ), 
           .CIN12(\op_r_23__N_1268[12] ), .CIN11(\op_r_23__N_1268[11] ), 
           .CIN10(\op_r_23__N_1268[10] ), .CIN9(\op_r_23__N_1268[9] ), .CIN8(\op_r_23__N_1268[8] ), 
           .CIN7(\op_r_23__N_1268[7] ), .CIN6(\op_r_23__N_1268[6] ), .CIN5(\op_r_23__N_1268[5] ), 
           .CIN4(\op_r_23__N_1268[4] ), .CIN3(\op_r_23__N_1268[3] ), .CIN2(\op_r_23__N_1268[2] ), 
           .CIN1(\op_r_23__N_1268[1] ), .CIN0(\op_r_23__N_1268[0] ), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(\op_r_23__N_1268[31] ), 
           .R12(\op_r_23__N_1268[30] ), .R11(\op_r_23__N_1268[29] ), .R10(\op_r_23__N_1268[28] ), 
           .R9(\op_r_23__N_1268[27] ), .R8(\op_r_23__N_1268[26] ), .R7(\op_r_23__N_1268[25] ), 
           .R6(\op_r_23__N_1268[24] ), .R5(\op_r_23__N_1268[23] ), .R4(\op_r_23__N_1268[22] ), 
           .R3(\op_r_23__N_1268[21] ), .R2(\op_r_23__N_1268[20] ), .R1(\op_r_23__N_1268[19] ), 
           .R0(\op_r_23__N_1268[18] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_alu_44.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_44.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_44.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_44.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_44.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_44.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_44.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_44.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_44.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_44.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_44.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_44.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_44.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_44.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_44.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_44.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_44.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_44.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_44.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_44.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_44.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_44.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_44.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_44.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_44.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_44.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_44.REG_FLAG_CLK = "NONE";
    defparam lat_alu_44.REG_FLAG_CE = "CE0";
    defparam lat_alu_44.REG_FLAG_RST = "RST0";
    defparam lat_alu_44.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_44.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_44.MASK01 = "0x00000000000000";
    defparam lat_alu_44.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_44.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_44.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_44.CLK0_DIV = "ENABLED";
    defparam lat_alu_44.CLK1_DIV = "ENABLED";
    defparam lat_alu_44.CLK2_DIV = "ENABLED";
    defparam lat_alu_44.CLK3_DIV = "ENABLED";
    defparam lat_alu_44.MCPAT = "0x00000000000000";
    defparam lat_alu_44.MASKPAT = "0x00000000000000";
    defparam lat_alu_44.RNDPAT = "0x00000000000000";
    defparam lat_alu_44.GSR = "DISABLED";
    defparam lat_alu_44.RESETMODE = "SYNC";
    defparam lat_alu_44.MULT9_MODE = "DISABLED";
    defparam lat_alu_44.LEGACY = "DISABLED";
    ALU54B lat_alu_24 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n14812), .SIGNEDIB(n14885), .SIGNEDCIN(n14958), .A35(n14811), 
           .A34(n14810), .A33(n14809), .A32(n14808), .A31(n14807), .A30(n14806), 
           .A29(n14805), .A28(n14804), .A27(n14803), .A26(n14802), .A25(n14801), 
           .A24(n14800), .A23(n14799), .A22(n14798), .A21(n14797), .A20(n14796), 
           .A19(n14795), .A18(n14794), .A17(n14793), .A16(n14792), .A15(n14791), 
           .A14(n14790), .A13(n14789), .A12(n14788), .A11(n14787), .A10(n14786), 
           .A9(n14785), .A8(n14784), .A7(n14783), .A6(n14782), .A5(n14781), 
           .A4(n14780), .A3(n14779), .A2(n14778), .A1(n14777), .A0(n14776), 
           .B35(n14884), .B34(n14883), .B33(n14882), .B32(n14881), .B31(n14880), 
           .B30(n14879), .B29(n14878), .B28(n14877), .B27(n14876), .B26(n14875), 
           .B25(n14874), .B24(n14873), .B23(n14872), .B22(n14871), .B21(n14870), 
           .B20(n14869), .B19(n14868), .B18(n14867), .B17(n14866), .B16(n14865), 
           .B15(n14864), .B14(n14863), .B13(n14862), .B12(n14861), .B11(n14860), 
           .B10(n14859), .B9(n14858), .B8(n14857), .B7(n14856), .B6(n14855), 
           .B5(n14854), .B4(n14853), .B3(n14852), .B2(n14851), .B1(n14850), 
           .B0(n14849), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n14848), .MA34(n14847), .MA33(n14846), .MA32(n14845), 
           .MA31(n14844), .MA30(n14843), .MA29(n14842), .MA28(n14841), 
           .MA27(n14840), .MA26(n14839), .MA25(n14838), .MA24(n14837), 
           .MA23(n14836), .MA22(n14835), .MA21(n14834), .MA20(n14833), 
           .MA19(n14832), .MA18(n14831), .MA17(n14830), .MA16(n14829), 
           .MA15(n14828), .MA14(n14827), .MA13(n14826), .MA12(n14825), 
           .MA11(n14824), .MA10(n14823), .MA9(n14822), .MA8(n14821), 
           .MA7(n14820), .MA6(n14819), .MA5(n14818), .MA4(n14817), .MA3(n14816), 
           .MA2(n14815), .MA1(n14814), .MA0(n14813), .MB35(n14921), 
           .MB34(n14920), .MB33(n14919), .MB32(n14918), .MB31(n14917), 
           .MB30(n14916), .MB29(n14915), .MB28(n14914), .MB27(n14913), 
           .MB26(n14912), .MB25(n14911), .MB24(n14910), .MB23(n14909), 
           .MB22(n14908), .MB21(n14907), .MB20(n14906), .MB19(n14905), 
           .MB18(n14904), .MB17(n14903), .MB16(n14902), .MB15(n14901), 
           .MB14(n14900), .MB13(n14899), .MB12(n14898), .MB11(n14897), 
           .MB10(n14896), .MB9(n14895), .MB8(n14894), .MB7(n14893), 
           .MB6(n14892), .MB5(n14891), .MB4(n14890), .MB3(n14889), .MB2(n14888), 
           .MB1(n14887), .MB0(n14886), .CIN53(n14957), .CIN52(n14956), 
           .CIN51(n14955), .CIN50(n14954), .CIN49(n14953), .CIN48(n14952), 
           .CIN47(n14951), .CIN46(n14950), .CIN45(n14949), .CIN44(n14948), 
           .CIN43(n14947), .CIN42(n14946), .CIN41(n14945), .CIN40(n14944), 
           .CIN39(n14943), .CIN38(n14942), .CIN37(n14941), .CIN36(n14940), 
           .CIN35(n14939), .CIN34(n14938), .CIN33(n14937), .CIN32(n14936), 
           .CIN31(n14935), .CIN30(n14934), .CIN29(n14933), .CIN28(n14932), 
           .CIN27(n14931), .CIN26(n14930), .CIN25(n14929), .CIN24(n14928), 
           .CIN23(n14927), .CIN22(n14926), .CIN21(n14925), .CIN20(n14924), 
           .CIN19(n14923), .CIN18(n14922), .CIN17(n9088), .CIN16(n9089), 
           .CIN15(n9090), .CIN14(n9091), .CIN13(n9092), .CIN12(n9093), 
           .CIN11(n9094), .CIN10(n9095), .CIN9(n9096), .CIN8(n9097), 
           .CIN7(n9098), .CIN6(n9099), .CIN5(n9100), .CIN4(n9101), .CIN3(n9102), 
           .CIN2(n9103), .CIN1(n9104), .CIN0(n9105), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R7(n9080), .R6(n9081), .R5(n9082), 
           .R4(n9083), .R3(n9084), .R2(n9085), .R1(n9086), .R0(n9087));
    defparam lat_alu_24.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_24.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_24.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_24.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_24.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_24.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_24.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_24.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_24.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_24.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_24.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_24.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_24.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_24.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_24.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_24.REG_FLAG_CLK = "NONE";
    defparam lat_alu_24.REG_FLAG_CE = "CE0";
    defparam lat_alu_24.REG_FLAG_RST = "RST0";
    defparam lat_alu_24.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_24.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_24.MASK01 = "0x00000000000000";
    defparam lat_alu_24.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_24.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_24.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_24.CLK0_DIV = "ENABLED";
    defparam lat_alu_24.CLK1_DIV = "ENABLED";
    defparam lat_alu_24.CLK2_DIV = "ENABLED";
    defparam lat_alu_24.CLK3_DIV = "ENABLED";
    defparam lat_alu_24.MCPAT = "0x00000000000000";
    defparam lat_alu_24.MASKPAT = "0x00000000000000";
    defparam lat_alu_24.RNDPAT = "0x00000000000000";
    defparam lat_alu_24.GSR = "DISABLED";
    defparam lat_alu_24.RESETMODE = "SYNC";
    defparam lat_alu_24.MULT9_MODE = "DISABLED";
    defparam lat_alu_24.LEGACY = "DISABLED";
    ALU54B lat_alu_23 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n14666), .SIGNEDIB(n14739), .SIGNEDCIN(GND_net), 
           .A35(n14665), .A34(n14664), .A33(n14663), .A32(n14662), .A31(n14661), 
           .A30(n14660), .A29(n14659), .A28(n14658), .A27(n14657), .A26(n14656), 
           .A25(n14655), .A24(n14654), .A23(n14653), .A22(n14652), .A21(n14651), 
           .A20(n14650), .A19(n14649), .A18(n14648), .A17(n14647), .A16(n14646), 
           .A15(n14645), .A14(n14644), .A13(n14643), .A12(n14642), .A11(n14641), 
           .A10(n14640), .A9(n14639), .A8(n14638), .A7(n14637), .A6(n14636), 
           .A5(n14635), .A4(n14634), .A3(n14633), .A2(n14632), .A1(n14631), 
           .A0(n14630), .B35(n14738), .B34(n14737), .B33(n14736), .B32(n14735), 
           .B31(n14734), .B30(n14733), .B29(n14732), .B28(n14731), .B27(n14730), 
           .B26(n14729), .B25(n14728), .B24(n14727), .B23(n14726), .B22(n14725), 
           .B21(n14724), .B20(n14723), .B19(n14722), .B18(n14721), .B17(n14720), 
           .B16(n14719), .B15(n14718), .B14(n14717), .B13(n14716), .B12(n14715), 
           .B11(n14714), .B10(n14713), .B9(n14712), .B8(n14711), .B7(n14710), 
           .B6(n14709), .B5(n14708), .B4(n14707), .B3(n14706), .B2(n14705), 
           .B1(n14704), .B0(n14703), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n14702), .MA34(n14701), .MA33(n14700), .MA32(n14699), 
           .MA31(n14698), .MA30(n14697), .MA29(n14696), .MA28(n14695), 
           .MA27(n14694), .MA26(n14693), .MA25(n14692), .MA24(n14691), 
           .MA23(n14690), .MA22(n14689), .MA21(n14688), .MA20(n14687), 
           .MA19(n14686), .MA18(n14685), .MA17(n14684), .MA16(n14683), 
           .MA15(n14682), .MA14(n14681), .MA13(n14680), .MA12(n14679), 
           .MA11(n14678), .MA10(n14677), .MA9(n14676), .MA8(n14675), 
           .MA7(n14674), .MA6(n14673), .MA5(n14672), .MA4(n14671), .MA3(n14670), 
           .MA2(n14669), .MA1(n14668), .MA0(n14667), .MB35(n14775), 
           .MB34(n14774), .MB33(n14773), .MB32(n14772), .MB31(n14771), 
           .MB30(n14770), .MB29(n14769), .MB28(n14768), .MB27(n14767), 
           .MB26(n14766), .MB25(n14765), .MB24(n14764), .MB23(n14763), 
           .MB22(n14762), .MB21(n14761), .MB20(n14760), .MB19(n14759), 
           .MB18(n14758), .MB17(n14757), .MB16(n14756), .MB15(n14755), 
           .MB14(n14754), .MB13(n14753), .MB12(n14752), .MB11(n14751), 
           .MB10(n14750), .MB9(n14749), .MB8(n14748), .MB7(n14747), 
           .MB6(n14746), .MB5(n14745), .MB4(n14744), .MB3(n14743), .MB2(n14742), 
           .MB1(n14741), .MB0(n14740), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n14957), 
           .R52(n14956), .R51(n14955), .R50(n14954), .R49(n14953), .R48(n14952), 
           .R47(n14951), .R46(n14950), .R45(n14949), .R44(n14948), .R43(n14947), 
           .R42(n14946), .R41(n14945), .R40(n14944), .R39(n14943), .R38(n14942), 
           .R37(n14941), .R36(n14940), .R35(n14939), .R34(n14938), .R33(n14937), 
           .R32(n14936), .R31(n14935), .R30(n14934), .R29(n14933), .R28(n14932), 
           .R27(n14931), .R26(n14930), .R25(n14929), .R24(n14928), .R23(n14927), 
           .R22(n14926), .R21(n14925), .R20(n14924), .R19(n14923), .R18(n14922), 
           .R17(n9088), .R16(n9089), .R15(n9090), .R14(n9091), .R13(n9092), 
           .R12(n9093), .R11(n9094), .R10(n9095), .R9(n9096), .R8(n9097), 
           .R7(n9098), .R6(n9099), .R5(n9100), .R4(n9101), .R3(n9102), 
           .R2(n9103), .R1(n9104), .R0(n9105), .SIGNEDR(n14958));
    defparam lat_alu_23.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_23.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_23.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_23.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_23.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_23.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_23.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_23.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_23.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_23.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_23.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_23.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_23.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_23.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_23.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_23.REG_FLAG_CLK = "NONE";
    defparam lat_alu_23.REG_FLAG_CE = "CE0";
    defparam lat_alu_23.REG_FLAG_RST = "RST0";
    defparam lat_alu_23.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_23.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_23.MASK01 = "0x00000000000000";
    defparam lat_alu_23.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_23.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_23.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_23.CLK0_DIV = "ENABLED";
    defparam lat_alu_23.CLK1_DIV = "ENABLED";
    defparam lat_alu_23.CLK2_DIV = "ENABLED";
    defparam lat_alu_23.CLK3_DIV = "ENABLED";
    defparam lat_alu_23.MCPAT = "0x00000000000000";
    defparam lat_alu_23.MASKPAT = "0x00000000000000";
    defparam lat_alu_23.RNDPAT = "0x00000000000000";
    defparam lat_alu_23.GSR = "DISABLED";
    defparam lat_alu_23.RESETMODE = "SYNC";
    defparam lat_alu_23.MULT9_MODE = "DISABLED";
    defparam lat_alu_23.LEGACY = "DISABLED";
    MULT18X18D lat_mult_22 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n319), .B16(n319), 
            .B15(n319), .B14(n319), .B13(n319), .B12(n319), .B11(n319), 
            .B10(n319), .B9(n319), .B8(n319), .B7(n319), .B6(n319), 
            .B5(n319), .B4(n319), .B3(n319), .B2(n319), .B1(n319), 
            .B0(n319), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14866), 
            .ROA16(n14865), .ROA15(n14864), .ROA14(n14863), .ROA13(n14862), 
            .ROA12(n14861), .ROA11(n14860), .ROA10(n14859), .ROA9(n14858), 
            .ROA8(n14857), .ROA7(n14856), .ROA6(n14855), .ROA5(n14854), 
            .ROA4(n14853), .ROA3(n14852), .ROA2(n14851), .ROA1(n14850), 
            .ROA0(n14849), .ROB17(n14884), .ROB16(n14883), .ROB15(n14882), 
            .ROB14(n14881), .ROB13(n14880), .ROB12(n14879), .ROB11(n14878), 
            .ROB10(n14877), .ROB9(n14876), .ROB8(n14875), .ROB7(n14874), 
            .ROB6(n14873), .ROB5(n14872), .ROB4(n14871), .ROB3(n14870), 
            .ROB2(n14869), .ROB1(n14868), .ROB0(n14867), .P35(n14921), 
            .P34(n14920), .P33(n14919), .P32(n14918), .P31(n14917), 
            .P30(n14916), .P29(n14915), .P28(n14914), .P27(n14913), 
            .P26(n14912), .P25(n14911), .P24(n14910), .P23(n14909), 
            .P22(n14908), .P21(n14907), .P20(n14906), .P19(n14905), 
            .P18(n14904), .P17(n14903), .P16(n14902), .P15(n14901), 
            .P14(n14900), .P13(n14899), .P12(n14898), .P11(n14897), 
            .P10(n14896), .P9(n14895), .P8(n14894), .P7(n14893), .P6(n14892), 
            .P5(n14891), .P4(n14890), .P3(n14889), .P2(n14888), .P1(n14887), 
            .P0(n14886), .SIGNEDP(n14885));
    defparam lat_mult_22.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_22.REG_INPUTA_CE = "CE0";
    defparam lat_mult_22.REG_INPUTA_RST = "RST0";
    defparam lat_mult_22.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_22.REG_INPUTB_CE = "CE0";
    defparam lat_mult_22.REG_INPUTB_RST = "RST0";
    defparam lat_mult_22.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_22.REG_INPUTC_CE = "CE0";
    defparam lat_mult_22.REG_INPUTC_RST = "RST0";
    defparam lat_mult_22.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_22.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_22.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_22.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_22.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_22.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_22.CLK0_DIV = "ENABLED";
    defparam lat_mult_22.CLK1_DIV = "ENABLED";
    defparam lat_mult_22.CLK2_DIV = "ENABLED";
    defparam lat_mult_22.CLK3_DIV = "ENABLED";
    defparam lat_mult_22.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_22.GSR = "DISABLED";
    defparam lat_mult_22.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_22.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_22.MULT_BYPASS = "DISABLED";
    defparam lat_mult_22.RESETMODE = "SYNC";
    MULT18X18D lat_mult_21 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n319), .B16(n319), 
            .B15(n319), .B14(n319), .B13(n319), .B12(n319), .B11(n319), 
            .B10(n319), .B9(n319), .B8(n319), .B7(n319), .B6(n319), 
            .B5(n319), .B4(n319), .B3(n319), .B2(n319), .B1(n319), 
            .B0(n319), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n14793), 
            .ROA16(n14792), .ROA15(n14791), .ROA14(n14790), .ROA13(n14789), 
            .ROA12(n14788), .ROA11(n14787), .ROA10(n14786), .ROA9(n14785), 
            .ROA8(n14784), .ROA7(n14783), .ROA6(n14782), .ROA5(n14781), 
            .ROA4(n14780), .ROA3(n14779), .ROA2(n14778), .ROA1(n14777), 
            .ROA0(n14776), .ROB17(n14811), .ROB16(n14810), .ROB15(n14809), 
            .ROB14(n14808), .ROB13(n14807), .ROB12(n14806), .ROB11(n14805), 
            .ROB10(n14804), .ROB9(n14803), .ROB8(n14802), .ROB7(n14801), 
            .ROB6(n14800), .ROB5(n14799), .ROB4(n14798), .ROB3(n14797), 
            .ROB2(n14796), .ROB1(n14795), .ROB0(n14794), .P35(n14848), 
            .P34(n14847), .P33(n14846), .P32(n14845), .P31(n14844), 
            .P30(n14843), .P29(n14842), .P28(n14841), .P27(n14840), 
            .P26(n14839), .P25(n14838), .P24(n14837), .P23(n14836), 
            .P22(n14835), .P21(n14834), .P20(n14833), .P19(n14832), 
            .P18(n14831), .P17(n14830), .P16(n14829), .P15(n14828), 
            .P14(n14827), .P13(n14826), .P12(n14825), .P11(n14824), 
            .P10(n14823), .P9(n14822), .P8(n14821), .P7(n14820), .P6(n14819), 
            .P5(n14818), .P4(n14817), .P3(n14816), .P2(n14815), .P1(n14814), 
            .P0(n14813), .SIGNEDP(n14812));
    defparam lat_mult_21.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_21.REG_INPUTA_CE = "CE0";
    defparam lat_mult_21.REG_INPUTA_RST = "RST0";
    defparam lat_mult_21.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_21.REG_INPUTB_CE = "CE0";
    defparam lat_mult_21.REG_INPUTB_RST = "RST0";
    defparam lat_mult_21.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_21.REG_INPUTC_CE = "CE0";
    defparam lat_mult_21.REG_INPUTC_RST = "RST0";
    defparam lat_mult_21.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_21.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_21.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_21.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_21.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_21.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_21.CLK0_DIV = "ENABLED";
    defparam lat_mult_21.CLK1_DIV = "ENABLED";
    defparam lat_mult_21.CLK2_DIV = "ENABLED";
    defparam lat_mult_21.CLK3_DIV = "ENABLED";
    defparam lat_mult_21.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_21.GSR = "DISABLED";
    defparam lat_mult_21.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_21.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_21.MULT_BYPASS = "DISABLED";
    defparam lat_mult_21.RESETMODE = "SYNC";
    MULT18X18D lat_mult_20 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n11579), 
            .B16(n11578), .B15(n11577), .B14(n11576), .B13(n11575), 
            .B12(n11574), .B11(n11573), .B10(n11572), .B9(n11571), .B8(n11570), 
            .B7(n11569), .B6(n11568), .B5(n11567), .B4(n11566), .B3(n11565), 
            .B2(n11564), .B1(n11563), .B0(n11562), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n14720), .ROA16(n14719), .ROA15(n14718), .ROA14(n14717), 
            .ROA13(n14716), .ROA12(n14715), .ROA11(n14714), .ROA10(n14713), 
            .ROA9(n14712), .ROA8(n14711), .ROA7(n14710), .ROA6(n14709), 
            .ROA5(n14708), .ROA4(n14707), .ROA3(n14706), .ROA2(n14705), 
            .ROA1(n14704), .ROA0(n14703), .ROB17(n14738), .ROB16(n14737), 
            .ROB15(n14736), .ROB14(n14735), .ROB13(n14734), .ROB12(n14733), 
            .ROB11(n14732), .ROB10(n14731), .ROB9(n14730), .ROB8(n14729), 
            .ROB7(n14728), .ROB6(n14727), .ROB5(n14726), .ROB4(n14725), 
            .ROB3(n14724), .ROB2(n14723), .ROB1(n14722), .ROB0(n14721), 
            .P35(n14775), .P34(n14774), .P33(n14773), .P32(n14772), 
            .P31(n14771), .P30(n14770), .P29(n14769), .P28(n14768), 
            .P27(n14767), .P26(n14766), .P25(n14765), .P24(n14764), 
            .P23(n14763), .P22(n14762), .P21(n14761), .P20(n14760), 
            .P19(n14759), .P18(n14758), .P17(n14757), .P16(n14756), 
            .P15(n14755), .P14(n14754), .P13(n14753), .P12(n14752), 
            .P11(n14751), .P10(n14750), .P9(n14749), .P8(n14748), .P7(n14747), 
            .P6(n14746), .P5(n14745), .P4(n14744), .P3(n14743), .P2(n14742), 
            .P1(n14741), .P0(n14740), .SIGNEDP(n14739));
    defparam lat_mult_20.REG_INPUTA_CLK = "NONE";
    defparam lat_mult_20.REG_INPUTA_CE = "CE0";
    defparam lat_mult_20.REG_INPUTA_RST = "RST0";
    defparam lat_mult_20.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_20.REG_INPUTB_CE = "CE0";
    defparam lat_mult_20.REG_INPUTB_RST = "RST0";
    defparam lat_mult_20.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_20.REG_INPUTC_CE = "CE0";
    defparam lat_mult_20.REG_INPUTC_RST = "RST0";
    defparam lat_mult_20.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_20.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_20.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_20.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_20.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_20.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_20.CLK0_DIV = "ENABLED";
    defparam lat_mult_20.CLK1_DIV = "ENABLED";
    defparam lat_mult_20.CLK2_DIV = "ENABLED";
    defparam lat_mult_20.CLK3_DIV = "ENABLED";
    defparam lat_mult_20.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_20.GSR = "DISABLED";
    defparam lat_mult_20.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_20.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_20.MULT_BYPASS = "DISABLED";
    defparam lat_mult_20.RESETMODE = "SYNC";
    MULT18X18D mult_978 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(n11579), 
            .B16(n11578), .B15(n11577), .B14(n11576), .B13(n11575), 
            .B12(n11574), .B11(n11573), .B10(n11572), .B9(n11571), .B8(n11570), 
            .B7(n11569), .B6(n11568), .B5(n11567), .B4(n11566), .B3(n11565), 
            .B2(n11564), .B1(n11563), .B0(n11562), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n14647), .ROA16(n14646), .ROA15(n14645), .ROA14(n14644), 
            .ROA13(n14643), .ROA12(n14642), .ROA11(n14641), .ROA10(n14640), 
            .ROA9(n14639), .ROA8(n14638), .ROA7(n14637), .ROA6(n14636), 
            .ROA5(n14635), .ROA4(n14634), .ROA3(n14633), .ROA2(n14632), 
            .ROA1(n14631), .ROA0(n14630), .ROB17(n14665), .ROB16(n14664), 
            .ROB15(n14663), .ROB14(n14662), .ROB13(n14661), .ROB12(n14660), 
            .ROB11(n14659), .ROB10(n14658), .ROB9(n14657), .ROB8(n14656), 
            .ROB7(n14655), .ROB6(n14654), .ROB5(n14653), .ROB4(n14652), 
            .ROB3(n14651), .ROB2(n14650), .ROB1(n14649), .ROB0(n14648), 
            .P35(n14702), .P34(n14701), .P33(n14700), .P32(n14699), 
            .P31(n14698), .P30(n14697), .P29(n14696), .P28(n14695), 
            .P27(n14694), .P26(n14693), .P25(n14692), .P24(n14691), 
            .P23(n14690), .P22(n14689), .P21(n14688), .P20(n14687), 
            .P19(n14686), .P18(n14685), .P17(n14684), .P16(n14683), 
            .P15(n14682), .P14(n14681), .P13(n14680), .P12(n14679), 
            .P11(n14678), .P10(n14677), .P9(n14676), .P8(n14675), .P7(n14674), 
            .P6(n14673), .P5(n14672), .P4(n14671), .P3(n14670), .P2(n14669), 
            .P1(n14668), .P0(n14667), .SIGNEDP(n14666));
    defparam mult_978.REG_INPUTA_CLK = "NONE";
    defparam mult_978.REG_INPUTA_CE = "CE0";
    defparam mult_978.REG_INPUTA_RST = "RST0";
    defparam mult_978.REG_INPUTB_CLK = "NONE";
    defparam mult_978.REG_INPUTB_CE = "CE0";
    defparam mult_978.REG_INPUTB_RST = "RST0";
    defparam mult_978.REG_INPUTC_CLK = "NONE";
    defparam mult_978.REG_INPUTC_CE = "CE0";
    defparam mult_978.REG_INPUTC_RST = "RST0";
    defparam mult_978.REG_PIPELINE_CLK = "NONE";
    defparam mult_978.REG_PIPELINE_CE = "CE0";
    defparam mult_978.REG_PIPELINE_RST = "RST0";
    defparam mult_978.REG_OUTPUT_CLK = "NONE";
    defparam mult_978.REG_OUTPUT_CE = "CE0";
    defparam mult_978.REG_OUTPUT_RST = "RST0";
    defparam mult_978.CLK0_DIV = "ENABLED";
    defparam mult_978.CLK1_DIV = "ENABLED";
    defparam mult_978.CLK2_DIV = "ENABLED";
    defparam mult_978.CLK3_DIV = "ENABLED";
    defparam mult_978.HIGHSPEED_CLK = "NONE";
    defparam mult_978.GSR = "DISABLED";
    defparam mult_978.CAS_MATCH_REG = "FALSE";
    defparam mult_978.SOURCEB_MODE = "B_SHIFT";
    defparam mult_978.MULT_BYPASS = "DISABLED";
    defparam mult_978.RESETMODE = "SYNC";
    LUT4 i12683_4_lut (.A(n34843), .B(delay_i_23__N_1202[0]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[0]), .Z(dout_i_23__N_5974[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12683_4_lut.init = 16'hcac0;
    LUT4 i13058_4_lut (.A(n34843), .B(delay_i_23__N_1202[1]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[1]), .Z(dout_i_23__N_5974[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13058_4_lut.init = 16'hcac0;
    LUT4 i13060_4_lut (.A(n34843), .B(delay_i_23__N_1202[2]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[2]), .Z(dout_i_23__N_5974[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13060_4_lut.init = 16'hcac0;
    LUT4 i13062_4_lut (.A(n34843), .B(delay_i_23__N_1202[3]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[3]), .Z(dout_i_23__N_5974[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13062_4_lut.init = 16'hcac0;
    LUT4 i13064_4_lut (.A(n34843), .B(delay_i_23__N_1202[4]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[4]), .Z(dout_i_23__N_5974[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13064_4_lut.init = 16'hcac0;
    LUT4 i13066_4_lut (.A(n34843), .B(delay_i_23__N_1202[5]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[5]), .Z(dout_i_23__N_5974[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13066_4_lut.init = 16'hcac0;
    LUT4 i13068_4_lut (.A(n34843), .B(delay_i_23__N_1202[6]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[6]), .Z(dout_i_23__N_5974[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13068_4_lut.init = 16'hcac0;
    LUT4 i13070_4_lut (.A(n34843), .B(delay_i_23__N_1202[7]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[7]), .Z(dout_i_23__N_5974[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13070_4_lut.init = 16'hcac0;
    LUT4 i13072_4_lut (.A(n34843), .B(delay_i_23__N_1202[8]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[8]), .Z(dout_i_23__N_5974[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13072_4_lut.init = 16'hcac0;
    LUT4 i13074_4_lut (.A(n34843), .B(delay_i_23__N_1202[9]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[9]), .Z(dout_i_23__N_5974[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13074_4_lut.init = 16'hcac0;
    LUT4 i13076_4_lut (.A(n34843), .B(delay_i_23__N_1202[10]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[10]), .Z(dout_i_23__N_5974[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13076_4_lut.init = 16'hcac0;
    LUT4 i13078_4_lut (.A(n34843), .B(delay_i_23__N_1202[11]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[11]), .Z(dout_i_23__N_5974[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13078_4_lut.init = 16'hcac0;
    LUT4 i13080_4_lut (.A(n34843), .B(delay_i_23__N_1202[12]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[12]), .Z(dout_i_23__N_5974[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13080_4_lut.init = 16'hcac0;
    LUT4 i13082_4_lut (.A(n34843), .B(delay_i_23__N_1202[13]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[13]), .Z(dout_i_23__N_5974[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13082_4_lut.init = 16'hcac0;
    LUT4 i13084_4_lut (.A(n34843), .B(delay_i_23__N_1202[14]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[14]), .Z(dout_i_23__N_5974[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13084_4_lut.init = 16'hcac0;
    LUT4 i13086_4_lut (.A(n34843), .B(delay_i_23__N_1202[15]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[15]), .Z(dout_i_23__N_5974[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13086_4_lut.init = 16'hcac0;
    LUT4 i13088_4_lut (.A(n34843), .B(delay_i_23__N_1202[16]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[16]), .Z(dout_i_23__N_5974[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13088_4_lut.init = 16'hcac0;
    LUT4 i13090_4_lut (.A(n34843), .B(delay_i_23__N_1202[17]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[17]), .Z(dout_i_23__N_5974[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13090_4_lut.init = 16'hcac0;
    LUT4 i13092_4_lut (.A(n34843), .B(delay_i_23__N_1202[18]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[18]), .Z(dout_i_23__N_5974[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13092_4_lut.init = 16'hcac0;
    LUT4 i13094_4_lut (.A(n34843), .B(delay_i_23__N_1202[19]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[19]), .Z(dout_i_23__N_5974[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13094_4_lut.init = 16'hcac0;
    LUT4 i13096_4_lut (.A(n34843), .B(delay_i_23__N_1202[20]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[20]), .Z(dout_i_23__N_5974[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13096_4_lut.init = 16'hcac0;
    LUT4 i13098_4_lut (.A(n34843), .B(delay_i_23__N_1202[21]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[21]), .Z(dout_i_23__N_5974[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13098_4_lut.init = 16'hcac0;
    LUT4 i13100_4_lut (.A(n34843), .B(delay_i_23__N_1202[22]), .C(\no5_state[0] ), 
         .D(op_i_23__N_1154[22]), .Z(dout_i_23__N_5974[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13100_4_lut.init = 16'hcac0;
    LUT4 i10877_4_lut (.A(op_i_23__N_1154[23]), .B(delay_i_23__N_1202[23]), 
         .C(\no5_state[0] ), .D(n34843), .Z(dout_i_23__N_5974[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i10877_4_lut.init = 16'hcac0;
    MULT18X18D lat_mult_40 (.A17(dout_i_23__N_5974[23]), .A16(dout_i_23__N_5974[23]), 
            .A15(dout_i_23__N_5974[23]), .A14(dout_i_23__N_5974[23]), .A13(dout_i_23__N_5974[23]), 
            .A12(dout_i_23__N_5974[23]), .A11(dout_i_23__N_5974[23]), .A10(dout_i_23__N_5974[23]), 
            .A9(dout_i_23__N_5974[23]), .A8(dout_i_23__N_5974[23]), .A7(dout_i_23__N_5974[23]), 
            .A6(dout_i_23__N_5974[23]), .A5(dout_i_23__N_5974[23]), .A4(dout_i_23__N_5974[22]), 
            .A3(dout_i_23__N_5974[21]), .A2(dout_i_23__N_5974[20]), .A1(dout_i_23__N_5974[19]), 
            .A0(dout_i_23__N_5974[18]), .B17(GND_net), .B16(GND_net), 
            .B15(GND_net), .B14(GND_net), .B13(GND_net), .B12(GND_net), 
            .B11(GND_net), .B10(GND_net), .B9(GND_net), .B8(VCC_net), 
            .B7(GND_net), .B6(GND_net), .B5(GND_net), .B4(GND_net), 
            .B3(GND_net), .B2(GND_net), .B1(GND_net), .B0(GND_net), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(n34738), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(rst_n_N_2), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n16104), .ROA16(n16103), 
            .ROA15(n16102), .ROA14(n16101), .ROA13(n16100), .ROA12(n16099), 
            .ROA11(n16098), .ROA10(n16097), .ROA9(n16096), .ROA8(n16095), 
            .ROA7(n16094), .ROA6(n16093), .ROA5(n16092), .ROA4(n16091), 
            .ROA3(n16090), .ROA2(n16089), .ROA1(n16088), .ROA0(n16087), 
            .ROB17(n16122), .ROB16(n16121), .ROB15(n16120), .ROB14(n16119), 
            .ROB13(n16118), .ROB12(n16117), .ROB11(n16116), .ROB10(n16115), 
            .ROB9(n16114), .ROB8(n16113), .ROB7(n16112), .ROB6(n16111), 
            .ROB5(n16110), .ROB4(n16109), .ROB3(n16108), .ROB2(n16107), 
            .ROB1(n16106), .ROB0(n16105), .P35(n16159), .P34(n16158), 
            .P33(n16157), .P32(n16156), .P31(n16155), .P30(n16154), 
            .P29(n16153), .P28(n16152), .P27(n16151), .P26(n16150), 
            .P25(n16149), .P24(n16148), .P23(n16147), .P22(n16146), 
            .P21(n16145), .P20(n16144), .P19(n16143), .P18(n16142), 
            .P17(n16141), .P16(n16140), .P15(n16139), .P14(n16138), 
            .P13(n16137), .P12(n16136), .P11(n16135), .P10(n16134), 
            .P9(n16133), .P8(n16132), .P7(n16131), .P6(n16130), .P5(n16129), 
            .P4(n16128), .P3(n16127), .P2(n16126), .P1(n16125), .P0(n16124), 
            .SIGNEDP(n16123));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(52[13:28])
    defparam lat_mult_40.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_40.REG_INPUTA_CE = "CE3";
    defparam lat_mult_40.REG_INPUTA_RST = "RST3";
    defparam lat_mult_40.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_40.REG_INPUTB_CE = "CE0";
    defparam lat_mult_40.REG_INPUTB_RST = "RST0";
    defparam lat_mult_40.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_40.REG_INPUTC_CE = "CE0";
    defparam lat_mult_40.REG_INPUTC_RST = "RST0";
    defparam lat_mult_40.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_40.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_40.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_40.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_40.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_40.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_40.CLK0_DIV = "ENABLED";
    defparam lat_mult_40.CLK1_DIV = "ENABLED";
    defparam lat_mult_40.CLK2_DIV = "ENABLED";
    defparam lat_mult_40.CLK3_DIV = "ENABLED";
    defparam lat_mult_40.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_40.GSR = "DISABLED";
    defparam lat_mult_40.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_40.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_40.MULT_BYPASS = "DISABLED";
    defparam lat_mult_40.RESETMODE = "ASYNC";
    LUT4 i12681_4_lut (.A(n34843), .B(delay_r_23__N_1178[0]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[0]), .Z(dout_r_23__N_5926[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12681_4_lut.init = 16'hcac0;
    LUT4 i13012_4_lut (.A(n34843), .B(delay_r_23__N_1178[1]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[1]), .Z(dout_r_23__N_5926[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13012_4_lut.init = 16'hcac0;
    LUT4 i13014_4_lut (.A(n34843), .B(delay_r_23__N_1178[2]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[2]), .Z(dout_r_23__N_5926[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13014_4_lut.init = 16'hcac0;
    LUT4 i13016_4_lut (.A(n34843), .B(delay_r_23__N_1178[3]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[3]), .Z(dout_r_23__N_5926[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13016_4_lut.init = 16'hcac0;
    LUT4 i13018_4_lut (.A(n34843), .B(delay_r_23__N_1178[4]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[4]), .Z(dout_r_23__N_5926[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13018_4_lut.init = 16'hcac0;
    LUT4 i13020_4_lut (.A(n34843), .B(delay_r_23__N_1178[5]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[5]), .Z(dout_r_23__N_5926[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13020_4_lut.init = 16'hcac0;
    LUT4 i13022_4_lut (.A(n34843), .B(delay_r_23__N_1178[6]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[6]), .Z(dout_r_23__N_5926[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13022_4_lut.init = 16'hcac0;
    LUT4 i13024_4_lut (.A(n34843), .B(delay_r_23__N_1178[7]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[7]), .Z(dout_r_23__N_5926[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13024_4_lut.init = 16'hcac0;
    LUT4 i13026_4_lut (.A(n34843), .B(delay_r_23__N_1178[8]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[8]), .Z(dout_r_23__N_5926[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13026_4_lut.init = 16'hcac0;
    LUT4 i13028_4_lut (.A(n34843), .B(delay_r_23__N_1178[9]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[9]), .Z(dout_r_23__N_5926[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13028_4_lut.init = 16'hcac0;
    LUT4 i13030_4_lut (.A(n34843), .B(delay_r_23__N_1178[10]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[10]), .Z(dout_r_23__N_5926[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13030_4_lut.init = 16'hcac0;
    LUT4 i13032_4_lut (.A(n34843), .B(delay_r_23__N_1178[11]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[11]), .Z(dout_r_23__N_5926[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13032_4_lut.init = 16'hcac0;
    LUT4 i13034_4_lut (.A(n34843), .B(delay_r_23__N_1178[12]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[12]), .Z(dout_r_23__N_5926[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13034_4_lut.init = 16'hcac0;
    LUT4 i13036_4_lut (.A(n34843), .B(delay_r_23__N_1178[13]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[13]), .Z(dout_r_23__N_5926[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13036_4_lut.init = 16'hcac0;
    LUT4 i13038_4_lut (.A(n34843), .B(delay_r_23__N_1178[14]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[14]), .Z(dout_r_23__N_5926[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13038_4_lut.init = 16'hcac0;
    LUT4 i13040_4_lut (.A(n34843), .B(delay_r_23__N_1178[15]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[15]), .Z(dout_r_23__N_5926[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13040_4_lut.init = 16'hcac0;
    LUT4 i13042_4_lut (.A(n34843), .B(delay_r_23__N_1178[16]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[16]), .Z(dout_r_23__N_5926[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13042_4_lut.init = 16'hcac0;
    LUT4 i13044_4_lut (.A(n34843), .B(delay_r_23__N_1178[17]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[17]), .Z(dout_r_23__N_5926[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13044_4_lut.init = 16'hcac0;
    LUT4 i13046_4_lut (.A(n34843), .B(delay_r_23__N_1178[18]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[18]), .Z(dout_r_23__N_5926[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13046_4_lut.init = 16'hcac0;
    LUT4 i13048_4_lut (.A(n34843), .B(delay_r_23__N_1178[19]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[19]), .Z(dout_r_23__N_5926[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13048_4_lut.init = 16'hcac0;
    LUT4 i13050_4_lut (.A(n34843), .B(delay_r_23__N_1178[20]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[20]), .Z(dout_r_23__N_5926[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13050_4_lut.init = 16'hcac0;
    LUT4 i13052_4_lut (.A(n34843), .B(delay_r_23__N_1178[21]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[21]), .Z(dout_r_23__N_5926[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13052_4_lut.init = 16'hcac0;
    LUT4 i13054_4_lut (.A(n34843), .B(delay_r_23__N_1178[22]), .C(\no5_state[0] ), 
         .D(op_r_23__N_1106[22]), .Z(dout_r_23__N_5926[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i13054_4_lut.init = 16'hcac0;
    LUT4 i10831_4_lut (.A(op_r_23__N_1106[23]), .B(delay_r_23__N_1178[23]), 
         .C(\no5_state[0] ), .D(n34843), .Z(dout_r_23__N_5926[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i10831_4_lut.init = 16'hcac0;
    LUT4 i12447_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[16] ), 
         .D(\op_i_23__N_1154[8]_adj_1 ), .Z(\out_i[8] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12447_4_lut_4_lut.init = 16'hc480;
    LUT4 i12567_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[21] ), 
         .D(\op_i_23__N_1154[13]_adj_2 ), .Z(\out_i[13] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12567_4_lut_4_lut.init = 16'hc480;
    LUT4 i12568_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[20] ), 
         .D(\op_i_23__N_1154[12]_adj_3 ), .Z(\out_i[12] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12568_4_lut_4_lut.init = 16'hc480;
    LUT4 i12569_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[19] ), 
         .D(\op_i_23__N_1154[11]_adj_4 ), .Z(\out_i[11] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12569_4_lut_4_lut.init = 16'hc480;
    LUT4 i12570_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[18] ), 
         .D(\op_i_23__N_1154[10]_adj_5 ), .Z(\out_i[10] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12570_4_lut_4_lut.init = 16'hc480;
    LUT4 i12503_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[17] ), 
         .D(\op_i_23__N_1154[9]_adj_6 ), .Z(\out_i[9] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12503_4_lut_4_lut.init = 16'hc480;
    LUT4 i12557_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[31] ), 
         .D(\op_i_23__N_1154[23]_adj_7 ), .Z(\out_i[23] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12557_4_lut_4_lut.init = 16'hc480;
    LUT4 i12558_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[30] ), 
         .D(\op_i_23__N_1154[22]_adj_8 ), .Z(\out_i[22] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12558_4_lut_4_lut.init = 16'hc480;
    LUT4 i12559_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[29] ), 
         .D(\op_i_23__N_1154[21]_adj_9 ), .Z(\out_i[21] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12559_4_lut_4_lut.init = 16'hc480;
    LUT4 i12560_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[28] ), 
         .D(\op_i_23__N_1154[20]_adj_10 ), .Z(\out_i[20] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12560_4_lut_4_lut.init = 16'hc480;
    LUT4 i12561_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[27] ), 
         .D(\op_i_23__N_1154[19]_adj_11 ), .Z(\out_i[19] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12561_4_lut_4_lut.init = 16'hc480;
    LUT4 i12562_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[26] ), 
         .D(\op_i_23__N_1154[18]_adj_12 ), .Z(\out_i[18] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12562_4_lut_4_lut.init = 16'hc480;
    LUT4 i12563_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[25] ), 
         .D(\op_i_23__N_1154[17]_adj_13 ), .Z(\out_i[17] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12563_4_lut_4_lut.init = 16'hc480;
    LUT4 i12564_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[24] ), 
         .D(\op_i_23__N_1154[16]_adj_14 ), .Z(\out_i[16] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12564_4_lut_4_lut.init = 16'hc480;
    LUT4 i12565_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[23] ), 
         .D(\op_i_23__N_1154[15]_adj_15 ), .Z(\out_i[15] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12565_4_lut_4_lut.init = 16'hc480;
    LUT4 i12566_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_i_23__N_1130[22] ), 
         .D(\op_i_23__N_1154[14]_adj_16 ), .Z(\out_i[14] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12566_4_lut_4_lut.init = 16'hc480;
    LUT4 i12451_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[16] ), 
         .D(\op_r_23__N_1106[8]_adj_17 ), .Z(\out_r[8] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12451_4_lut_4_lut.init = 16'hc480;
    LUT4 i12571_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[17] ), 
         .D(\op_r_23__N_1106[9]_adj_18 ), .Z(\out_r[9] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12571_4_lut_4_lut.init = 16'hc480;
    LUT4 i12572_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[18] ), 
         .D(\op_r_23__N_1106[10]_adj_19 ), .Z(\out_r[10] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12572_4_lut_4_lut.init = 16'hc480;
    LUT4 i12573_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[19] ), 
         .D(\op_r_23__N_1106[11]_adj_20 ), .Z(\out_r[11] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12573_4_lut_4_lut.init = 16'hc480;
    LUT4 i12574_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[20] ), 
         .D(\op_r_23__N_1106[12]_adj_21 ), .Z(\out_r[12] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12574_4_lut_4_lut.init = 16'hc480;
    LUT4 i12575_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[21] ), 
         .D(\op_r_23__N_1106[13]_adj_22 ), .Z(\out_r[13] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12575_4_lut_4_lut.init = 16'hc480;
    LUT4 i12576_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[22] ), 
         .D(\op_r_23__N_1106[14]_adj_23 ), .Z(\out_r[14] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12576_4_lut_4_lut.init = 16'hc480;
    LUT4 i12577_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[23] ), 
         .D(\op_r_23__N_1106[15]_adj_24 ), .Z(\out_r[15] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12577_4_lut_4_lut.init = 16'hc480;
    LUT4 i12578_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[24] ), 
         .D(\op_r_23__N_1106[16]_adj_25 ), .Z(\out_r[16] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12578_4_lut_4_lut.init = 16'hc480;
    LUT4 i12579_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[25] ), 
         .D(\op_r_23__N_1106[17]_adj_26 ), .Z(\out_r[17] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12579_4_lut_4_lut.init = 16'hc480;
    LUT4 i12580_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[26] ), 
         .D(\op_r_23__N_1106[18]_adj_27 ), .Z(\out_r[18] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12580_4_lut_4_lut.init = 16'hc480;
    LUT4 i12581_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[27] ), 
         .D(\op_r_23__N_1106[19]_adj_28 ), .Z(\out_r[19] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12581_4_lut_4_lut.init = 16'hc480;
    LUT4 i12582_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[28] ), 
         .D(\op_r_23__N_1106[20]_adj_29 ), .Z(\out_r[20] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12582_4_lut_4_lut.init = 16'hc480;
    LUT4 i12583_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[29] ), 
         .D(\op_r_23__N_1106[21]_adj_30 ), .Z(\out_r[21] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12583_4_lut_4_lut.init = 16'hc480;
    LUT4 i12584_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[30] ), 
         .D(\op_r_23__N_1106[22]_adj_31 ), .Z(\out_r[22] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12584_4_lut_4_lut.init = 16'hc480;
    LUT4 i12585_4_lut_4_lut (.A(s5_count), .B(r4_valid), .C(\op_r_23__N_1082[31] ), 
         .D(\op_r_23__N_1106[23]_adj_32 ), .Z(\out_r[23] )) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/radix2.v(24[5] 68[12])
    defparam i12585_4_lut_4_lut.init = 16'hc480;
    
endmodule
//
// Verilog Description of module ROM_16
//

module ROM_16 (clk_c, n34737, n30203, \rom16_w_i[5] , \count[4] , 
            n30207, n33013, n30197, n34736, n32928, \count[5] , 
            n34735, \rom16_w_i[1] , \rom16_w_i[6] , n20089, \rom16_w_r[1] , 
            n28589, \rom16_w_r[2] , n20095, \rom16_w_r[3] , n20103, 
            \rom16_w_r[4] , n28591, \rom16_w_r[5] , \rom16_w_r[8] , 
            n17, GND_net, VCC_net, in_valid_reg, n34713, \rom16_w_i[8] , 
            n34727, \rom16_w_i[0] , \rom16_w_r[6] , n30499, \rom16_w_i[2] , 
            \rom16_w_i[3] , n33030, \rom16_w_i[4] , n34729, \rom16_w_i[7] , 
            n34730, n34789, \rom16_w_r[9] , n33051, n28598, \rom16_w_r[0] , 
            n34757, n34733, \op_i_23__N_1130[17] , \din_i_reg[9] , n31698, 
            \op_i_23__N_1130[16] , \din_i_reg[8] , n31700, \op_i_23__N_1130[19] , 
            \din_i_reg[11] , n31694, \op_i_23__N_1130[18] , \din_i_reg[10] , 
            n31696, \op_i_23__N_1130[21] , \din_i_reg[13] , n31690, 
            \op_i_23__N_1130[20] , \din_i_reg[12] , n31692, \op_i_23__N_1130[23] , 
            \din_i_reg[15] , n31686, \op_i_23__N_1130[22] , \din_i_reg[14] , 
            n31688, \op_i_23__N_1130[25] , \din_i_reg[17] , n31682, 
            \op_i_23__N_1130[24] , \din_i_reg[16] , n31684, \op_i_23__N_1130[27] , 
            \din_i_reg[23] , n31678, \op_i_23__N_1130[26] , \din_i_reg[18] , 
            n31680, \op_i_23__N_1130[29] , n31674, \op_i_23__N_1130[28] , 
            n31676, \op_i_23__N_1130[31] , n31670, \op_i_23__N_1130[30] , 
            n31672, \op_r_23__N_1082[17] , \din_r_reg[9] , n31731, \op_r_23__N_1082[16] , 
            \din_r_reg[8] , n31733, \rom16_w_r[7] , \op_r_23__N_1082[30] , 
            \din_r_reg[23] , n31705, \op_r_23__N_1082[31] , n31703, 
            \op_r_23__N_1082[28] , n31709, \op_r_23__N_1082[29] , n31707, 
            \op_r_23__N_1082[26] , \din_r_reg[18] , n31713, \op_r_23__N_1082[27] , 
            n31711, \op_r_23__N_1082[24] , \din_r_reg[16] , n31717, 
            \op_r_23__N_1082[25] , \din_r_reg[17] , n31715, \op_r_23__N_1082[22] , 
            \din_r_reg[14] , n31721, \op_r_23__N_1082[23] , \din_r_reg[15] , 
            n31719, \op_r_23__N_1082[20] , \din_r_reg[12] , n31725, 
            \op_r_23__N_1082[21] , \din_r_reg[13] , n31723, \op_r_23__N_1082[18] , 
            \din_r_reg[10] , n31729, \op_r_23__N_1082[19] , \din_r_reg[11] , 
            n31727, n34759) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n34737;
    output n30203;
    output \rom16_w_i[5] ;
    output \count[4] ;
    output n30207;
    output n33013;
    output n30197;
    output n34736;
    output n32928;
    output \count[5] ;
    output n34735;
    output \rom16_w_i[1] ;
    output \rom16_w_i[6] ;
    output n20089;
    output \rom16_w_r[1] ;
    output n28589;
    output \rom16_w_r[2] ;
    output n20095;
    output \rom16_w_r[3] ;
    output n20103;
    output \rom16_w_r[4] ;
    output n28591;
    output \rom16_w_r[5] ;
    output \rom16_w_r[8] ;
    output n17;
    input GND_net;
    input VCC_net;
    input in_valid_reg;
    output n34713;
    output \rom16_w_i[8] ;
    output n34727;
    output \rom16_w_i[0] ;
    output \rom16_w_r[6] ;
    output n30499;
    output \rom16_w_i[2] ;
    output \rom16_w_i[3] ;
    output n33030;
    output \rom16_w_i[4] ;
    output n34729;
    output \rom16_w_i[7] ;
    output n34730;
    output n34789;
    output \rom16_w_r[9] ;
    output n33051;
    output n28598;
    output \rom16_w_r[0] ;
    output n34757;
    output n34733;
    input \op_i_23__N_1130[17] ;
    input \din_i_reg[9] ;
    output n31698;
    input \op_i_23__N_1130[16] ;
    input \din_i_reg[8] ;
    output n31700;
    input \op_i_23__N_1130[19] ;
    input \din_i_reg[11] ;
    output n31694;
    input \op_i_23__N_1130[18] ;
    input \din_i_reg[10] ;
    output n31696;
    input \op_i_23__N_1130[21] ;
    input \din_i_reg[13] ;
    output n31690;
    input \op_i_23__N_1130[20] ;
    input \din_i_reg[12] ;
    output n31692;
    input \op_i_23__N_1130[23] ;
    input \din_i_reg[15] ;
    output n31686;
    input \op_i_23__N_1130[22] ;
    input \din_i_reg[14] ;
    output n31688;
    input \op_i_23__N_1130[25] ;
    input \din_i_reg[17] ;
    output n31682;
    input \op_i_23__N_1130[24] ;
    input \din_i_reg[16] ;
    output n31684;
    input \op_i_23__N_1130[27] ;
    input \din_i_reg[23] ;
    output n31678;
    input \op_i_23__N_1130[26] ;
    input \din_i_reg[18] ;
    output n31680;
    input \op_i_23__N_1130[29] ;
    output n31674;
    input \op_i_23__N_1130[28] ;
    output n31676;
    input \op_i_23__N_1130[31] ;
    output n31670;
    input \op_i_23__N_1130[30] ;
    output n31672;
    input \op_r_23__N_1082[17] ;
    input \din_r_reg[9] ;
    output n31731;
    input \op_r_23__N_1082[16] ;
    input \din_r_reg[8] ;
    output n31733;
    output \rom16_w_r[7] ;
    input \op_r_23__N_1082[30] ;
    input \din_r_reg[23] ;
    output n31705;
    input \op_r_23__N_1082[31] ;
    output n31703;
    input \op_r_23__N_1082[28] ;
    output n31709;
    input \op_r_23__N_1082[29] ;
    output n31707;
    input \op_r_23__N_1082[26] ;
    input \din_r_reg[18] ;
    output n31713;
    input \op_r_23__N_1082[27] ;
    output n31711;
    input \op_r_23__N_1082[24] ;
    input \din_r_reg[16] ;
    output n31717;
    input \op_r_23__N_1082[25] ;
    input \din_r_reg[17] ;
    output n31715;
    input \op_r_23__N_1082[22] ;
    input \din_r_reg[14] ;
    output n31721;
    input \op_r_23__N_1082[23] ;
    input \din_r_reg[15] ;
    output n31719;
    input \op_r_23__N_1082[20] ;
    input \din_r_reg[12] ;
    output n31725;
    input \op_r_23__N_1082[21] ;
    input \din_r_reg[13] ;
    output n31723;
    input \op_r_23__N_1082[18] ;
    input \din_r_reg[10] ;
    output n31729;
    input \op_r_23__N_1082[19] ;
    input \din_r_reg[11] ;
    output n31727;
    output n34759;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire valid, valid_N_3705, n34764;
    wire [5:0]count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(11[11:16])
    
    wire n34766, n28590, n34550, clk_c_enable_2289;
    wire [5:0]n29;
    
    wire n8, n34790, n33003, n34791, n34792, n29803, n7, n33043, 
        n33190, n33015, n33116, n34728, n34763, n34748, n34549, 
        n34758, n25, n34552, n34555, n34558, n32389, n32388, n32387, 
        n34559, n34556, n20105, n34783, n34744, n34743, n34746, 
        n34745, n34793, n34797, n34796, n30015, n34553, n34804, 
        n34781, n34803, n34784, n28370;
    
    FD1S3AX valid_47 (.D(valid_N_3705), .CK(clk_c), .Q(valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=106, LSE_RLINE=113 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(117[10] 126[8])
    defparam valid_47.GSR = "ENABLED";
    LUT4 i12489_2_lut_rep_375_3_lut_4_lut_4_lut (.A(n34764), .B(count[1]), 
         .C(count[2]), .D(n34766), .Z(n34737)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i12489_2_lut_rep_375_3_lut_4_lut_4_lut.init = 16'hfbcb;
    LUT4 i12493_2_lut_3_lut_4_lut_4_lut (.A(n34764), .B(count[1]), .C(count[2]), 
         .D(n34766), .Z(n30203)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B (C+(D))+!B !(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i12493_2_lut_3_lut_4_lut_4_lut.init = 16'hefe3;
    LUT4 i16333_3_lut_4_lut_4_lut (.A(n34764), .B(n34766), .C(count[1]), 
         .D(count[2]), .Z(\rom16_w_i[5] )) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;
    defparam i16333_3_lut_4_lut_4_lut.init = 16'h0770;
    LUT4 i10910_4_lut_4_lut (.A(\count[4] ), .B(count[3]), .C(count[2]), 
         .D(count[1]), .Z(n28590)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i10910_4_lut_4_lut.init = 16'hebbe;
    LUT4 count_0__bdd_4_lut_16453_4_lut (.A(\count[4] ), .B(count[3]), .C(count[1]), 
         .D(count[2]), .Z(n34550)) /* synthesis lut_function=(A+!(B (C)+!B !(C+!(D)))) */ ;
    defparam count_0__bdd_4_lut_16453_4_lut.init = 16'hbebf;
    FD1P3AX count_690__i0 (.D(n29[0]), .SP(clk_c_enable_2289), .CK(clk_c), 
            .Q(count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690__i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n30207), .B(n8), .C(n34790), .D(n33003), .Z(n33013)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h2220;
    LUT4 i1_4_lut_adj_21 (.A(n30203), .B(n30197), .C(n34737), .D(n34736), 
         .Z(n32928)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_21.init = 16'h8000;
    LUT4 i1_4_lut_adj_22 (.A(n34791), .B(\count[5] ), .C(count[0]), .D(n34792), 
         .Z(n29803)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_4_lut_adj_22.init = 16'hffbf;
    LUT4 count_5__I_0_52_i7_2_lut (.A(count[1]), .B(count[2]), .Z(n7)) /* synthesis lut_function=((B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(34[5:10])
    defparam count_5__I_0_52_i7_2_lut.init = 16'hdddd;
    LUT4 i12497_4_lut (.A(n33043), .B(n33190), .C(count[3]), .D(count[0]), 
         .Z(n30207)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;
    defparam i12497_4_lut.init = 16'h8aaa;
    LUT4 i1_4_lut_adj_23 (.A(count[0]), .B(n33015), .C(n34792), .D(n33116), 
         .Z(n8)) /* synthesis lut_function=(!(A+(B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_23.init = 16'h1511;
    LUT4 i16339_4_lut (.A(n8), .B(n30197), .C(n34728), .D(n34735), .Z(\rom16_w_i[1] )) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i16339_4_lut.init = 16'hbfff;
    LUT4 i16344_4_lut (.A(n34763), .B(n34737), .C(n34748), .D(n29803), 
         .Z(\rom16_w_i[6] )) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i16344_4_lut.init = 16'h7fff;
    LUT4 i12509_2_lut (.A(\count[5] ), .B(n20089), .Z(\rom16_w_r[1] )) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i12509_2_lut.init = 16'h2222;
    LUT4 count_0__bdd_4_lut_16450 (.A(\count[4] ), .B(count[3]), .C(count[1]), 
         .D(count[2]), .Z(n34549)) /* synthesis lut_function=(A+(B ((D)+!C)+!B !(C+!(D)))) */ ;
    defparam count_0__bdd_4_lut_16450.init = 16'hefae;
    LUT4 i12511_2_lut (.A(\count[5] ), .B(n28589), .Z(\rom16_w_r[2] )) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i12511_2_lut.init = 16'h2222;
    LUT4 i12513_2_lut (.A(\count[5] ), .B(n20095), .Z(\rom16_w_r[3] )) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i12513_2_lut.init = 16'h2222;
    LUT4 i12515_2_lut (.A(\count[5] ), .B(n20103), .Z(\rom16_w_r[4] )) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i12515_2_lut.init = 16'h2222;
    LUT4 i12517_2_lut (.A(\count[5] ), .B(n28591), .Z(\rom16_w_r[5] )) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i12517_2_lut.init = 16'h2222;
    LUT4 i1_3_lut (.A(\count[5] ), .B(n34758), .C(\count[4] ), .Z(\rom16_w_r[8] )) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_3_lut.init = 16'hfdfd;
    LUT4 i1_4_lut_adj_24 (.A(count[3]), .B(count[2]), .C(count[1]), .D(count[0]), 
         .Z(n25)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam i1_4_lut_adj_24.init = 16'h1734;
    LUT4 count_0__bdd_4_lut_16454 (.A(count[0]), .B(\count[4] ), .C(count[3]), 
         .D(count[2]), .Z(n34552)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C+(D)))) */ ;
    defparam count_0__bdd_4_lut_16454.init = 16'heccf;
    LUT4 n20077_bdd_2_lut (.A(\count[4] ), .B(count[1]), .Z(n34555)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n20077_bdd_2_lut.init = 16'heeee;
    LUT4 count_0__bdd_4_lut_16460 (.A(\count[4] ), .B(count[1]), .C(count[2]), 
         .D(count[3]), .Z(n34558)) /* synthesis lut_function=(A+!(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam count_0__bdd_4_lut_16460.init = 16'hbeeb;
    LUT4 i16347_2_lut (.A(\count[4] ), .B(n25), .Z(n17)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i16347_2_lut.init = 16'hbbbb;
    CCU2C count_690_add_4_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32389), .S0(n29[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690_add_4_7.INIT0 = 16'haaa0;
    defparam count_690_add_4_7.INIT1 = 16'h0000;
    defparam count_690_add_4_7.INJECT1_0 = "NO";
    defparam count_690_add_4_7.INJECT1_1 = "NO";
    CCU2C count_690_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(\count[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n32388), .COUT(n32389), .S0(n29[3]), .S1(n29[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690_add_4_5.INIT0 = 16'haaa0;
    defparam count_690_add_4_5.INIT1 = 16'haaa0;
    defparam count_690_add_4_5.INJECT1_0 = "NO";
    defparam count_690_add_4_5.INJECT1_1 = "NO";
    CCU2C count_690_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32387), .COUT(n32388), .S0(n29[1]), .S1(n29[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690_add_4_3.INIT0 = 16'haaa0;
    defparam count_690_add_4_3.INIT1 = 16'haaa0;
    defparam count_690_add_4_3.INJECT1_0 = "NO";
    defparam count_690_add_4_3.INJECT1_1 = "NO";
    CCU2C count_690_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(in_valid_reg), .B1(valid), .C1(count[0]), 
          .D1(VCC_net), .COUT(n32387), .S1(n29[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690_add_4_1.INIT0 = 16'h0000;
    defparam count_690_add_4_1.INIT1 = 16'h1e1e;
    defparam count_690_add_4_1.INJECT1_0 = "NO";
    defparam count_690_add_4_1.INJECT1_1 = "NO";
    PFUMX i16461 (.BLUT(n34559), .ALUT(n34558), .C0(count[0]), .Z(n28589));
    PFUMX i16457 (.BLUT(n34556), .ALUT(n34555), .C0(count[0]), .Z(n20095));
    LUT4 i1_2_lut_rep_351 (.A(n33013), .B(n32928), .Z(n34713)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_351.init = 16'h8888;
    LUT4 i52_1_lut_2_lut (.A(n33013), .B(n32928), .Z(\rom16_w_i[8] )) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i52_1_lut_2_lut.init = 16'h7777;
    LUT4 i1_3_lut_rep_365 (.A(n34735), .B(n8), .C(n30207), .Z(n34727)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_365.init = 16'h2020;
    LUT4 i13313_1_lut_3_lut (.A(n34735), .B(n8), .C(n30207), .Z(\rom16_w_i[0] )) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i13313_1_lut_3_lut.init = 16'hdfdf;
    LUT4 i12519_2_lut_4_lut (.A(n20105), .B(n34783), .C(count[0]), .D(\count[5] ), 
         .Z(\rom16_w_r[6] )) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam i12519_2_lut_4_lut.init = 16'h3500;
    LUT4 i12789_2_lut_4_lut (.A(n34763), .B(n34744), .C(n34743), .D(n8), 
         .Z(n30499)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i12789_2_lut_4_lut.init = 16'h0080;
    LUT4 i16335_3_lut_4_lut (.A(n34748), .B(n29803), .C(n30207), .D(n30197), 
         .Z(\rom16_w_i[2] )) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i16335_3_lut_4_lut.init = 16'h7fff;
    LUT4 i16337_3_lut_4_lut (.A(n34748), .B(n29803), .C(n30197), .D(n34735), 
         .Z(\rom16_w_i[3] )) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i16337_3_lut_4_lut.init = 16'h7fff;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n34748), .B(n29803), .C(n30197), .D(n34737), 
         .Z(n33030)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i16341_2_lut_3_lut_4_lut (.A(n34746), .B(n34745), .C(n30197), 
         .D(n8), .Z(\rom16_w_i[4] )) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i16341_2_lut_3_lut_4_lut.init = 16'hff7f;
    LUT4 i1_2_lut_rep_366_3_lut_4_lut (.A(n34746), .B(n34745), .C(n29803), 
         .D(n34748), .Z(n34728)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_366_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_rep_373_4_lut (.A(n34766), .B(n7), .C(n34744), .D(n34763), 
         .Z(n34735)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_3_lut_rep_373_4_lut.init = 16'he000;
    LUT4 i12537_2_lut_rep_367_3_lut_4_lut (.A(n34766), .B(n34793), .C(n8), 
         .D(n34746), .Z(n34729)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i12537_2_lut_rep_367_3_lut_4_lut.init = 16'h0e00;
    LUT4 i12528_1_lut_2_lut_3_lut_4_lut (.A(n34766), .B(n34797), .C(n30197), 
         .D(n29803), .Z(\rom16_w_i[7] )) /* synthesis lut_function=(!(A (C (D))+!A !(B+!(C (D))))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i12528_1_lut_2_lut_3_lut_4_lut.init = 16'h4fff;
    LUT4 valid_I_0_3_lut_4_lut (.A(n34766), .B(n34797), .C(valid), .D(in_valid_reg), 
         .Z(valid_N_3705)) /* synthesis lut_function=(A (C+(D))+!A (B (D)+!B (C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam valid_I_0_3_lut_4_lut.init = 16'hffb0;
    LUT4 i12527_2_lut_rep_368_3_lut_4_lut (.A(n34766), .B(n34797), .C(n30197), 
         .D(n29803), .Z(n34730)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i12527_2_lut_rep_368_3_lut_4_lut.init = 16'hb000;
    LUT4 i1_3_lut_4_lut (.A(count[0]), .B(n34791), .C(\count[5] ), .D(n34789), 
         .Z(\rom16_w_r[9] )) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n34790), .B(n34793), .C(n34746), .D(n34766), 
         .Z(n33051)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_3_lut_4_lut_4_lut.init = 16'he0c0;
    LUT4 i1_2_lut_rep_384_4_lut (.A(count[0]), .B(\count[5] ), .C(n34792), 
         .D(n7), .Z(n34746)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_384_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_382_4_lut (.A(count[0]), .B(\count[5] ), .C(n34792), 
         .D(n34793), .Z(n34744)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_382_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_4_lut (.A(count[0]), .B(\count[5] ), .C(n34792), .D(n34797), 
         .Z(n33043)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_4_lut.init = 16'hf7ff;
    LUT4 i1_2_lut_rep_381_4_lut (.A(n34796), .B(count[0]), .C(\count[4] ), 
         .D(n7), .Z(n34743)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_381_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_383_4_lut (.A(n34796), .B(count[0]), .C(\count[4] ), 
         .D(n34793), .Z(n34745)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_383_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_386_4_lut (.A(n34796), .B(count[0]), .C(\count[4] ), 
         .D(n34797), .Z(n34748)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_386_4_lut.init = 16'hf7ff;
    LUT4 i2408_3_lut_4_lut_4_lut (.A(\count[4] ), .B(count[3]), .C(count[2]), 
         .D(count[1]), .Z(n20105)) /* synthesis lut_function=(A+(B ((D)+!C)+!B !(D))) */ ;
    defparam i2408_3_lut_4_lut_4_lut.init = 16'heebf;
    LUT4 in_valid_I_0_2_lut_rep_410 (.A(in_valid_reg), .B(valid), .Z(clk_c_enable_2289)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[8:25])
    defparam in_valid_I_0_2_lut_rep_410.init = 16'heeee;
    LUT4 i12305_3_lut_4_lut (.A(in_valid_reg), .B(valid), .C(n29[5]), 
         .D(\count[5] ), .Z(n30015)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[8:25])
    defparam i12305_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i16455 (.BLUT(n34553), .ALUT(n34552), .C0(count[1]), .Z(n20089));
    LUT4 i16353_4_lut_then_4_lut (.A(count[0]), .B(\count[4] ), .C(n34797), 
         .D(\count[5] ), .Z(n34804)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i16353_4_lut_then_4_lut.init = 16'hefff;
    LUT4 i10895_2_lut_4_lut_4_lut (.A(count[3]), .B(count[2]), .C(\count[4] ), 
         .D(n34781), .Z(n28598)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i10895_2_lut_4_lut_4_lut.init = 16'hfaf9;
    LUT4 i10663_2_lut_rep_419 (.A(count[1]), .B(count[0]), .Z(n34781)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10663_2_lut_rep_419.init = 16'heeee;
    LUT4 i10664_3_lut_rep_396_3_lut_4_lut (.A(count[1]), .B(count[0]), .C(count[2]), 
         .D(count[3]), .Z(n34758)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam i10664_3_lut_rep_396_3_lut_4_lut.init = 16'hfe01;
    LUT4 i16353_4_lut_else_4_lut (.A(count[0]), .B(\count[4] ), .C(n7), 
         .D(\count[5] ), .Z(n34803)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i16353_4_lut_else_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_4_lut_4_lut (.A(count[3]), .B(count[2]), .C(n34784), 
         .D(n34781), .Z(\rom16_w_r[0] )) /* synthesis lut_function=(A (B (C))+!A !(B ((D)+!C)+!B !(C (D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h90c0;
    LUT4 i10903_3_lut_rep_395_4_lut_4_lut (.A(count[3]), .B(count[2]), .C(count[0]), 
         .D(count[1]), .Z(n34757)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;
    defparam i10903_3_lut_rep_395_4_lut_4_lut.init = 16'h6663;
    LUT4 i2393_2_lut_rep_421 (.A(\count[4] ), .B(count[2]), .Z(n34783)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2393_2_lut_rep_421.init = 16'heeee;
    LUT4 i2409_3_lut_rep_371_4_lut (.A(\count[4] ), .B(count[2]), .C(count[0]), 
         .D(n20105), .Z(n34733)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i2409_3_lut_rep_371_4_lut.init = 16'hefe0;
    LUT4 i1_2_lut_rep_422 (.A(\count[4] ), .B(\count[5] ), .Z(n34784)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_422.init = 16'h4444;
    LUT4 i13953_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[17] ), 
         .D(\din_i_reg[9] ), .Z(n31698)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13953_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13955_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[16] ), 
         .D(\din_i_reg[8] ), .Z(n31700)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13955_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13949_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[19] ), 
         .D(\din_i_reg[11] ), .Z(n31694)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13949_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13951_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[18] ), 
         .D(\din_i_reg[10] ), .Z(n31696)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13951_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13945_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[21] ), 
         .D(\din_i_reg[13] ), .Z(n31690)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13945_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13947_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[20] ), 
         .D(\din_i_reg[12] ), .Z(n31692)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13947_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13941_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[23] ), 
         .D(\din_i_reg[15] ), .Z(n31686)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13941_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13943_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[22] ), 
         .D(\din_i_reg[14] ), .Z(n31688)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13943_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13937_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[25] ), 
         .D(\din_i_reg[17] ), .Z(n31682)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13937_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13939_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[24] ), 
         .D(\din_i_reg[16] ), .Z(n31684)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13939_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13933_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[27] ), 
         .D(\din_i_reg[23] ), .Z(n31678)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13933_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13935_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[26] ), 
         .D(\din_i_reg[18] ), .Z(n31680)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13935_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13929_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[29] ), 
         .D(\din_i_reg[23] ), .Z(n31674)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13929_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13931_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[28] ), 
         .D(\din_i_reg[23] ), .Z(n31676)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13931_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13925_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[31] ), 
         .D(\din_i_reg[23] ), .Z(n31670)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13925_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13927_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_i_23__N_1130[30] ), 
         .D(\din_i_reg[23] ), .Z(n31672)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13927_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13986_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[17] ), 
         .D(\din_r_reg[9] ), .Z(n31731)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13986_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13988_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[16] ), 
         .D(\din_r_reg[8] ), .Z(n31733)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13988_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_3_lut (.A(\count[4] ), .B(\count[5] ), .C(n25), .Z(\rom16_w_r[7] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 i13960_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[30] ), 
         .D(\din_r_reg[23] ), .Z(n31705)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13960_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13958_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[31] ), 
         .D(\din_r_reg[23] ), .Z(n31703)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13958_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13964_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[28] ), 
         .D(\din_r_reg[23] ), .Z(n31709)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13964_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13962_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[29] ), 
         .D(\din_r_reg[23] ), .Z(n31707)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13962_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13968_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[26] ), 
         .D(\din_r_reg[18] ), .Z(n31713)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13968_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13966_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[27] ), 
         .D(\din_r_reg[23] ), .Z(n31711)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13966_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13972_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[24] ), 
         .D(\din_r_reg[16] ), .Z(n31717)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13972_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13970_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[25] ), 
         .D(\din_r_reg[17] ), .Z(n31715)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13970_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13976_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[22] ), 
         .D(\din_r_reg[14] ), .Z(n31721)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13976_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13974_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[23] ), 
         .D(\din_r_reg[15] ), .Z(n31719)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13974_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13980_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[20] ), 
         .D(\din_r_reg[12] ), .Z(n31725)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13980_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13978_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[21] ), 
         .D(\din_r_reg[13] ), .Z(n31723)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13978_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13984_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[18] ), 
         .D(\din_r_reg[10] ), .Z(n31729)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13984_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13982_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(\op_r_23__N_1082[19] ), 
         .D(\din_r_reg[11] ), .Z(n31727)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13982_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2380_2_lut_rep_427 (.A(\count[4] ), .B(count[3]), .Z(n34789)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i2380_2_lut_rep_427.init = 16'hbbbb;
    LUT4 n20077_bdd_4_lut_4_lut (.A(\count[4] ), .B(count[3]), .C(count[2]), 
         .D(count[1]), .Z(n34556)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;
    defparam n20077_bdd_4_lut_4_lut.init = 16'hfabf;
    LUT4 count_0__bdd_4_lut_16459_4_lut (.A(\count[4] ), .B(count[3]), .C(count[2]), 
         .D(count[0]), .Z(n34553)) /* synthesis lut_function=(A+!(B (C+(D))+!B (D))) */ ;
    defparam count_0__bdd_4_lut_16459_4_lut.init = 16'haabf;
    LUT4 i1_3_lut_4_lut_adj_25 (.A(\count[4] ), .B(count[3]), .C(\count[5] ), 
         .D(n7), .Z(n33015)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_3_lut_4_lut_adj_25.init = 16'hffbf;
    LUT4 i1_3_lut_rep_428 (.A(\count[5] ), .B(\count[4] ), .C(count[0]), 
         .Z(n34790)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_3_lut_rep_428.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_401_4_lut (.A(\count[5] ), .B(\count[4] ), .C(count[0]), 
         .D(n34793), .Z(n34763)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_401_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_429 (.A(count[1]), .B(count[2]), .Z(n34791)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_429.init = 16'heeee;
    LUT4 i12796_2_lut_rep_397_3_lut (.A(count[1]), .B(count[2]), .C(count[0]), 
         .Z(n34759)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i12796_2_lut_rep_397_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_26 (.A(count[1]), .B(count[2]), .C(\count[4] ), 
         .D(\count[5] ), .Z(n33190)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_26.init = 16'hfeff;
    LUT4 i1_2_lut_rep_430 (.A(\count[4] ), .B(count[3]), .Z(n34792)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_2_lut_rep_430.init = 16'heeee;
    LUT4 count_0__bdd_4_lut_4_lut (.A(\count[4] ), .B(count[3]), .C(count[2]), 
         .D(count[1]), .Z(n34559)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam count_0__bdd_4_lut_4_lut.init = 16'hfaef;
    LUT4 i1_3_lut_rep_402_4_lut (.A(\count[4] ), .B(count[3]), .C(\count[5] ), 
         .D(count[0]), .Z(n34764)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_3_lut_rep_402_4_lut.init = 16'hefff;
    LUT4 i10671_2_lut_3_lut_4_lut (.A(\count[4] ), .B(count[3]), .C(count[2]), 
         .D(count[1]), .Z(n28370)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i10671_2_lut_3_lut_4_lut.init = 16'heeef;
    LUT4 count_5__I_0_55_i7_2_lut_rep_431 (.A(count[1]), .B(count[2]), .Z(n34793)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam count_5__I_0_55_i7_2_lut_rep_431.init = 16'hbbbb;
    LUT4 i1_3_lut_4_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), 
         .Z(n33003)) /* synthesis lut_function=(A+!(B+(C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(49[5:10])
    defparam i1_3_lut_4_lut_3_lut.init = 16'habab;
    LUT4 i1_2_lut_rep_434 (.A(\count[5] ), .B(count[3]), .Z(n34796)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_434.init = 16'h8888;
    LUT4 i1_3_lut_rep_404_4_lut (.A(\count[5] ), .B(count[3]), .C(\count[4] ), 
         .D(count[0]), .Z(n34766)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_3_lut_rep_404_4_lut.init = 16'hf7ff;
    LUT4 i12523_2_lut_rep_435 (.A(count[1]), .B(count[2]), .Z(n34797)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12523_2_lut_rep_435.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_27 (.A(count[1]), .B(count[2]), .C(\count[5] ), 
         .Z(n33116)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_27.init = 16'h8080;
    LUT4 i1_2_lut_rep_374_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(n29803), 
         .D(n34766), .Z(n34736)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_rep_374_3_lut_4_lut.init = 16'hf070;
    PFUMX i10891 (.BLUT(n28370), .ALUT(n28590), .C0(count[0]), .Z(n28591));
    PFUMX i16451 (.BLUT(n34550), .ALUT(n34549), .C0(count[0]), .Z(n20103));
    PFUMX i16466 (.BLUT(n34803), .ALUT(n34804), .C0(count[3]), .Z(n30197));
    FD1S3AX count_690__i5 (.D(n30015), .CK(clk_c), .Q(\count[5] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690__i5.GSR = "ENABLED";
    FD1P3AX count_690__i1 (.D(n29[1]), .SP(clk_c_enable_2289), .CK(clk_c), 
            .Q(count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690__i1.GSR = "ENABLED";
    FD1P3AX count_690__i2 (.D(n29[2]), .SP(clk_c_enable_2289), .CK(clk_c), 
            .Q(count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690__i2.GSR = "ENABLED";
    FD1P3AX count_690__i3 (.D(n29[3]), .SP(clk_c_enable_2289), .CK(clk_c), 
            .Q(count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690__i3.GSR = "ENABLED";
    FD1P3AX count_690__i4 (.D(n29[4]), .SP(clk_c_enable_2289), .CK(clk_c), 
            .Q(\count[4] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_16.v(13[39:48])
    defparam count_690__i4.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module shift_16
//

module shift_16 (clk_c, in_valid_reg, VCC_net, \op_i_23__N_1154[7] , 
            \op_i_23__N_1154[6] , \op_i_23__N_1154[5] , \op_i_23__N_1154[4] , 
            \op_i_23__N_1154[3] , \op_i_23__N_1154[2] , \op_i_23__N_1154[1] , 
            \op_r_23__N_1106[7] , \op_r_23__N_1106[6] , \op_r_23__N_1106[5] , 
            \op_r_23__N_1106[4] , \op_r_23__N_1106[3] , \op_r_23__N_1106[2] , 
            \op_r_23__N_1106[1] , \op_i_23__N_1154[0] , \op_r_23__N_1106[0] , 
            \dout_r_23__N_2506[8] , \dout_r_23__N_2506[9] , \dout_r_23__N_2506[10] , 
            \dout_r_23__N_2506[11] , \dout_r_23__N_2506[12] , \dout_r_23__N_2506[13] , 
            \dout_r_23__N_2506[14] , \dout_r_23__N_2506[15] , \dout_r_23__N_2506[16] , 
            \dout_r_23__N_2506[17] , \dout_r_23__N_2506[18] , \dout_r_23__N_2506[19] , 
            \dout_r_23__N_2506[20] , \dout_r_23__N_2506[21] , \dout_r_23__N_2506[22] , 
            \dout_r_23__N_2506[23] , \shift_16_dout_i[23] , \shift_16_dout_i[22] , 
            \shift_16_dout_i[21] , \shift_16_dout_i[20] , \shift_16_dout_i[19] , 
            \shift_16_dout_i[18] , \shift_16_dout_i[17] , \shift_16_dout_i[16] , 
            \shift_16_dout_i[15] , \shift_16_dout_i[14] , \shift_16_dout_i[13] , 
            \shift_16_dout_i[12] , \shift_16_dout_i[11] , \shift_16_dout_i[10] , 
            \shift_16_dout_i[9] , \shift_16_dout_i[8] , \shift_16_dout_r[23] , 
            \shift_16_dout_r[22] , \shift_16_dout_r[21] , \shift_16_dout_r[20] , 
            \shift_16_dout_r[19] , \shift_16_dout_r[18] , \shift_16_dout_r[17] , 
            \shift_16_dout_r[16] , \shift_16_dout_r[15] , \shift_16_dout_r[13] , 
            \shift_16_dout_r[12] , \shift_16_dout_r[11] , \shift_16_dout_r[10] , 
            \shift_16_dout_r[9] , \shift_16_dout_r[8] , \shift_16_dout_r[14] , 
            \count[5] , \count[4] , \dout_i_23__N_3274[8] , \dout_i_23__N_3274[9] , 
            \dout_i_23__N_3274[10] , \dout_i_23__N_3274[11] , \dout_i_23__N_3274[12] , 
            \dout_i_23__N_3274[13] , \dout_i_23__N_3274[14] , \dout_i_23__N_3274[15] , 
            \dout_i_23__N_3274[16] , \dout_i_23__N_3274[17] , \dout_i_23__N_3274[18] , 
            \dout_i_23__N_3274[19] , \dout_i_23__N_3274[20] , \dout_i_23__N_3274[21] , 
            \dout_i_23__N_3274[22] , \dout_i_23__N_3274[23] ) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input in_valid_reg;
    input VCC_net;
    output \op_i_23__N_1154[7] ;
    output \op_i_23__N_1154[6] ;
    output \op_i_23__N_1154[5] ;
    output \op_i_23__N_1154[4] ;
    output \op_i_23__N_1154[3] ;
    output \op_i_23__N_1154[2] ;
    output \op_i_23__N_1154[1] ;
    output \op_r_23__N_1106[7] ;
    output \op_r_23__N_1106[6] ;
    output \op_r_23__N_1106[5] ;
    output \op_r_23__N_1106[4] ;
    output \op_r_23__N_1106[3] ;
    output \op_r_23__N_1106[2] ;
    output \op_r_23__N_1106[1] ;
    output \op_i_23__N_1154[0] ;
    output \op_r_23__N_1106[0] ;
    input \dout_r_23__N_2506[8] ;
    input \dout_r_23__N_2506[9] ;
    input \dout_r_23__N_2506[10] ;
    input \dout_r_23__N_2506[11] ;
    input \dout_r_23__N_2506[12] ;
    input \dout_r_23__N_2506[13] ;
    input \dout_r_23__N_2506[14] ;
    input \dout_r_23__N_2506[15] ;
    input \dout_r_23__N_2506[16] ;
    input \dout_r_23__N_2506[17] ;
    input \dout_r_23__N_2506[18] ;
    input \dout_r_23__N_2506[19] ;
    input \dout_r_23__N_2506[20] ;
    input \dout_r_23__N_2506[21] ;
    input \dout_r_23__N_2506[22] ;
    input \dout_r_23__N_2506[23] ;
    output \shift_16_dout_i[23] ;
    output \shift_16_dout_i[22] ;
    output \shift_16_dout_i[21] ;
    output \shift_16_dout_i[20] ;
    output \shift_16_dout_i[19] ;
    output \shift_16_dout_i[18] ;
    output \shift_16_dout_i[17] ;
    output \shift_16_dout_i[16] ;
    output \shift_16_dout_i[15] ;
    output \shift_16_dout_i[14] ;
    output \shift_16_dout_i[13] ;
    output \shift_16_dout_i[12] ;
    output \shift_16_dout_i[11] ;
    output \shift_16_dout_i[10] ;
    output \shift_16_dout_i[9] ;
    output \shift_16_dout_i[8] ;
    output \shift_16_dout_r[23] ;
    output \shift_16_dout_r[22] ;
    output \shift_16_dout_r[21] ;
    output \shift_16_dout_r[20] ;
    output \shift_16_dout_r[19] ;
    output \shift_16_dout_r[18] ;
    output \shift_16_dout_r[17] ;
    output \shift_16_dout_r[16] ;
    output \shift_16_dout_r[15] ;
    output \shift_16_dout_r[13] ;
    output \shift_16_dout_r[12] ;
    output \shift_16_dout_r[11] ;
    output \shift_16_dout_r[10] ;
    output \shift_16_dout_r[9] ;
    output \shift_16_dout_r[8] ;
    output \shift_16_dout_r[14] ;
    input \count[5] ;
    input \count[4] ;
    input \dout_i_23__N_3274[8] ;
    input \dout_i_23__N_3274[9] ;
    input \dout_i_23__N_3274[10] ;
    input \dout_i_23__N_3274[11] ;
    input \dout_i_23__N_3274[12] ;
    input \dout_i_23__N_3274[13] ;
    input \dout_i_23__N_3274[14] ;
    input \dout_i_23__N_3274[15] ;
    input \dout_i_23__N_3274[16] ;
    input \dout_i_23__N_3274[17] ;
    input \dout_i_23__N_3274[18] ;
    input \dout_i_23__N_3274[19] ;
    input \dout_i_23__N_3274[20] ;
    input \dout_i_23__N_3274[21] ;
    input \dout_i_23__N_3274[22] ;
    input \dout_i_23__N_3274[23] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire valid;
    wire [383:0]dout_i_23__N_3274;
    
    wire clk_c_enable_1772, n29834;
    wire [383:0]dout_r_23__N_2506;
    
    wire n29919, n29920, n29921, n29922, n29923, n29924, n29925, 
        n29926, n29927, n29928, n29929, n29930, n29931, n29932, 
        n29933, n29934, n29935, n29936, n29937, n29938, n29939, 
        n29940, n29941, n29942, n29943, n29944, n29945, n29946, 
        n29947, n29948, n29949, n29950, n29951, n29953, n29954, 
        n29955, n29956, n29957, n29958, n29959, n29960, n29952, 
        n29961, n29962, n29963, n29964, n29965, n29966;
    
    FD1P3AX valid_26 (.D(VCC_net), .SP(in_valid_reg), .CK(clk_c), .Q(valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam valid_26.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i7 (.D(\op_i_23__N_1154[7] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i7.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i6 (.D(\op_i_23__N_1154[6] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i6.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i5 (.D(\op_i_23__N_1154[5] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i5.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i4 (.D(\op_i_23__N_1154[4] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i4.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i3 (.D(\op_i_23__N_1154[3] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i3.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i2 (.D(\op_i_23__N_1154[2] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i2.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i1 (.D(\op_i_23__N_1154[1] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i1.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i7 (.D(\op_r_23__N_1106[7] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i7.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i6 (.D(\op_r_23__N_1106[6] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i6.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i5 (.D(\op_r_23__N_1106[5] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i5.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i4 (.D(\op_r_23__N_1106[4] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i4.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i3 (.D(\op_r_23__N_1106[3] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i3.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i2 (.D(\op_r_23__N_1106[2] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i2.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i1 (.D(\op_r_23__N_1106[1] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i1.GSR = "ENABLED";
    FD1P3IX shift_reg_i_i0_i0 (.D(\op_i_23__N_1154[0] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_i_23__N_3274[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i0.GSR = "ENABLED";
    FD1P3IX shift_reg_r_i0_i0 (.D(\op_r_23__N_1106[0] ), .SP(clk_c_enable_1772), 
            .CD(n29834), .CK(clk_c), .Q(dout_r_23__N_2506[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i0.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i8 (.D(\dout_r_23__N_2506[8] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i8.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i9 (.D(\dout_r_23__N_2506[9] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i9.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i10 (.D(\dout_r_23__N_2506[10] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i10.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i11 (.D(\dout_r_23__N_2506[11] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i11.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i12 (.D(\dout_r_23__N_2506[12] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i12.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i13 (.D(\dout_r_23__N_2506[13] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i13.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i14 (.D(\dout_r_23__N_2506[14] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i14.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i15 (.D(\dout_r_23__N_2506[15] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i15.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i16 (.D(\dout_r_23__N_2506[16] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i16.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i17 (.D(\dout_r_23__N_2506[17] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i17.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i18 (.D(\dout_r_23__N_2506[18] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i18.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i19 (.D(\dout_r_23__N_2506[19] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i19.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i20 (.D(\dout_r_23__N_2506[20] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i20.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i21 (.D(\dout_r_23__N_2506[21] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i21.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i22 (.D(\dout_r_23__N_2506[22] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i22.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i23 (.D(\dout_r_23__N_2506[23] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i23.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i24 (.D(dout_r_23__N_2506[24]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i24.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i25 (.D(dout_r_23__N_2506[25]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i25.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i26 (.D(dout_r_23__N_2506[26]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i26.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i27 (.D(dout_r_23__N_2506[27]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i27.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i28 (.D(dout_r_23__N_2506[28]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i28.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i29 (.D(dout_r_23__N_2506[29]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i29.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i30 (.D(dout_r_23__N_2506[30]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i30.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i31 (.D(dout_r_23__N_2506[31]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i31.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i32 (.D(dout_r_23__N_2506[32]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i32.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i33 (.D(dout_r_23__N_2506[33]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i33.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i34 (.D(dout_r_23__N_2506[34]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i34.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i35 (.D(dout_r_23__N_2506[35]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i35.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i36 (.D(dout_r_23__N_2506[36]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i36.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i37 (.D(dout_r_23__N_2506[37]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i37.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i38 (.D(dout_r_23__N_2506[38]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i38.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i39 (.D(dout_r_23__N_2506[39]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i39.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i40 (.D(dout_r_23__N_2506[40]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i40.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i41 (.D(dout_r_23__N_2506[41]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i41.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i42 (.D(dout_r_23__N_2506[42]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i42.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i43 (.D(dout_r_23__N_2506[43]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i43.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i44 (.D(dout_r_23__N_2506[44]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i44.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i45 (.D(dout_r_23__N_2506[45]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i45.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i46 (.D(dout_r_23__N_2506[46]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i46.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i47 (.D(dout_r_23__N_2506[47]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i47.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i48 (.D(dout_r_23__N_2506[48]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i48.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i49 (.D(dout_r_23__N_2506[49]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i49.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i50 (.D(dout_r_23__N_2506[50]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i50.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i51 (.D(dout_r_23__N_2506[51]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i51.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i52 (.D(dout_r_23__N_2506[52]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i52.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i53 (.D(dout_r_23__N_2506[53]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[77])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i53.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i54 (.D(dout_r_23__N_2506[54]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[78])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i54.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i55 (.D(dout_r_23__N_2506[55]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[79])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i55.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i56 (.D(dout_r_23__N_2506[56]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i56.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i57 (.D(dout_r_23__N_2506[57]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i57.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i58 (.D(dout_r_23__N_2506[58]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i58.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i59 (.D(dout_r_23__N_2506[59]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i59.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i60 (.D(dout_r_23__N_2506[60]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i60.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i61 (.D(dout_r_23__N_2506[61]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[85])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i61.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i62 (.D(dout_r_23__N_2506[62]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[86])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i62.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i63 (.D(dout_r_23__N_2506[63]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[87])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i63.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i64 (.D(dout_r_23__N_2506[64]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i64.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i65 (.D(dout_r_23__N_2506[65]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i65.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i66 (.D(dout_r_23__N_2506[66]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i66.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i67 (.D(dout_r_23__N_2506[67]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i67.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i68 (.D(dout_r_23__N_2506[68]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i68.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i69 (.D(dout_r_23__N_2506[69]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[93])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i69.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i70 (.D(dout_r_23__N_2506[70]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[94])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i70.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i71 (.D(dout_r_23__N_2506[71]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[95])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i71.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i72 (.D(dout_r_23__N_2506[72]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[96])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i72.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i73 (.D(dout_r_23__N_2506[73]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[97])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i73.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i74 (.D(dout_r_23__N_2506[74]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[98])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i74.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i75 (.D(dout_r_23__N_2506[75]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[99])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i75.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i76 (.D(dout_r_23__N_2506[76]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[100])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i76.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i77 (.D(dout_r_23__N_2506[77]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[101])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i77.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i78 (.D(dout_r_23__N_2506[78]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[102])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i78.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i79 (.D(dout_r_23__N_2506[79]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[103])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i79.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i80 (.D(dout_r_23__N_2506[80]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[104])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i80.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i81 (.D(dout_r_23__N_2506[81]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[105])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i81.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i82 (.D(dout_r_23__N_2506[82]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[106])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i82.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i83 (.D(dout_r_23__N_2506[83]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[107])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i83.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i84 (.D(dout_r_23__N_2506[84]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[108])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i84.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i85 (.D(dout_r_23__N_2506[85]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[109])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i85.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i86 (.D(dout_r_23__N_2506[86]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[110])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i86.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i87 (.D(dout_r_23__N_2506[87]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[111])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i87.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i88 (.D(dout_r_23__N_2506[88]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[112])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i88.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i89 (.D(dout_r_23__N_2506[89]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[113])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i89.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i90 (.D(dout_r_23__N_2506[90]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[114])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i90.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i91 (.D(dout_r_23__N_2506[91]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[115])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i91.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i92 (.D(dout_r_23__N_2506[92]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[116])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i92.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i93 (.D(dout_r_23__N_2506[93]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[117])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i93.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i94 (.D(dout_r_23__N_2506[94]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[118])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i94.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i95 (.D(dout_r_23__N_2506[95]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[119])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i95.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i96 (.D(dout_r_23__N_2506[96]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[120])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i96.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i97 (.D(dout_r_23__N_2506[97]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[121])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i97.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i98 (.D(dout_r_23__N_2506[98]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[122])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i98.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i99 (.D(dout_r_23__N_2506[99]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[123])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i99.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i100 (.D(dout_r_23__N_2506[100]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[124])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i100.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i101 (.D(dout_r_23__N_2506[101]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[125])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i101.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i102 (.D(dout_r_23__N_2506[102]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[126])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i102.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i103 (.D(dout_r_23__N_2506[103]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[127])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i103.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i104 (.D(dout_r_23__N_2506[104]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[128])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i104.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i105 (.D(dout_r_23__N_2506[105]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[129])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i105.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i106 (.D(dout_r_23__N_2506[106]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[130])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i106.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i107 (.D(dout_r_23__N_2506[107]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[131])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i107.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i108 (.D(dout_r_23__N_2506[108]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[132])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i108.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i109 (.D(dout_r_23__N_2506[109]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[133])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i109.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i110 (.D(dout_r_23__N_2506[110]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[134])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i110.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i111 (.D(dout_r_23__N_2506[111]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[135])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i111.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i112 (.D(dout_r_23__N_2506[112]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[136])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i112.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i113 (.D(dout_r_23__N_2506[113]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[137])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i113.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i114 (.D(dout_r_23__N_2506[114]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[138])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i114.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i115 (.D(dout_r_23__N_2506[115]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[139])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i115.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i116 (.D(dout_r_23__N_2506[116]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[140])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i116.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i117 (.D(dout_r_23__N_2506[117]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[141])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i117.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i118 (.D(dout_r_23__N_2506[118]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[142])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i118.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i119 (.D(dout_r_23__N_2506[119]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[143])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i119.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i120 (.D(dout_r_23__N_2506[120]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[144])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i120.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i121 (.D(dout_r_23__N_2506[121]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[145])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i121.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i122 (.D(dout_r_23__N_2506[122]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[146])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i122.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i123 (.D(dout_r_23__N_2506[123]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[147])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i123.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i124 (.D(dout_r_23__N_2506[124]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[148])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i124.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i125 (.D(dout_r_23__N_2506[125]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[149])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i125.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i126 (.D(dout_r_23__N_2506[126]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[150])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i126.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i127 (.D(dout_r_23__N_2506[127]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[151])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i127.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i128 (.D(dout_r_23__N_2506[128]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[152])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i128.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i129 (.D(dout_r_23__N_2506[129]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[153])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i129.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i130 (.D(dout_r_23__N_2506[130]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[154])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i130.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i131 (.D(dout_r_23__N_2506[131]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[155])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i131.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i132 (.D(dout_r_23__N_2506[132]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[156])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i132.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i133 (.D(dout_r_23__N_2506[133]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[157])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i133.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i134 (.D(dout_r_23__N_2506[134]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[158])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i134.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i135 (.D(dout_r_23__N_2506[135]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[159])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i135.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i136 (.D(dout_r_23__N_2506[136]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[160])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i136.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i137 (.D(dout_r_23__N_2506[137]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[161])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i137.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i138 (.D(dout_r_23__N_2506[138]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[162])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i138.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i139 (.D(dout_r_23__N_2506[139]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[163])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i139.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i140 (.D(dout_r_23__N_2506[140]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[164])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i140.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i141 (.D(dout_r_23__N_2506[141]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[165])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i141.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i142 (.D(dout_r_23__N_2506[142]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[166])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i142.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i143 (.D(dout_r_23__N_2506[143]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[167])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i143.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i144 (.D(dout_r_23__N_2506[144]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[168])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i144.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i145 (.D(dout_r_23__N_2506[145]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[169])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i145.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i146 (.D(dout_r_23__N_2506[146]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[170])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i146.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i147 (.D(dout_r_23__N_2506[147]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[171])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i147.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i148 (.D(dout_r_23__N_2506[148]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[172])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i148.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i149 (.D(dout_r_23__N_2506[149]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[173])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i149.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i150 (.D(dout_r_23__N_2506[150]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[174])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i150.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i151 (.D(dout_r_23__N_2506[151]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[175])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i151.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i152 (.D(dout_r_23__N_2506[152]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[176])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i152.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i153 (.D(dout_r_23__N_2506[153]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[177])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i153.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i154 (.D(dout_r_23__N_2506[154]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[178])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i154.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i155 (.D(dout_r_23__N_2506[155]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[179])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i155.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i156 (.D(dout_r_23__N_2506[156]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[180])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i156.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i157 (.D(dout_r_23__N_2506[157]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[181])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i157.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i158 (.D(dout_r_23__N_2506[158]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[182])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i158.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i159 (.D(dout_r_23__N_2506[159]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[183])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i159.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i160 (.D(dout_r_23__N_2506[160]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[184])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i160.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i161 (.D(dout_r_23__N_2506[161]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[185])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i161.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i162 (.D(dout_r_23__N_2506[162]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[186])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i162.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i163 (.D(dout_r_23__N_2506[163]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[187])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i163.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i164 (.D(dout_r_23__N_2506[164]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[188])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i164.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i165 (.D(dout_r_23__N_2506[165]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[189])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i165.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i166 (.D(dout_r_23__N_2506[166]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[190])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i166.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i167 (.D(dout_r_23__N_2506[167]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[191])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i167.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i168 (.D(dout_r_23__N_2506[168]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[192])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i168.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i169 (.D(dout_r_23__N_2506[169]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[193])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i169.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i170 (.D(dout_r_23__N_2506[170]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[194])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i170.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i171 (.D(dout_r_23__N_2506[171]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[195])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i171.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i172 (.D(dout_r_23__N_2506[172]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[196])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i172.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i173 (.D(dout_r_23__N_2506[173]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[197])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i173.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i174 (.D(dout_r_23__N_2506[174]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[198])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i174.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i175 (.D(dout_r_23__N_2506[175]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[199])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i175.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i176 (.D(dout_r_23__N_2506[176]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[200])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i176.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i177 (.D(dout_r_23__N_2506[177]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[201])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i177.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i178 (.D(dout_r_23__N_2506[178]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[202])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i178.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i179 (.D(dout_r_23__N_2506[179]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[203])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i179.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i180 (.D(dout_r_23__N_2506[180]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[204])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i180.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i181 (.D(dout_r_23__N_2506[181]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[205])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i181.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i182 (.D(dout_r_23__N_2506[182]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[206])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i182.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i183 (.D(dout_r_23__N_2506[183]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[207])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i183.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i184 (.D(dout_r_23__N_2506[184]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[208])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i184.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i185 (.D(dout_r_23__N_2506[185]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[209])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i185.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i186 (.D(dout_r_23__N_2506[186]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[210])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i186.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i187 (.D(dout_r_23__N_2506[187]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[211])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i187.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i188 (.D(dout_r_23__N_2506[188]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[212])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i188.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i189 (.D(dout_r_23__N_2506[189]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[213])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i189.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i190 (.D(dout_r_23__N_2506[190]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[214])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i190.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i191 (.D(dout_r_23__N_2506[191]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[215])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i191.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i192 (.D(dout_r_23__N_2506[192]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[216])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i192.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i193 (.D(dout_r_23__N_2506[193]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[217])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i193.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i194 (.D(dout_r_23__N_2506[194]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[218])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i194.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i195 (.D(dout_r_23__N_2506[195]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[219])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i195.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i196 (.D(dout_r_23__N_2506[196]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[220])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i196.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i197 (.D(dout_r_23__N_2506[197]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[221])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i197.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i198 (.D(dout_r_23__N_2506[198]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[222])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i198.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i199 (.D(dout_r_23__N_2506[199]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[223])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i199.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i200 (.D(dout_r_23__N_2506[200]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[224])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i200.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i201 (.D(dout_r_23__N_2506[201]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[225])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i201.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i202 (.D(dout_r_23__N_2506[202]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[226])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i202.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i203 (.D(dout_r_23__N_2506[203]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[227])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i203.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i204 (.D(dout_r_23__N_2506[204]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[228])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i204.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i205 (.D(dout_r_23__N_2506[205]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[229])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i205.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i206 (.D(dout_r_23__N_2506[206]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[230])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i206.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i207 (.D(dout_r_23__N_2506[207]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[231])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i207.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i208 (.D(dout_r_23__N_2506[208]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[232])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i208.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i209 (.D(dout_r_23__N_2506[209]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[233])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i209.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i210 (.D(dout_r_23__N_2506[210]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[234])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i210.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i211 (.D(dout_r_23__N_2506[211]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[235])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i211.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i212 (.D(dout_r_23__N_2506[212]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[236])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i212.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i213 (.D(dout_r_23__N_2506[213]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[237])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i213.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i214 (.D(dout_r_23__N_2506[214]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[238])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i214.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i215 (.D(dout_r_23__N_2506[215]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[239])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i215.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i216 (.D(dout_r_23__N_2506[216]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[240])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i216.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i217 (.D(dout_r_23__N_2506[217]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[241])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i217.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i218 (.D(dout_r_23__N_2506[218]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[242])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i218.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i219 (.D(dout_r_23__N_2506[219]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[243])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i219.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i220 (.D(dout_r_23__N_2506[220]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[244])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i220.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i221 (.D(dout_r_23__N_2506[221]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[245])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i221.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i222 (.D(dout_r_23__N_2506[222]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[246])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i222.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i223 (.D(dout_r_23__N_2506[223]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[247])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i223.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i224 (.D(dout_r_23__N_2506[224]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[248])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i224.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i225 (.D(dout_r_23__N_2506[225]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[249])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i225.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i226 (.D(dout_r_23__N_2506[226]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[250])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i226.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i227 (.D(dout_r_23__N_2506[227]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[251])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i227.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i228 (.D(dout_r_23__N_2506[228]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[252])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i228.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i229 (.D(dout_r_23__N_2506[229]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[253])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i229.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i230 (.D(dout_r_23__N_2506[230]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[254])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i230.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i231 (.D(dout_r_23__N_2506[231]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[255])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i231.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i232 (.D(dout_r_23__N_2506[232]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[256])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i232.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i233 (.D(dout_r_23__N_2506[233]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[257])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i233.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i234 (.D(dout_r_23__N_2506[234]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[258])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i234.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i235 (.D(dout_r_23__N_2506[235]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[259])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i235.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i236 (.D(dout_r_23__N_2506[236]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[260])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i236.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i237 (.D(dout_r_23__N_2506[237]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[261])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i237.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i238 (.D(dout_r_23__N_2506[238]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[262])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i238.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i239 (.D(dout_r_23__N_2506[239]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[263])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i239.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i240 (.D(dout_r_23__N_2506[240]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[264])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i240.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i241 (.D(dout_r_23__N_2506[241]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[265])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i241.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i242 (.D(dout_r_23__N_2506[242]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[266])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i242.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i243 (.D(dout_r_23__N_2506[243]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[267])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i243.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i244 (.D(dout_r_23__N_2506[244]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[268])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i244.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i245 (.D(dout_r_23__N_2506[245]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[269])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i245.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i246 (.D(dout_r_23__N_2506[246]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[270])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i246.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i247 (.D(dout_r_23__N_2506[247]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[271])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i247.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i248 (.D(dout_r_23__N_2506[248]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[272])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i248.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i249 (.D(dout_r_23__N_2506[249]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[273])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i249.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i250 (.D(dout_r_23__N_2506[250]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[274])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i250.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i251 (.D(dout_r_23__N_2506[251]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[275])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i251.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i252 (.D(dout_r_23__N_2506[252]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[276])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i252.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i253 (.D(dout_r_23__N_2506[253]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[277])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i253.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i254 (.D(dout_r_23__N_2506[254]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[278])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i254.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i255 (.D(dout_r_23__N_2506[255]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[279])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i255.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i256 (.D(dout_r_23__N_2506[256]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[280])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i256.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i257 (.D(dout_r_23__N_2506[257]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[281])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i257.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i258 (.D(dout_r_23__N_2506[258]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[282])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i258.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i259 (.D(dout_r_23__N_2506[259]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[283])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i259.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i260 (.D(dout_r_23__N_2506[260]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[284])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i260.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i261 (.D(dout_r_23__N_2506[261]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[285])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i261.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i262 (.D(dout_r_23__N_2506[262]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[286])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i262.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i263 (.D(dout_r_23__N_2506[263]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[287])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i263.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i264 (.D(dout_r_23__N_2506[264]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[288])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i264.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i265 (.D(dout_r_23__N_2506[265]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[289])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i265.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i266 (.D(dout_r_23__N_2506[266]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[290])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i266.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i267 (.D(dout_r_23__N_2506[267]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[291])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i267.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i268 (.D(dout_r_23__N_2506[268]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[292])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i268.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i269 (.D(dout_r_23__N_2506[269]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[293])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i269.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i270 (.D(dout_r_23__N_2506[270]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[294])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i270.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i271 (.D(dout_r_23__N_2506[271]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[295])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i271.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i272 (.D(dout_r_23__N_2506[272]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[296])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i272.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i273 (.D(dout_r_23__N_2506[273]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[297])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i273.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i274 (.D(dout_r_23__N_2506[274]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[298])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i274.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i275 (.D(dout_r_23__N_2506[275]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[299])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i275.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i276 (.D(dout_r_23__N_2506[276]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[300])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i276.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i277 (.D(dout_r_23__N_2506[277]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[301])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i277.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i278 (.D(dout_r_23__N_2506[278]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[302])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i278.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i279 (.D(dout_r_23__N_2506[279]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[303])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i279.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i280 (.D(dout_r_23__N_2506[280]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[304])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i280.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i281 (.D(dout_r_23__N_2506[281]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[305])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i281.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i282 (.D(dout_r_23__N_2506[282]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[306])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i282.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i283 (.D(dout_r_23__N_2506[283]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[307])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i283.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i284 (.D(dout_r_23__N_2506[284]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[308])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i284.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i285 (.D(dout_r_23__N_2506[285]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[309])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i285.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i286 (.D(dout_r_23__N_2506[286]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[310])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i286.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i287 (.D(dout_r_23__N_2506[287]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[311])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i287.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i288 (.D(dout_r_23__N_2506[288]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[312])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i288.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i289 (.D(dout_r_23__N_2506[289]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[313])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i289.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i290 (.D(dout_r_23__N_2506[290]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[314])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i290.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i291 (.D(dout_r_23__N_2506[291]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[315])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i291.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i292 (.D(dout_r_23__N_2506[292]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[316])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i292.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i293 (.D(dout_r_23__N_2506[293]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[317])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i293.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i294 (.D(dout_r_23__N_2506[294]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[318])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i294.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i295 (.D(dout_r_23__N_2506[295]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[319])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i295.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i296 (.D(dout_r_23__N_2506[296]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[320])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i296.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i297 (.D(dout_r_23__N_2506[297]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[321])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i297.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i298 (.D(dout_r_23__N_2506[298]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[322])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i298.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i299 (.D(dout_r_23__N_2506[299]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[323])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i299.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i300 (.D(dout_r_23__N_2506[300]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[324])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i300.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i301 (.D(dout_r_23__N_2506[301]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[325])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i301.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i302 (.D(dout_r_23__N_2506[302]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[326])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i302.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i303 (.D(dout_r_23__N_2506[303]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[327])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i303.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i304 (.D(dout_r_23__N_2506[304]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[328])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i304.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i305 (.D(dout_r_23__N_2506[305]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[329])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i305.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i306 (.D(dout_r_23__N_2506[306]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[330])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i306.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i307 (.D(dout_r_23__N_2506[307]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[331])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i307.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i308 (.D(dout_r_23__N_2506[308]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[332])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i308.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i309 (.D(dout_r_23__N_2506[309]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[333])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i309.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i310 (.D(dout_r_23__N_2506[310]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[334])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i310.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i311 (.D(dout_r_23__N_2506[311]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[335])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i311.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i312 (.D(dout_r_23__N_2506[312]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[336])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i312.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i313 (.D(dout_r_23__N_2506[313]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[337])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i313.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i314 (.D(dout_r_23__N_2506[314]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[338])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i314.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i315 (.D(dout_r_23__N_2506[315]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[339])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i315.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i316 (.D(dout_r_23__N_2506[316]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[340])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i316.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i317 (.D(dout_r_23__N_2506[317]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[341])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i317.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i318 (.D(dout_r_23__N_2506[318]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[342])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i318.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i319 (.D(dout_r_23__N_2506[319]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[343])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i319.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i320 (.D(dout_r_23__N_2506[320]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[344])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i320.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i321 (.D(dout_r_23__N_2506[321]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[345])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i321.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i322 (.D(dout_r_23__N_2506[322]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[346])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i322.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i323 (.D(dout_r_23__N_2506[323]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[347])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i323.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i324 (.D(dout_r_23__N_2506[324]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[348])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i324.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i325 (.D(dout_r_23__N_2506[325]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[349])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i325.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i326 (.D(dout_r_23__N_2506[326]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[350])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i326.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i327 (.D(dout_r_23__N_2506[327]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[351])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i327.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i328 (.D(dout_r_23__N_2506[328]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[352])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i328.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i329 (.D(dout_r_23__N_2506[329]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[353])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i329.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i330 (.D(dout_r_23__N_2506[330]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[354])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i330.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i331 (.D(dout_r_23__N_2506[331]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[355])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i331.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i332 (.D(dout_r_23__N_2506[332]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[356])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i332.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i333 (.D(dout_r_23__N_2506[333]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[357])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i333.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i334 (.D(dout_r_23__N_2506[334]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[358])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i334.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i335 (.D(dout_r_23__N_2506[335]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[359])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i335.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i336 (.D(dout_r_23__N_2506[336]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[360])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i336.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i337 (.D(dout_r_23__N_2506[337]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[361])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i337.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i338 (.D(dout_r_23__N_2506[338]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[362])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i338.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i339 (.D(dout_r_23__N_2506[339]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[363])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i339.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i340 (.D(dout_r_23__N_2506[340]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[364])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i340.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i341 (.D(dout_r_23__N_2506[341]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[365])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i341.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i342 (.D(dout_r_23__N_2506[342]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[366])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i342.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i343 (.D(dout_r_23__N_2506[343]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[367])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i343.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i344 (.D(dout_r_23__N_2506[344]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[368])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i344.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i345 (.D(dout_r_23__N_2506[345]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[369])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i345.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i346 (.D(dout_r_23__N_2506[346]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[370])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i346.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i347 (.D(dout_r_23__N_2506[347]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[371])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i347.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i348 (.D(dout_r_23__N_2506[348]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[372])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i348.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i349 (.D(dout_r_23__N_2506[349]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[373])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i349.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i350 (.D(dout_r_23__N_2506[350]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[374])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i350.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i351 (.D(dout_r_23__N_2506[351]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[375])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i351.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i352 (.D(dout_r_23__N_2506[352]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[376])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i352.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i353 (.D(dout_r_23__N_2506[353]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[377])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i353.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i354 (.D(dout_r_23__N_2506[354]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[378])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i354.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i355 (.D(dout_r_23__N_2506[355]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[379])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i355.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i356 (.D(dout_r_23__N_2506[356]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[380])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i356.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i357 (.D(dout_r_23__N_2506[357]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[381])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i357.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i358 (.D(dout_r_23__N_2506[358]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[382])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i358.GSR = "ENABLED";
    FD1P3AX shift_reg_r_i0_i359 (.D(dout_r_23__N_2506[359]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_r_23__N_2506[383])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i359.GSR = "ENABLED";
    LUT4 i153_2_lut_rep_413 (.A(valid), .B(in_valid_reg), .Z(clk_c_enable_1772)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i153_2_lut_rep_413.init = 16'heeee;
    LUT4 i12209_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[383]), 
         .D(\shift_16_dout_i[23] ), .Z(n29919)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12209_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12210_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[382]), 
         .D(\shift_16_dout_i[22] ), .Z(n29920)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12210_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12211_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[381]), 
         .D(\shift_16_dout_i[21] ), .Z(n29921)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12211_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12212_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[380]), 
         .D(\shift_16_dout_i[20] ), .Z(n29922)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12212_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12213_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[379]), 
         .D(\shift_16_dout_i[19] ), .Z(n29923)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12213_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12214_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[378]), 
         .D(\shift_16_dout_i[18] ), .Z(n29924)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12214_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12215_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[377]), 
         .D(\shift_16_dout_i[17] ), .Z(n29925)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12215_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12216_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[376]), 
         .D(\shift_16_dout_i[16] ), .Z(n29926)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12216_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12217_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[375]), 
         .D(\shift_16_dout_i[15] ), .Z(n29927)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12217_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12218_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[374]), 
         .D(\shift_16_dout_i[14] ), .Z(n29928)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12218_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12219_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[373]), 
         .D(\shift_16_dout_i[13] ), .Z(n29929)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12219_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12220_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[372]), 
         .D(\shift_16_dout_i[12] ), .Z(n29930)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12220_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12221_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[371]), 
         .D(\shift_16_dout_i[11] ), .Z(n29931)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12221_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12222_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[370]), 
         .D(\shift_16_dout_i[10] ), .Z(n29932)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12222_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12223_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[369]), 
         .D(\shift_16_dout_i[9] ), .Z(n29933)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12223_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12224_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[368]), 
         .D(\shift_16_dout_i[8] ), .Z(n29934)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12224_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12225_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[367]), 
         .D(\op_i_23__N_1154[7] ), .Z(n29935)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12225_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12226_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[366]), 
         .D(\op_i_23__N_1154[6] ), .Z(n29936)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12226_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12227_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[365]), 
         .D(\op_i_23__N_1154[5] ), .Z(n29937)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12227_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12228_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[364]), 
         .D(\op_i_23__N_1154[4] ), .Z(n29938)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12228_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12229_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[363]), 
         .D(\op_i_23__N_1154[3] ), .Z(n29939)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12229_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12230_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[362]), 
         .D(\op_i_23__N_1154[2] ), .Z(n29940)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12230_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12231_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[361]), 
         .D(\op_i_23__N_1154[1] ), .Z(n29941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12231_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12232_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_i_23__N_3274[360]), 
         .D(\op_i_23__N_1154[0] ), .Z(n29942)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12232_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12233_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[383]), 
         .D(\shift_16_dout_r[23] ), .Z(n29943)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12233_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12234_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[382]), 
         .D(\shift_16_dout_r[22] ), .Z(n29944)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12234_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12235_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[381]), 
         .D(\shift_16_dout_r[21] ), .Z(n29945)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12235_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12236_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[380]), 
         .D(\shift_16_dout_r[20] ), .Z(n29946)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12236_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12237_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[379]), 
         .D(\shift_16_dout_r[19] ), .Z(n29947)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12237_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12238_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[378]), 
         .D(\shift_16_dout_r[18] ), .Z(n29948)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12238_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12239_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[377]), 
         .D(\shift_16_dout_r[17] ), .Z(n29949)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12239_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12240_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[376]), 
         .D(\shift_16_dout_r[16] ), .Z(n29950)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12240_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12241_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[375]), 
         .D(\shift_16_dout_r[15] ), .Z(n29951)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12241_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12243_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[373]), 
         .D(\shift_16_dout_r[13] ), .Z(n29953)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12243_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12244_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[372]), 
         .D(\shift_16_dout_r[12] ), .Z(n29954)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12244_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12245_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[371]), 
         .D(\shift_16_dout_r[11] ), .Z(n29955)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12245_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12246_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[370]), 
         .D(\shift_16_dout_r[10] ), .Z(n29956)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12246_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12247_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[369]), 
         .D(\shift_16_dout_r[9] ), .Z(n29957)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12247_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12248_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[368]), 
         .D(\shift_16_dout_r[8] ), .Z(n29958)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12248_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12249_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[367]), 
         .D(\op_r_23__N_1106[7] ), .Z(n29959)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12249_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12250_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[366]), 
         .D(\op_r_23__N_1106[6] ), .Z(n29960)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12250_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12242_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[374]), 
         .D(\shift_16_dout_r[14] ), .Z(n29952)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12242_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12251_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[365]), 
         .D(\op_r_23__N_1106[5] ), .Z(n29961)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12251_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12252_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[364]), 
         .D(\op_r_23__N_1106[4] ), .Z(n29962)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12252_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12253_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[363]), 
         .D(\op_r_23__N_1106[3] ), .Z(n29963)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12253_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12254_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[362]), 
         .D(\op_r_23__N_1106[2] ), .Z(n29964)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12254_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12255_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[361]), 
         .D(\op_r_23__N_1106[1] ), .Z(n29965)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12255_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12256_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(dout_r_23__N_2506[360]), 
         .D(\op_r_23__N_1106[0] ), .Z(n29966)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12256_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12125_2_lut_3_lut_4_lut (.A(valid), .B(in_valid_reg), .C(\count[5] ), 
         .D(\count[4] ), .Z(n29834)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(42[10] 47[8])
    defparam i12125_2_lut_3_lut_4_lut.init = 16'he0ee;
    FD1P3AX shift_reg_i_i0_i8 (.D(\dout_i_23__N_3274[8] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i8.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i9 (.D(\dout_i_23__N_3274[9] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i9.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i10 (.D(\dout_i_23__N_3274[10] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i10.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i11 (.D(\dout_i_23__N_3274[11] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i11.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i12 (.D(\dout_i_23__N_3274[12] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i12.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i13 (.D(\dout_i_23__N_3274[13] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i13.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i14 (.D(\dout_i_23__N_3274[14] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i14.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i15 (.D(\dout_i_23__N_3274[15] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i15.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i16 (.D(\dout_i_23__N_3274[16] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i16.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i17 (.D(\dout_i_23__N_3274[17] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i17.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i18 (.D(\dout_i_23__N_3274[18] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i18.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i19 (.D(\dout_i_23__N_3274[19] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i19.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i20 (.D(\dout_i_23__N_3274[20] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i20.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i21 (.D(\dout_i_23__N_3274[21] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i21.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i22 (.D(\dout_i_23__N_3274[22] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i22.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i23 (.D(\dout_i_23__N_3274[23] ), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i23.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i24 (.D(dout_i_23__N_3274[24]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i24.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i25 (.D(dout_i_23__N_3274[25]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i25.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i26 (.D(dout_i_23__N_3274[26]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i26.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i27 (.D(dout_i_23__N_3274[27]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i27.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i28 (.D(dout_i_23__N_3274[28]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i28.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i29 (.D(dout_i_23__N_3274[29]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i29.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i30 (.D(dout_i_23__N_3274[30]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i30.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i31 (.D(dout_i_23__N_3274[31]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i31.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i32 (.D(dout_i_23__N_3274[32]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i32.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i33 (.D(dout_i_23__N_3274[33]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i33.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i34 (.D(dout_i_23__N_3274[34]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i34.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i35 (.D(dout_i_23__N_3274[35]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i35.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i36 (.D(dout_i_23__N_3274[36]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i36.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i37 (.D(dout_i_23__N_3274[37]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i37.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i38 (.D(dout_i_23__N_3274[38]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i38.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i39 (.D(dout_i_23__N_3274[39]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i39.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i40 (.D(dout_i_23__N_3274[40]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i40.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i41 (.D(dout_i_23__N_3274[41]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i41.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i42 (.D(dout_i_23__N_3274[42]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i42.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i43 (.D(dout_i_23__N_3274[43]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i43.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i44 (.D(dout_i_23__N_3274[44]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i44.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i45 (.D(dout_i_23__N_3274[45]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i45.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i46 (.D(dout_i_23__N_3274[46]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i46.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i47 (.D(dout_i_23__N_3274[47]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i47.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i48 (.D(dout_i_23__N_3274[48]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i48.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i49 (.D(dout_i_23__N_3274[49]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i49.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i50 (.D(dout_i_23__N_3274[50]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i50.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i51 (.D(dout_i_23__N_3274[51]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i51.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i52 (.D(dout_i_23__N_3274[52]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i52.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i53 (.D(dout_i_23__N_3274[53]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[77])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i53.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i54 (.D(dout_i_23__N_3274[54]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[78])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i54.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i55 (.D(dout_i_23__N_3274[55]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[79])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i55.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i56 (.D(dout_i_23__N_3274[56]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i56.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i57 (.D(dout_i_23__N_3274[57]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i57.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i58 (.D(dout_i_23__N_3274[58]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i58.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i59 (.D(dout_i_23__N_3274[59]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i59.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i60 (.D(dout_i_23__N_3274[60]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i60.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i61 (.D(dout_i_23__N_3274[61]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[85])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i61.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i62 (.D(dout_i_23__N_3274[62]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[86])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i62.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i63 (.D(dout_i_23__N_3274[63]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[87])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i63.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i64 (.D(dout_i_23__N_3274[64]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i64.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i65 (.D(dout_i_23__N_3274[65]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i65.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i66 (.D(dout_i_23__N_3274[66]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i66.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i67 (.D(dout_i_23__N_3274[67]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i67.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i68 (.D(dout_i_23__N_3274[68]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i68.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i69 (.D(dout_i_23__N_3274[69]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[93])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i69.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i70 (.D(dout_i_23__N_3274[70]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[94])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i70.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i71 (.D(dout_i_23__N_3274[71]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[95])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i71.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i72 (.D(dout_i_23__N_3274[72]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[96])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i72.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i73 (.D(dout_i_23__N_3274[73]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[97])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i73.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i74 (.D(dout_i_23__N_3274[74]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[98])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i74.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i75 (.D(dout_i_23__N_3274[75]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[99])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i75.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i76 (.D(dout_i_23__N_3274[76]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[100])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i76.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i77 (.D(dout_i_23__N_3274[77]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[101])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i77.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i78 (.D(dout_i_23__N_3274[78]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[102])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i78.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i79 (.D(dout_i_23__N_3274[79]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[103])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i79.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i80 (.D(dout_i_23__N_3274[80]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[104])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i80.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i81 (.D(dout_i_23__N_3274[81]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[105])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i81.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i82 (.D(dout_i_23__N_3274[82]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[106])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i82.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i83 (.D(dout_i_23__N_3274[83]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[107])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i83.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i84 (.D(dout_i_23__N_3274[84]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[108])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i84.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i85 (.D(dout_i_23__N_3274[85]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[109])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i85.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i86 (.D(dout_i_23__N_3274[86]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[110])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i86.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i87 (.D(dout_i_23__N_3274[87]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[111])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i87.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i88 (.D(dout_i_23__N_3274[88]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[112])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i88.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i89 (.D(dout_i_23__N_3274[89]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[113])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i89.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i90 (.D(dout_i_23__N_3274[90]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[114])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i90.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i91 (.D(dout_i_23__N_3274[91]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[115])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i91.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i92 (.D(dout_i_23__N_3274[92]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[116])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i92.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i93 (.D(dout_i_23__N_3274[93]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[117])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i93.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i94 (.D(dout_i_23__N_3274[94]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[118])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i94.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i95 (.D(dout_i_23__N_3274[95]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[119])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i95.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i96 (.D(dout_i_23__N_3274[96]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[120])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i96.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i97 (.D(dout_i_23__N_3274[97]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[121])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i97.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i98 (.D(dout_i_23__N_3274[98]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[122])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i98.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i99 (.D(dout_i_23__N_3274[99]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[123])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i99.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i100 (.D(dout_i_23__N_3274[100]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[124])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i100.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i101 (.D(dout_i_23__N_3274[101]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[125])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i101.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i102 (.D(dout_i_23__N_3274[102]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[126])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i102.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i103 (.D(dout_i_23__N_3274[103]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[127])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i103.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i104 (.D(dout_i_23__N_3274[104]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[128])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i104.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i105 (.D(dout_i_23__N_3274[105]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[129])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i105.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i106 (.D(dout_i_23__N_3274[106]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[130])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i106.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i107 (.D(dout_i_23__N_3274[107]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[131])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i107.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i108 (.D(dout_i_23__N_3274[108]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[132])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i108.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i109 (.D(dout_i_23__N_3274[109]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[133])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i109.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i110 (.D(dout_i_23__N_3274[110]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[134])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i110.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i111 (.D(dout_i_23__N_3274[111]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[135])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i111.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i112 (.D(dout_i_23__N_3274[112]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[136])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i112.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i113 (.D(dout_i_23__N_3274[113]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[137])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i113.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i114 (.D(dout_i_23__N_3274[114]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[138])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i114.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i115 (.D(dout_i_23__N_3274[115]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[139])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i115.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i116 (.D(dout_i_23__N_3274[116]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[140])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i116.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i117 (.D(dout_i_23__N_3274[117]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[141])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i117.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i118 (.D(dout_i_23__N_3274[118]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[142])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i118.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i119 (.D(dout_i_23__N_3274[119]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[143])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i119.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i120 (.D(dout_i_23__N_3274[120]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[144])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i120.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i121 (.D(dout_i_23__N_3274[121]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[145])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i121.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i122 (.D(dout_i_23__N_3274[122]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[146])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i122.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i123 (.D(dout_i_23__N_3274[123]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[147])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i123.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i124 (.D(dout_i_23__N_3274[124]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[148])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i124.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i125 (.D(dout_i_23__N_3274[125]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[149])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i125.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i126 (.D(dout_i_23__N_3274[126]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[150])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i126.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i127 (.D(dout_i_23__N_3274[127]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[151])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i127.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i128 (.D(dout_i_23__N_3274[128]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[152])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i128.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i129 (.D(dout_i_23__N_3274[129]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[153])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i129.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i130 (.D(dout_i_23__N_3274[130]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[154])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i130.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i131 (.D(dout_i_23__N_3274[131]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[155])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i131.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i132 (.D(dout_i_23__N_3274[132]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[156])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i132.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i133 (.D(dout_i_23__N_3274[133]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[157])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i133.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i134 (.D(dout_i_23__N_3274[134]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[158])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i134.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i135 (.D(dout_i_23__N_3274[135]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[159])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i135.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i136 (.D(dout_i_23__N_3274[136]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[160])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i136.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i137 (.D(dout_i_23__N_3274[137]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[161])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i137.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i138 (.D(dout_i_23__N_3274[138]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[162])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i138.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i139 (.D(dout_i_23__N_3274[139]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[163])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i139.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i140 (.D(dout_i_23__N_3274[140]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[164])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i140.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i141 (.D(dout_i_23__N_3274[141]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[165])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i141.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i142 (.D(dout_i_23__N_3274[142]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[166])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i142.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i143 (.D(dout_i_23__N_3274[143]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[167])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i143.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i144 (.D(dout_i_23__N_3274[144]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[168])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i144.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i145 (.D(dout_i_23__N_3274[145]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[169])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i145.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i146 (.D(dout_i_23__N_3274[146]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[170])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i146.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i147 (.D(dout_i_23__N_3274[147]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[171])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i147.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i148 (.D(dout_i_23__N_3274[148]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[172])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i148.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i149 (.D(dout_i_23__N_3274[149]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[173])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i149.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i150 (.D(dout_i_23__N_3274[150]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[174])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i150.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i151 (.D(dout_i_23__N_3274[151]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[175])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i151.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i152 (.D(dout_i_23__N_3274[152]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[176])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i152.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i153 (.D(dout_i_23__N_3274[153]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[177])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i153.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i154 (.D(dout_i_23__N_3274[154]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[178])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i154.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i155 (.D(dout_i_23__N_3274[155]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[179])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i155.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i156 (.D(dout_i_23__N_3274[156]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[180])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i156.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i157 (.D(dout_i_23__N_3274[157]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[181])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i157.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i158 (.D(dout_i_23__N_3274[158]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[182])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i158.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i159 (.D(dout_i_23__N_3274[159]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[183])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i159.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i160 (.D(dout_i_23__N_3274[160]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[184])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i160.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i161 (.D(dout_i_23__N_3274[161]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[185])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i161.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i162 (.D(dout_i_23__N_3274[162]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[186])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i162.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i163 (.D(dout_i_23__N_3274[163]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[187])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i163.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i164 (.D(dout_i_23__N_3274[164]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[188])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i164.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i165 (.D(dout_i_23__N_3274[165]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[189])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i165.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i166 (.D(dout_i_23__N_3274[166]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[190])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i166.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i167 (.D(dout_i_23__N_3274[167]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[191])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i167.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i168 (.D(dout_i_23__N_3274[168]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[192])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i168.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i169 (.D(dout_i_23__N_3274[169]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[193])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i169.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i170 (.D(dout_i_23__N_3274[170]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[194])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i170.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i171 (.D(dout_i_23__N_3274[171]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[195])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i171.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i172 (.D(dout_i_23__N_3274[172]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[196])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i172.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i173 (.D(dout_i_23__N_3274[173]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[197])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i173.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i174 (.D(dout_i_23__N_3274[174]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[198])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i174.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i175 (.D(dout_i_23__N_3274[175]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[199])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i175.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i176 (.D(dout_i_23__N_3274[176]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[200])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i176.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i177 (.D(dout_i_23__N_3274[177]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[201])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i177.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i178 (.D(dout_i_23__N_3274[178]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[202])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i178.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i179 (.D(dout_i_23__N_3274[179]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[203])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i179.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i180 (.D(dout_i_23__N_3274[180]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[204])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i180.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i181 (.D(dout_i_23__N_3274[181]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[205])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i181.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i182 (.D(dout_i_23__N_3274[182]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[206])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i182.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i183 (.D(dout_i_23__N_3274[183]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[207])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i183.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i184 (.D(dout_i_23__N_3274[184]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[208])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i184.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i185 (.D(dout_i_23__N_3274[185]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[209])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i185.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i186 (.D(dout_i_23__N_3274[186]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[210])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i186.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i187 (.D(dout_i_23__N_3274[187]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[211])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i187.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i188 (.D(dout_i_23__N_3274[188]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[212])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i188.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i189 (.D(dout_i_23__N_3274[189]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[213])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i189.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i190 (.D(dout_i_23__N_3274[190]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[214])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i190.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i191 (.D(dout_i_23__N_3274[191]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[215])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i191.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i192 (.D(dout_i_23__N_3274[192]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[216])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i192.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i193 (.D(dout_i_23__N_3274[193]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[217])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i193.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i194 (.D(dout_i_23__N_3274[194]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[218])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i194.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i195 (.D(dout_i_23__N_3274[195]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[219])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i195.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i196 (.D(dout_i_23__N_3274[196]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[220])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i196.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i197 (.D(dout_i_23__N_3274[197]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[221])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i197.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i198 (.D(dout_i_23__N_3274[198]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[222])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i198.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i199 (.D(dout_i_23__N_3274[199]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[223])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i199.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i200 (.D(dout_i_23__N_3274[200]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[224])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i200.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i201 (.D(dout_i_23__N_3274[201]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[225])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i201.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i202 (.D(dout_i_23__N_3274[202]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[226])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i202.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i203 (.D(dout_i_23__N_3274[203]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[227])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i203.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i204 (.D(dout_i_23__N_3274[204]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[228])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i204.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i205 (.D(dout_i_23__N_3274[205]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[229])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i205.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i206 (.D(dout_i_23__N_3274[206]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[230])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i206.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i207 (.D(dout_i_23__N_3274[207]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[231])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i207.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i208 (.D(dout_i_23__N_3274[208]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[232])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i208.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i209 (.D(dout_i_23__N_3274[209]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[233])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i209.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i210 (.D(dout_i_23__N_3274[210]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[234])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i210.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i211 (.D(dout_i_23__N_3274[211]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[235])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i211.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i212 (.D(dout_i_23__N_3274[212]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[236])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i212.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i213 (.D(dout_i_23__N_3274[213]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[237])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i213.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i214 (.D(dout_i_23__N_3274[214]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[238])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i214.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i215 (.D(dout_i_23__N_3274[215]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[239])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i215.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i216 (.D(dout_i_23__N_3274[216]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[240])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i216.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i217 (.D(dout_i_23__N_3274[217]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[241])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i217.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i218 (.D(dout_i_23__N_3274[218]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[242])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i218.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i219 (.D(dout_i_23__N_3274[219]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[243])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i219.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i220 (.D(dout_i_23__N_3274[220]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[244])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i220.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i221 (.D(dout_i_23__N_3274[221]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[245])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i221.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i222 (.D(dout_i_23__N_3274[222]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[246])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i222.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i223 (.D(dout_i_23__N_3274[223]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[247])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i223.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i224 (.D(dout_i_23__N_3274[224]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[248])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i224.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i225 (.D(dout_i_23__N_3274[225]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[249])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i225.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i226 (.D(dout_i_23__N_3274[226]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[250])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i226.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i227 (.D(dout_i_23__N_3274[227]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[251])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i227.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i228 (.D(dout_i_23__N_3274[228]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[252])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i228.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i229 (.D(dout_i_23__N_3274[229]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[253])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i229.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i230 (.D(dout_i_23__N_3274[230]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[254])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i230.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i231 (.D(dout_i_23__N_3274[231]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[255])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i231.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i232 (.D(dout_i_23__N_3274[232]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[256])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i232.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i233 (.D(dout_i_23__N_3274[233]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[257])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i233.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i234 (.D(dout_i_23__N_3274[234]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[258])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i234.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i235 (.D(dout_i_23__N_3274[235]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[259])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i235.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i236 (.D(dout_i_23__N_3274[236]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[260])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i236.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i237 (.D(dout_i_23__N_3274[237]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[261])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i237.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i238 (.D(dout_i_23__N_3274[238]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[262])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i238.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i239 (.D(dout_i_23__N_3274[239]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[263])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i239.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i240 (.D(dout_i_23__N_3274[240]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[264])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i240.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i241 (.D(dout_i_23__N_3274[241]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[265])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i241.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i242 (.D(dout_i_23__N_3274[242]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[266])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i242.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i243 (.D(dout_i_23__N_3274[243]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[267])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i243.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i244 (.D(dout_i_23__N_3274[244]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[268])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i244.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i245 (.D(dout_i_23__N_3274[245]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[269])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i245.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i246 (.D(dout_i_23__N_3274[246]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[270])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i246.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i247 (.D(dout_i_23__N_3274[247]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[271])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i247.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i248 (.D(dout_i_23__N_3274[248]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[272])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i248.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i249 (.D(dout_i_23__N_3274[249]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[273])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i249.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i250 (.D(dout_i_23__N_3274[250]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[274])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i250.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i251 (.D(dout_i_23__N_3274[251]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[275])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i251.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i252 (.D(dout_i_23__N_3274[252]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[276])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i252.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i253 (.D(dout_i_23__N_3274[253]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[277])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i253.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i254 (.D(dout_i_23__N_3274[254]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[278])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i254.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i255 (.D(dout_i_23__N_3274[255]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[279])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i255.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i256 (.D(dout_i_23__N_3274[256]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[280])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i256.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i257 (.D(dout_i_23__N_3274[257]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[281])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i257.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i258 (.D(dout_i_23__N_3274[258]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[282])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i258.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i259 (.D(dout_i_23__N_3274[259]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[283])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i259.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i260 (.D(dout_i_23__N_3274[260]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[284])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i260.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i261 (.D(dout_i_23__N_3274[261]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[285])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i261.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i262 (.D(dout_i_23__N_3274[262]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[286])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i262.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i263 (.D(dout_i_23__N_3274[263]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[287])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i263.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i264 (.D(dout_i_23__N_3274[264]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[288])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i264.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i265 (.D(dout_i_23__N_3274[265]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[289])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i265.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i266 (.D(dout_i_23__N_3274[266]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[290])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i266.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i267 (.D(dout_i_23__N_3274[267]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[291])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i267.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i268 (.D(dout_i_23__N_3274[268]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[292])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i268.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i269 (.D(dout_i_23__N_3274[269]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[293])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i269.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i270 (.D(dout_i_23__N_3274[270]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[294])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i270.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i271 (.D(dout_i_23__N_3274[271]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[295])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i271.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i272 (.D(dout_i_23__N_3274[272]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[296])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i272.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i273 (.D(dout_i_23__N_3274[273]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[297])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i273.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i274 (.D(dout_i_23__N_3274[274]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[298])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i274.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i275 (.D(dout_i_23__N_3274[275]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[299])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i275.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i276 (.D(dout_i_23__N_3274[276]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[300])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i276.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i277 (.D(dout_i_23__N_3274[277]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[301])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i277.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i278 (.D(dout_i_23__N_3274[278]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[302])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i278.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i279 (.D(dout_i_23__N_3274[279]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[303])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i279.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i280 (.D(dout_i_23__N_3274[280]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[304])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i280.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i281 (.D(dout_i_23__N_3274[281]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[305])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i281.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i282 (.D(dout_i_23__N_3274[282]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[306])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i282.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i283 (.D(dout_i_23__N_3274[283]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[307])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i283.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i284 (.D(dout_i_23__N_3274[284]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[308])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i284.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i285 (.D(dout_i_23__N_3274[285]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[309])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i285.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i286 (.D(dout_i_23__N_3274[286]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[310])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i286.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i287 (.D(dout_i_23__N_3274[287]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[311])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i287.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i288 (.D(dout_i_23__N_3274[288]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[312])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i288.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i289 (.D(dout_i_23__N_3274[289]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[313])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i289.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i290 (.D(dout_i_23__N_3274[290]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[314])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i290.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i291 (.D(dout_i_23__N_3274[291]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[315])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i291.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i292 (.D(dout_i_23__N_3274[292]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[316])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i292.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i293 (.D(dout_i_23__N_3274[293]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[317])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i293.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i294 (.D(dout_i_23__N_3274[294]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[318])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i294.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i295 (.D(dout_i_23__N_3274[295]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[319])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i295.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i296 (.D(dout_i_23__N_3274[296]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[320])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i296.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i297 (.D(dout_i_23__N_3274[297]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[321])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i297.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i298 (.D(dout_i_23__N_3274[298]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[322])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i298.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i299 (.D(dout_i_23__N_3274[299]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[323])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i299.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i300 (.D(dout_i_23__N_3274[300]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[324])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i300.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i301 (.D(dout_i_23__N_3274[301]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[325])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i301.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i302 (.D(dout_i_23__N_3274[302]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[326])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i302.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i303 (.D(dout_i_23__N_3274[303]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[327])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i303.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i304 (.D(dout_i_23__N_3274[304]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[328])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i304.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i305 (.D(dout_i_23__N_3274[305]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[329])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i305.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i306 (.D(dout_i_23__N_3274[306]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[330])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i306.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i307 (.D(dout_i_23__N_3274[307]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[331])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i307.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i308 (.D(dout_i_23__N_3274[308]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[332])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i308.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i309 (.D(dout_i_23__N_3274[309]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[333])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i309.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i310 (.D(dout_i_23__N_3274[310]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[334])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i310.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i311 (.D(dout_i_23__N_3274[311]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[335])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i311.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i312 (.D(dout_i_23__N_3274[312]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[336])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i312.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i313 (.D(dout_i_23__N_3274[313]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[337])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i313.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i314 (.D(dout_i_23__N_3274[314]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[338])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i314.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i315 (.D(dout_i_23__N_3274[315]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[339])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i315.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i316 (.D(dout_i_23__N_3274[316]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[340])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i316.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i317 (.D(dout_i_23__N_3274[317]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[341])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i317.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i318 (.D(dout_i_23__N_3274[318]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[342])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i318.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i319 (.D(dout_i_23__N_3274[319]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[343])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i319.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i320 (.D(dout_i_23__N_3274[320]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[344])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i320.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i321 (.D(dout_i_23__N_3274[321]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[345])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i321.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i322 (.D(dout_i_23__N_3274[322]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[346])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i322.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i323 (.D(dout_i_23__N_3274[323]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[347])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i323.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i324 (.D(dout_i_23__N_3274[324]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[348])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i324.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i325 (.D(dout_i_23__N_3274[325]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[349])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i325.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i326 (.D(dout_i_23__N_3274[326]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[350])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i326.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i327 (.D(dout_i_23__N_3274[327]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[351])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i327.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i328 (.D(dout_i_23__N_3274[328]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[352])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i328.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i329 (.D(dout_i_23__N_3274[329]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[353])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i329.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i330 (.D(dout_i_23__N_3274[330]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[354])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i330.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i331 (.D(dout_i_23__N_3274[331]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[355])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i331.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i332 (.D(dout_i_23__N_3274[332]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[356])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i332.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i333 (.D(dout_i_23__N_3274[333]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[357])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i333.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i334 (.D(dout_i_23__N_3274[334]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[358])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i334.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i335 (.D(dout_i_23__N_3274[335]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[359])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i335.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i336 (.D(dout_i_23__N_3274[336]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[360])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i336.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i337 (.D(dout_i_23__N_3274[337]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[361])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i337.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i338 (.D(dout_i_23__N_3274[338]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[362])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i338.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i339 (.D(dout_i_23__N_3274[339]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[363])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i339.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i340 (.D(dout_i_23__N_3274[340]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[364])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i340.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i341 (.D(dout_i_23__N_3274[341]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[365])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i341.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i342 (.D(dout_i_23__N_3274[342]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[366])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i342.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i343 (.D(dout_i_23__N_3274[343]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[367])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i343.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i344 (.D(dout_i_23__N_3274[344]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[368])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i344.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i345 (.D(dout_i_23__N_3274[345]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[369])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i345.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i346 (.D(dout_i_23__N_3274[346]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[370])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i346.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i347 (.D(dout_i_23__N_3274[347]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[371])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i347.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i348 (.D(dout_i_23__N_3274[348]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[372])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i348.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i349 (.D(dout_i_23__N_3274[349]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[373])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i349.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i350 (.D(dout_i_23__N_3274[350]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[374])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i350.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i351 (.D(dout_i_23__N_3274[351]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[375])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i351.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i352 (.D(dout_i_23__N_3274[352]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[376])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i352.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i353 (.D(dout_i_23__N_3274[353]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[377])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i353.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i354 (.D(dout_i_23__N_3274[354]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[378])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i354.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i355 (.D(dout_i_23__N_3274[355]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[379])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i355.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i356 (.D(dout_i_23__N_3274[356]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[380])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i356.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i357 (.D(dout_i_23__N_3274[357]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[381])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i357.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i358 (.D(dout_i_23__N_3274[358]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[382])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i358.GSR = "ENABLED";
    FD1P3AX shift_reg_i_i0_i359 (.D(dout_i_23__N_3274[359]), .SP(clk_c_enable_1772), 
            .CK(clk_c), .Q(dout_i_23__N_3274[383])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i359.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i360 (.D(n29966), .CK(clk_c), .Q(\op_r_23__N_1106[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i360.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i361 (.D(n29965), .CK(clk_c), .Q(\op_r_23__N_1106[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i361.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i362 (.D(n29964), .CK(clk_c), .Q(\op_r_23__N_1106[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i362.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i363 (.D(n29963), .CK(clk_c), .Q(\op_r_23__N_1106[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i363.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i364 (.D(n29962), .CK(clk_c), .Q(\op_r_23__N_1106[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i364.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i365 (.D(n29961), .CK(clk_c), .Q(\op_r_23__N_1106[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i365.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i366 (.D(n29960), .CK(clk_c), .Q(\op_r_23__N_1106[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i366.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i367 (.D(n29959), .CK(clk_c), .Q(\op_r_23__N_1106[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i367.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i368 (.D(n29958), .CK(clk_c), .Q(\shift_16_dout_r[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i368.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i369 (.D(n29957), .CK(clk_c), .Q(\shift_16_dout_r[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i369.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i370 (.D(n29956), .CK(clk_c), .Q(\shift_16_dout_r[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i370.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i371 (.D(n29955), .CK(clk_c), .Q(\shift_16_dout_r[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i371.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i372 (.D(n29954), .CK(clk_c), .Q(\shift_16_dout_r[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i372.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i373 (.D(n29953), .CK(clk_c), .Q(\shift_16_dout_r[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i373.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i374 (.D(n29952), .CK(clk_c), .Q(\shift_16_dout_r[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i374.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i375 (.D(n29951), .CK(clk_c), .Q(\shift_16_dout_r[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i375.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i376 (.D(n29950), .CK(clk_c), .Q(\shift_16_dout_r[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i376.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i377 (.D(n29949), .CK(clk_c), .Q(\shift_16_dout_r[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i377.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i378 (.D(n29948), .CK(clk_c), .Q(\shift_16_dout_r[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i378.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i379 (.D(n29947), .CK(clk_c), .Q(\shift_16_dout_r[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i379.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i380 (.D(n29946), .CK(clk_c), .Q(\shift_16_dout_r[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i380.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i381 (.D(n29945), .CK(clk_c), .Q(\shift_16_dout_r[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i381.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i382 (.D(n29944), .CK(clk_c), .Q(\shift_16_dout_r[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i382.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i383 (.D(n29943), .CK(clk_c), .Q(\shift_16_dout_r[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_r_i0_i383.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i360 (.D(n29942), .CK(clk_c), .Q(\op_i_23__N_1154[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i360.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i361 (.D(n29941), .CK(clk_c), .Q(\op_i_23__N_1154[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i361.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i362 (.D(n29940), .CK(clk_c), .Q(\op_i_23__N_1154[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i362.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i363 (.D(n29939), .CK(clk_c), .Q(\op_i_23__N_1154[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i363.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i364 (.D(n29938), .CK(clk_c), .Q(\op_i_23__N_1154[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i364.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i365 (.D(n29937), .CK(clk_c), .Q(\op_i_23__N_1154[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i365.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i366 (.D(n29936), .CK(clk_c), .Q(\op_i_23__N_1154[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i366.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i367 (.D(n29935), .CK(clk_c), .Q(\op_i_23__N_1154[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i367.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i368 (.D(n29934), .CK(clk_c), .Q(\shift_16_dout_i[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i368.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i369 (.D(n29933), .CK(clk_c), .Q(\shift_16_dout_i[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i369.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i370 (.D(n29932), .CK(clk_c), .Q(\shift_16_dout_i[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i370.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i371 (.D(n29931), .CK(clk_c), .Q(\shift_16_dout_i[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i371.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i372 (.D(n29930), .CK(clk_c), .Q(\shift_16_dout_i[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i372.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i373 (.D(n29929), .CK(clk_c), .Q(\shift_16_dout_i[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i373.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i374 (.D(n29928), .CK(clk_c), .Q(\shift_16_dout_i[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i374.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i375 (.D(n29927), .CK(clk_c), .Q(\shift_16_dout_i[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i375.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i376 (.D(n29926), .CK(clk_c), .Q(\shift_16_dout_i[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i376.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i377 (.D(n29925), .CK(clk_c), .Q(\shift_16_dout_i[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i377.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i378 (.D(n29924), .CK(clk_c), .Q(\shift_16_dout_i[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i378.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i379 (.D(n29923), .CK(clk_c), .Q(\shift_16_dout_i[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i379.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i380 (.D(n29922), .CK(clk_c), .Q(\shift_16_dout_i[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i380.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i381 (.D(n29921), .CK(clk_c), .Q(\shift_16_dout_i[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i381.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i382 (.D(n29920), .CK(clk_c), .Q(\shift_16_dout_i[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i382.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i383 (.D(n29919), .CK(clk_c), .Q(\shift_16_dout_i[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=97, LSE_RLINE=104 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_16.v(36[5] 47[8])
    defparam shift_reg_i_i0_i383.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module ROM_2
//

module ROM_2 (clk_c, clk_c_enable_2299, clk_c_enable_2300, n34839, n34801, 
            n34843, \s_count[1] , GND_net, VCC_net, \count[1] , n34800, 
            \state_1__N_5843[1] , n30179, valid, n34738, n34795, \rom2_w_r[8] , 
            n34769) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input clk_c_enable_2299;
    output clk_c_enable_2300;
    output n34839;
    output n34801;
    output n34843;
    output \s_count[1] ;
    input GND_net;
    input VCC_net;
    output \count[1] ;
    output n34800;
    output \state_1__N_5843[1] ;
    output n30179;
    input valid;
    output n34738;
    output n34795;
    output \rom2_w_r[8] ;
    output n34769;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    wire [5:0]n51;
    wire [5:0]n29;
    wire [1:0]s_count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(12[11:18])
    wire [1:0]n13;
    wire [5:0]count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(11[11:16])
    
    wire n32395, n32394, n32393;
    
    FD1P3AX count_696__i0 (.D(n29[0]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(n51[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i0.GSR = "ENABLED";
    FD1P3AX s_count_695__i0 (.D(n13[0]), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(s_count[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(33[24:35])
    defparam s_count_695__i0.GSR = "ENABLED";
    FD1P3AX count_696__i1_rep_443 (.D(n29[1]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(n34839)) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i1_rep_443.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_447 (.A(count[3]), .B(count[5]), .C(n34839), .D(n34801), 
         .Z(n34843)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i1_2_lut_rep_447.init = 16'hfffe;
    LUT4 i14028_2_lut (.A(\s_count[1] ), .B(s_count[0]), .Z(n13[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(33[24:35])
    defparam i14028_2_lut.init = 16'h6666;
    LUT4 i14026_1_lut (.A(s_count[0]), .Z(n13[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(33[24:35])
    defparam i14026_1_lut.init = 16'h5555;
    CCU2C count_696_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32395), .S0(n29[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696_add_4_7.INIT0 = 16'haaa0;
    defparam count_696_add_4_7.INIT1 = 16'h0000;
    defparam count_696_add_4_7.INJECT1_0 = "NO";
    defparam count_696_add_4_7.INJECT1_1 = "NO";
    CCU2C count_696_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32394), .COUT(n32395), .S0(n29[3]), .S1(n29[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696_add_4_5.INIT0 = 16'haaa0;
    defparam count_696_add_4_5.INIT1 = 16'haaa0;
    defparam count_696_add_4_5.INJECT1_0 = "NO";
    defparam count_696_add_4_5.INJECT1_1 = "NO";
    CCU2C count_696_add_4_3 (.A0(\count[1] ), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32393), .COUT(n32394), .S0(n29[1]), .S1(n29[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696_add_4_3.INIT0 = 16'haaa0;
    defparam count_696_add_4_3.INIT1 = 16'haaa0;
    defparam count_696_add_4_3.INJECT1_0 = "NO";
    defparam count_696_add_4_3.INJECT1_1 = "NO";
    CCU2C count_696_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n51[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32393), .S1(n29[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696_add_4_1.INIT0 = 16'h0000;
    defparam count_696_add_4_1.INIT1 = 16'h555f;
    defparam count_696_add_4_1.INJECT1_0 = "NO";
    defparam count_696_add_4_1.INJECT1_1 = "NO";
    LUT4 i14_2_lut_3_lut_4_lut (.A(n34801), .B(n34800), .C(\s_count[1] ), 
         .D(\count[1] ), .Z(\state_1__N_5843[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i14_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i12469_2_lut_3_lut_4_lut (.A(n34801), .B(n34800), .C(\s_count[1] ), 
         .D(n34839), .Z(n30179)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i12469_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i260_2_lut_rep_376_3_lut_4_lut (.A(n34801), .B(n34800), .C(valid), 
         .D(\count[1] ), .Z(n34738)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i260_2_lut_rep_376_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12545_2_lut_rep_433 (.A(s_count[0]), .B(\s_count[1] ), .Z(n34795)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12545_2_lut_rep_433.init = 16'h8888;
    LUT4 i12546_1_lut_2_lut (.A(s_count[0]), .B(\s_count[1] ), .Z(\rom2_w_r[8] )) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i12546_1_lut_2_lut.init = 16'h7777;
    LUT4 i1_2_lut_rep_438 (.A(count[3]), .B(count[5]), .Z(n34800)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i1_2_lut_rep_438.init = 16'heeee;
    LUT4 i1_2_lut_rep_388_3_lut_4_lut (.A(count[3]), .B(count[5]), .C(n34839), 
         .D(n34801), .Z(clk_c_enable_2300)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i1_2_lut_rep_388_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_439 (.A(count[4]), .B(count[2]), .Z(n34801)) /* synthesis lut_function=(A+(B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i1_2_lut_rep_439.init = 16'heeee;
    LUT4 i1_2_lut_rep_407_3_lut_4_lut (.A(count[4]), .B(count[2]), .C(count[5]), 
         .D(count[3]), .Z(n34769)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(26[9:19])
    defparam i1_2_lut_rep_407_3_lut_4_lut.init = 16'hfffe;
    FD1P3AX count_696__i1 (.D(n29[1]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(\count[1] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i1.GSR = "ENABLED";
    FD1P3AX count_696__i2 (.D(n29[2]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i2.GSR = "ENABLED";
    FD1P3AX count_696__i3 (.D(n29[3]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i3.GSR = "ENABLED";
    FD1P3AX count_696__i4 (.D(n29[4]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i4.GSR = "ENABLED";
    FD1P3AX count_696__i5 (.D(n29[5]), .SP(clk_c_enable_2299), .CK(clk_c), 
            .Q(count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(18[22:31])
    defparam count_696__i5.GSR = "ENABLED";
    FD1P3AX s_count_695__i1 (.D(n13[1]), .SP(clk_c_enable_2300), .CK(clk_c), 
            .Q(\s_count[1] ));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_2.v(33[24:35])
    defparam s_count_695__i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module shift_1
//

module shift_1 (rst_n_c, rst_n_N_2, valid, clk_c, n34738, n34843, 
            dout_i_23__N_5974, shift_1_dout_i, dout_r_23__N_5926, shift_1_dout_r) /* synthesis syn_module_defined=1 */ ;
    input rst_n_c;
    output rst_n_N_2;
    output valid;
    input clk_c;
    input n34738;
    input n34843;
    input [23:0]dout_i_23__N_5974;
    output [23:0]shift_1_dout_i;
    input [23:0]dout_r_23__N_5926;
    output [23:0]shift_1_dout_r;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    
    wire n29873, n29872, n29874, n29875, n29876, n29877, n29878, 
        n29879, n29880, n29881, n29882, n29883, n29884, n29885, 
        n29886, n29887, n29888, n29889, n29890, n29891, n29892, 
        n29893, n29894, n29895, n29896, n29897, n29898, n29899, 
        n29900, n29901, n29902, n29903, n29904, n29905, n29906, 
        n29907, n29908, n29909, n29910, n29911, n29912, n29913, 
        n29914, n29915, n29916, n29917, n29918, n29871;
    
    LUT4 rst_n_I_0_1_lut (.A(rst_n_c), .Z(rst_n_N_2)) /* synthesis lut_function=(!(A)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(265[8:14])
    defparam rst_n_I_0_1_lut.init = 16'h5555;
    FD1S3AX valid_26 (.D(n34738), .CK(clk_c), .Q(valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam valid_26.GSR = "ENABLED";
    LUT4 i12163_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[21]), 
         .D(shift_1_dout_i[21]), .Z(n29873)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12163_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12162_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[22]), 
         .D(shift_1_dout_i[22]), .Z(n29872)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12162_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12164_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[20]), 
         .D(shift_1_dout_i[20]), .Z(n29874)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12164_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12165_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[19]), 
         .D(shift_1_dout_i[19]), .Z(n29875)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12165_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12166_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[18]), 
         .D(shift_1_dout_i[18]), .Z(n29876)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12166_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12167_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[17]), 
         .D(shift_1_dout_i[17]), .Z(n29877)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12167_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12168_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[16]), 
         .D(shift_1_dout_i[16]), .Z(n29878)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12168_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12169_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[15]), 
         .D(shift_1_dout_i[15]), .Z(n29879)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12169_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12170_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[14]), 
         .D(shift_1_dout_i[14]), .Z(n29880)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12170_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12171_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[13]), 
         .D(shift_1_dout_i[13]), .Z(n29881)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12171_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12172_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[12]), 
         .D(shift_1_dout_i[12]), .Z(n29882)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12172_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12173_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[11]), 
         .D(shift_1_dout_i[11]), .Z(n29883)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12173_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12174_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[10]), 
         .D(shift_1_dout_i[10]), .Z(n29884)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12174_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12175_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[9]), 
         .D(shift_1_dout_i[9]), .Z(n29885)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12175_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12176_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[8]), 
         .D(shift_1_dout_i[8]), .Z(n29886)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12176_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12177_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[7]), 
         .D(shift_1_dout_i[7]), .Z(n29887)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12177_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12178_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[6]), 
         .D(shift_1_dout_i[6]), .Z(n29888)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12178_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12179_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[5]), 
         .D(shift_1_dout_i[5]), .Z(n29889)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12179_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12180_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[4]), 
         .D(shift_1_dout_i[4]), .Z(n29890)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12181_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[3]), 
         .D(shift_1_dout_i[3]), .Z(n29891)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12181_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12182_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[2]), 
         .D(shift_1_dout_i[2]), .Z(n29892)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12182_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12183_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[1]), 
         .D(shift_1_dout_i[1]), .Z(n29893)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12183_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12184_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[0]), 
         .D(shift_1_dout_i[0]), .Z(n29894)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12185_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[23]), 
         .D(shift_1_dout_r[23]), .Z(n29895)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12186_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[22]), 
         .D(shift_1_dout_r[22]), .Z(n29896)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12186_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12187_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[21]), 
         .D(shift_1_dout_r[21]), .Z(n29897)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12187_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12188_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[20]), 
         .D(shift_1_dout_r[20]), .Z(n29898)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12189_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[19]), 
         .D(shift_1_dout_r[19]), .Z(n29899)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12189_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12190_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[18]), 
         .D(shift_1_dout_r[18]), .Z(n29900)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12191_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[17]), 
         .D(shift_1_dout_r[17]), .Z(n29901)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12192_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[16]), 
         .D(shift_1_dout_r[16]), .Z(n29902)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12193_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[15]), 
         .D(shift_1_dout_r[15]), .Z(n29903)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12193_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12194_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[14]), 
         .D(shift_1_dout_r[14]), .Z(n29904)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12194_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12195_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[13]), 
         .D(shift_1_dout_r[13]), .Z(n29905)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12195_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12196_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[12]), 
         .D(shift_1_dout_r[12]), .Z(n29906)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12196_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12197_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[11]), 
         .D(shift_1_dout_r[11]), .Z(n29907)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12197_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12198_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[10]), 
         .D(shift_1_dout_r[10]), .Z(n29908)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12198_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12199_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[9]), 
         .D(shift_1_dout_r[9]), .Z(n29909)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12199_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12200_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[8]), 
         .D(shift_1_dout_r[8]), .Z(n29910)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12200_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12201_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[7]), 
         .D(shift_1_dout_r[7]), .Z(n29911)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12201_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12202_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[6]), 
         .D(shift_1_dout_r[6]), .Z(n29912)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12202_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12203_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[5]), 
         .D(shift_1_dout_r[5]), .Z(n29913)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12203_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12204_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[4]), 
         .D(shift_1_dout_r[4]), .Z(n29914)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12204_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12205_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[3]), 
         .D(shift_1_dout_r[3]), .Z(n29915)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12205_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12206_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[2]), 
         .D(shift_1_dout_r[2]), .Z(n29916)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12206_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12207_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[1]), 
         .D(shift_1_dout_r[1]), .Z(n29917)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12207_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12208_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_r_23__N_5926[0]), 
         .D(shift_1_dout_r[0]), .Z(n29918)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12208_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12161_3_lut_4_lut (.A(valid), .B(n34843), .C(dout_i_23__N_5974[23]), 
         .D(shift_1_dout_i[23]), .Z(n29871)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(41[14] 46[8])
    defparam i12161_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX shift_reg_r_i0_i0 (.D(n29918), .CK(clk_c), .Q(shift_1_dout_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i0.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i1 (.D(n29917), .CK(clk_c), .Q(shift_1_dout_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i1.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i2 (.D(n29916), .CK(clk_c), .Q(shift_1_dout_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i2.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i3 (.D(n29915), .CK(clk_c), .Q(shift_1_dout_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i3.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i4 (.D(n29914), .CK(clk_c), .Q(shift_1_dout_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i4.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i5 (.D(n29913), .CK(clk_c), .Q(shift_1_dout_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i5.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i6 (.D(n29912), .CK(clk_c), .Q(shift_1_dout_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i6.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i7 (.D(n29911), .CK(clk_c), .Q(shift_1_dout_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i7.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i8 (.D(n29910), .CK(clk_c), .Q(shift_1_dout_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i8.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i9 (.D(n29909), .CK(clk_c), .Q(shift_1_dout_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i9.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i10 (.D(n29908), .CK(clk_c), .Q(shift_1_dout_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i10.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i11 (.D(n29907), .CK(clk_c), .Q(shift_1_dout_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i11.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i12 (.D(n29906), .CK(clk_c), .Q(shift_1_dout_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i12.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i13 (.D(n29905), .CK(clk_c), .Q(shift_1_dout_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i13.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i14 (.D(n29904), .CK(clk_c), .Q(shift_1_dout_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i14.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i15 (.D(n29903), .CK(clk_c), .Q(shift_1_dout_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i15.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i16 (.D(n29902), .CK(clk_c), .Q(shift_1_dout_r[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i16.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i17 (.D(n29901), .CK(clk_c), .Q(shift_1_dout_r[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i17.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i18 (.D(n29900), .CK(clk_c), .Q(shift_1_dout_r[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i18.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i19 (.D(n29899), .CK(clk_c), .Q(shift_1_dout_r[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i19.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i20 (.D(n29898), .CK(clk_c), .Q(shift_1_dout_r[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i20.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i21 (.D(n29897), .CK(clk_c), .Q(shift_1_dout_r[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i21.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i22 (.D(n29896), .CK(clk_c), .Q(shift_1_dout_r[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i22.GSR = "ENABLED";
    FD1S3AX shift_reg_r_i0_i23 (.D(n29895), .CK(clk_c), .Q(shift_1_dout_r[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_r_i0_i23.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i0 (.D(n29894), .CK(clk_c), .Q(shift_1_dout_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i0.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i1 (.D(n29893), .CK(clk_c), .Q(shift_1_dout_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i1.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i2 (.D(n29892), .CK(clk_c), .Q(shift_1_dout_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i2.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i3 (.D(n29891), .CK(clk_c), .Q(shift_1_dout_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i3.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i4 (.D(n29890), .CK(clk_c), .Q(shift_1_dout_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i4.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i5 (.D(n29889), .CK(clk_c), .Q(shift_1_dout_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i5.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i6 (.D(n29888), .CK(clk_c), .Q(shift_1_dout_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i6.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i7 (.D(n29887), .CK(clk_c), .Q(shift_1_dout_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i7.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i8 (.D(n29886), .CK(clk_c), .Q(shift_1_dout_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i8.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i9 (.D(n29885), .CK(clk_c), .Q(shift_1_dout_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i9.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i10 (.D(n29884), .CK(clk_c), .Q(shift_1_dout_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i10.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i11 (.D(n29883), .CK(clk_c), .Q(shift_1_dout_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i11.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i12 (.D(n29882), .CK(clk_c), .Q(shift_1_dout_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i12.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i13 (.D(n29881), .CK(clk_c), .Q(shift_1_dout_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i13.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i14 (.D(n29880), .CK(clk_c), .Q(shift_1_dout_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i14.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i15 (.D(n29879), .CK(clk_c), .Q(shift_1_dout_i[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i15.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i16 (.D(n29878), .CK(clk_c), .Q(shift_1_dout_i[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i16.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i17 (.D(n29877), .CK(clk_c), .Q(shift_1_dout_i[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i17.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i18 (.D(n29876), .CK(clk_c), .Q(shift_1_dout_i[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i18.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i19 (.D(n29875), .CK(clk_c), .Q(shift_1_dout_i[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i19.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i20 (.D(n29874), .CK(clk_c), .Q(shift_1_dout_i[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i20.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i21 (.D(n29873), .CK(clk_c), .Q(shift_1_dout_i[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i21.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i22 (.D(n29872), .CK(clk_c), .Q(shift_1_dout_i[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i22.GSR = "ENABLED";
    FD1S3AX shift_reg_i_i0_i23 (.D(n29871), .CK(clk_c), .Q(shift_1_dout_i[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=232, LSE_RLINE=239 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/shift_1.v(36[5] 46[8])
    defparam shift_reg_i_i0_i23.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module ROM_4
//

module ROM_4 (n29820, n29819, n34520, \rom4_state[0] , state_1__N_5502, 
            clk_c, clk_c_enable_2305, s_count, \rom4_w_i[12] , GND_net, 
            VCC_net, n29826, n29828, n29827, n34841, \rom4_w_r[1] , 
            n34776, \rom4_w_r[8] , n34777, \rom4_w_r[5] , n34799, 
            clk_c_enable_2299, n6514, n3, n30041) /* synthesis syn_module_defined=1 */ ;
    output n29820;
    output n29819;
    output n34520;
    output \rom4_state[0] ;
    output state_1__N_5502;
    input clk_c;
    input clk_c_enable_2305;
    output [2:0]s_count;
    output \rom4_w_i[12] ;
    input GND_net;
    input VCC_net;
    output n29826;
    output n29828;
    output n29827;
    output n34841;
    output \rom4_w_r[1] ;
    output n34776;
    output \rom4_w_r[8] ;
    output n34777;
    output \rom4_w_r[5] ;
    output n34799;
    output clk_c_enable_2299;
    output n6514;
    output n3;
    input n30041;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/fft.v(13[7:10])
    wire [5:0]count;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(11[11:16])
    wire [5:0]n51;
    wire [5:0]n29;
    
    wire n32398, n32397, n32396, n30042;
    
    LUT4 i12111_3_lut (.A(n29820), .B(n29819), .C(n34520), .Z(\rom4_state[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(14[1] 57[4])
    defparam i12111_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(count[2]), .B(count[5]), .C(count[3]), .D(count[4]), 
         .Z(state_1__N_5502)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    FD1P3AX count_694__i0 (.D(n29[0]), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(n51[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694__i0.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(s_count[2]), .B(s_count[1]), .C(s_count[0]), .Z(\rom4_w_i[12] )) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_3_lut.init = 16'ha8a8;
    CCU2C count_694_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n32398), .S0(n29[5]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694_add_4_7.INIT0 = 16'haaa0;
    defparam count_694_add_4_7.INIT1 = 16'h0000;
    defparam count_694_add_4_7.INJECT1_0 = "NO";
    defparam count_694_add_4_7.INJECT1_1 = "NO";
    CCU2C count_694_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32397), .COUT(n32398), .S0(n29[3]), .S1(n29[4]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694_add_4_5.INIT0 = 16'haaa0;
    defparam count_694_add_4_5.INIT1 = 16'haaa0;
    defparam count_694_add_4_5.INJECT1_0 = "NO";
    defparam count_694_add_4_5.INJECT1_1 = "NO";
    CCU2C count_694_add_4_3 (.A0(n51[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n32396), .COUT(n32397), .S0(n29[1]), .S1(n29[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694_add_4_3.INIT0 = 16'haaa0;
    defparam count_694_add_4_3.INIT1 = 16'haaa0;
    defparam count_694_add_4_3.INJECT1_0 = "NO";
    defparam count_694_add_4_3.INJECT1_1 = "NO";
    CCU2C count_694_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n51[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n32396), .S1(n29[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694_add_4_1.INIT0 = 16'h0000;
    defparam count_694_add_4_1.INIT1 = 16'h555f;
    defparam count_694_add_4_1.INJECT1_0 = "NO";
    defparam count_694_add_4_1.INJECT1_1 = "NO";
    LUT4 i16387_3_lut_3_lut (.A(state_1__N_5502), .B(s_count[2]), .C(n29820), 
         .Z(n29820)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i16387_3_lut_3_lut.init = 16'h2020;
    LUT4 i16355_3_lut_2_lut (.A(state_1__N_5502), .B(s_count[2]), .Z(n34520)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i16355_3_lut_2_lut.init = 16'h2222;
    LUT4 i16391_3_lut_3_lut (.A(state_1__N_5502), .B(s_count[2]), .C(n29819), 
         .Z(n29819)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam i16391_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i16363_3_lut_2_lut (.A(s_count[2]), .B(state_1__N_5502), .Z(n29826)) /* synthesis lut_function=(A (B)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(27[10] 34[8])
    defparam i16363_3_lut_2_lut.init = 16'h8888;
    LUT4 i16371_3_lut_3_lut (.A(s_count[2]), .B(state_1__N_5502), .C(n29828), 
         .Z(n29828)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(27[10] 34[8])
    defparam i16371_3_lut_3_lut.init = 16'h8080;
    LUT4 i16375_4_lut_2_lut_3_lut (.A(s_count[2]), .B(state_1__N_5502), 
         .C(n29827), .Z(n29827)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(27[10] 34[8])
    defparam i16375_4_lut_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i2351_2_lut_rep_445 (.A(n29828), .B(n29827), .C(n29826), .D(\rom4_state[0] ), 
         .Z(n34841)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(14[1] 57[4])
    defparam i2351_2_lut_rep_445.init = 16'h35ca;
    LUT4 i1_2_lut_3_lut (.A(s_count[1]), .B(s_count[0]), .C(s_count[2]), 
         .Z(\rom4_w_r[1] )) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i12332_3_lut_4_lut (.A(s_count[1]), .B(s_count[0]), .C(state_1__N_5502), 
         .D(s_count[2]), .Z(n30042)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i12332_3_lut_4_lut.init = 16'h7f80;
    LUT4 i21_2_lut_rep_414 (.A(s_count[0]), .B(s_count[1]), .Z(n34776)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i21_2_lut_rep_414.init = 16'h6666;
    LUT4 i16324_2_lut_3_lut (.A(s_count[0]), .B(s_count[1]), .C(s_count[2]), 
         .Z(\rom4_w_r[8] )) /* synthesis lut_function=(A (B+!(C))+!A !(B (C))) */ ;
    defparam i16324_2_lut_3_lut.init = 16'h9f9f;
    LUT4 i1_2_lut_rep_415 (.A(s_count[2]), .B(s_count[0]), .Z(n34777)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_415.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_20 (.A(s_count[2]), .B(s_count[0]), .C(s_count[1]), 
         .Z(\rom4_w_r[5] )) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_20.init = 16'h0808;
    LUT4 i12119_3_lut_rep_437 (.A(n29828), .B(n29827), .C(n29826), .Z(n34799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(14[1] 57[4])
    defparam i12119_3_lut_rep_437.init = 16'hcaca;
    LUT4 i2351_2_lut_rep_406_4_lut (.A(n29828), .B(n29827), .C(n29826), 
         .D(\rom4_state[0] ), .Z(clk_c_enable_2299)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(14[1] 57[4])
    defparam i2351_2_lut_rep_406_4_lut.init = 16'h35ca;
    LUT4 i252_2_lut_4_lut (.A(n29828), .B(n29827), .C(n29826), .D(\rom4_state[0] ), 
         .Z(n6514)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(14[1] 57[4])
    defparam i252_2_lut_4_lut.init = 16'h00ca;
    LUT4 equal_374_i3_2_lut_4_lut (.A(n29828), .B(n29827), .C(n29826), 
         .D(\rom4_state[0] ), .Z(n3)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(14[1] 57[4])
    defparam equal_374_i3_2_lut_4_lut.init = 16'hcaff;
    FD1S3AX s_count_693__i2 (.D(n30042), .CK(clk_c), .Q(s_count[2]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(33[24:35])
    defparam s_count_693__i2.GSR = "ENABLED";
    FD1S3AX s_count_693__i0 (.D(n30041), .CK(clk_c), .Q(s_count[0]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(33[24:35])
    defparam s_count_693__i0.GSR = "ENABLED";
    FD1P3AX count_694__i1 (.D(n29[1]), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(n51[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694__i1.GSR = "ENABLED";
    FD1P3AX count_694__i2 (.D(n29[2]), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694__i2.GSR = "ENABLED";
    FD1P3AX count_694__i3 (.D(n29[3]), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694__i3.GSR = "ENABLED";
    FD1P3AX count_694__i4 (.D(n29[4]), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694__i4.GSR = "ENABLED";
    FD1P3AX count_694__i5 (.D(n29[5]), .SP(clk_c_enable_2305), .CK(clk_c), 
            .Q(count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(17[22:31])
    defparam count_694__i5.GSR = "ENABLED";
    FD1P3AX s_count_693__i1 (.D(n34776), .SP(state_1__N_5502), .CK(clk_c), 
            .Q(s_count[1]));   // d:/ci/rtl_fpga/sd4/fft/impl1/source/rom_4.v(33[24:35])
    defparam s_count_693__i1.GSR = "ENABLED";
    
endmodule
