module transistors (
	input a,
	output b
);

// and gate
not(b,a);

endmodule