// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Wed Jul 23 21:37:01 2025
//
// Verilog Description of module matrix_inv
//

module matrix_inv (clk, reset, a, b, c, d, a_inv, b_inv, c_inv, 
            d_inv, error) /* synthesis syn_module_defined=1 */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(8[8:18])
    input clk;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[20:23])
    input reset;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[25:30])
    input [15:0]a;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    input [15:0]b;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    input [15:0]c;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    input [15:0]d;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    output [15:0]a_inv;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    output [15:0]b_inv;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    output [15:0]c_inv;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    output [15:0]d_inv;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    output error;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(19[26:31])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[20:23])
    
    wire GND_net, VCC_net, reset_c, a_c_15, a_c_14, a_c_13, a_c_12, 
        a_c_11, a_c_10, a_c_9, a_c_8, a_c_7, a_c_6, a_c_5, a_c_4, 
        a_c_3, a_c_2, a_c_1, a_c_0, b_c_15, b_c_14, b_c_13, b_c_12, 
        b_c_11, b_c_10, b_c_9, b_c_8, b_c_7, b_c_6, b_c_5, b_c_4, 
        b_c_3, b_c_2, b_c_1, b_c_0, c_c_15, c_c_14, c_c_13, c_c_12, 
        c_c_11, c_c_10, c_c_9, c_c_8, c_c_7, c_c_6, c_c_5, c_c_4, 
        c_c_3, c_c_2, c_c_1, c_c_0, d_c_15, d_c_14, d_c_13, d_c_12, 
        d_c_11, d_c_10, d_c_9, d_c_8, d_c_7, d_c_6, d_c_5, d_c_4, 
        d_c_3, d_c_2, d_c_1, d_c_0, a_inv_c_15, a_inv_c_14, a_inv_c_13, 
        a_inv_c_12, a_inv_c_11, a_inv_c_10, a_inv_c_9, a_inv_c_8, 
        a_inv_c_7, a_inv_c_6, a_inv_c_5, a_inv_c_4, a_inv_c_3, a_inv_c_2, 
        a_inv_c_1, a_inv_c_0, b_inv_c_15, b_inv_c_14, b_inv_c_13, 
        b_inv_c_12, b_inv_c_11, b_inv_c_10, b_inv_c_9, b_inv_c_8, 
        b_inv_c_7, b_inv_c_6, b_inv_c_5, b_inv_c_4, b_inv_c_3, b_inv_c_2, 
        b_inv_c_1, b_inv_c_0, c_inv_c_15, c_inv_c_14, c_inv_c_13, 
        c_inv_c_12, c_inv_c_11, c_inv_c_10, c_inv_c_9, c_inv_c_8, 
        c_inv_c_7, c_inv_c_6, c_inv_c_5, c_inv_c_4, c_inv_c_3, c_inv_c_2, 
        c_inv_c_1, c_inv_c_0, d_inv_c_15, d_inv_c_14, d_inv_c_13, 
        d_inv_c_12, d_inv_c_11, d_inv_c_10, d_inv_c_9, d_inv_c_8, 
        d_inv_c_7, d_inv_c_6, d_inv_c_5, d_inv_c_4, d_inv_c_3, d_inv_c_2, 
        d_inv_c_1, d_inv_c_0, error_c;
    wire [31:0]det_q4_28;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(31[34:43])
    
    wire n10519, n10560, n10520, n10559, n10521, n10558, n10522, 
        n10557, n10523, n10556, n10524, n10555, n10525, n10554, 
        n10526, n10553;
    wire [15:0]b_reg;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(32[41:46])
    wire [15:0]c_reg;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(32[48:53])
    
    wire n10527, n10552, n10528, n10551, n10529, n10550, n10530, 
        n10549, n10531, n10548, n10532, n10547, n10533, n10546, 
        n10534, n10545, det_zero, n10313, n10011, n10314, n10010, 
        n10315, n9817, n9816, n9815, n9814, n9813, n9812, n9811, 
        n9810, n9809, n9808, n9807, n9806, n9805, n9804, n9803, 
        n9802, n10027, n10026, n10025, n10024, n10023, n10022, 
        n10021, n10020, n10019, n10018, n10017, error_recip, n10535, 
        n10213;
    wire [31:0]b_s;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[24:27])
    wire [31:0]c_s;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[24:27])
    wire [47:0]prod_a;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[35:41])
    
    wire n10544, n10536, n10216, n10543, n10537, n10542, n10226, 
        n10772, n10009, n10773, n10008, n10774, n10007, n10775, 
        n10006, n10776, n10005, n10777, n10004, n10778, n10003, 
        n10779, n9801, n9800, n9799, n9798;
    wire [47:0]prod_b;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[35:41])
    
    wire n9797, n10214, n10538, n9796, n9795, n9794, n9793, n9792, 
        n9791, n9790, n9789, n9788, n9787, n9786, n10541, n10539, 
        n10540, n10108, n10109, n10110, n10111, n10112, n10113, 
        n10114, n10115, n10116, n10117, n10118, n10119, n10120, 
        n10121, n10122;
    wire [47:0]prod_c;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[35:41])
    
    wire n10123, n10228, n10124, n10125, n10126, n10127, n10128, 
        n10129, n64, n63, n10215, n62, n61, n60, n59, n58, 
        n57, n56, n55, n54, n53, n52, n51, n50, n49, n48, 
        n47, n46;
    wire [47:0]prod_d;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[35:41])
    
    wire n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, 
        n35, n34, n33, n10237;
    wire [31:0]det_q4_28_31__N_33;
    wire [31:0]det_q4_28_31__N_65;
    wire [31:0]det_q4_28_31__N_1;
    
    wire n1036, n1037, n1033, n1039, n1038, n1035, n1034, n1040, 
        n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
        n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
        n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
        n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
        n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
        n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
        n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
        n10075, n10074, n10073, n10072, n10071, n10070, n10069, 
        n10068, n10067, n10066, n10065, n10064, n10063, n10062, 
        n10061, n10060, n9785, n9784, n9783, n9782, n9781, n9780, 
        n9779, n9778, n9777, n9776, n9775, n9774, n9773, n9772, 
        n9771, n9770, n9769, n9768, n9767, n9766, n9765, n9764, 
        n9763, n9762, n9761, n9760, n9759, n9758, n9757, n9756, 
        n9755, n9754, n130, n10715, n128, n10714, n126, n10713, 
        n124, n10712, n122, n10711, n120, n10710, n118, n10709, 
        n116, n10708, n114, n10707, n112, n10706, n110, n10705, 
        n108, n10704, n106, n10703, n104, n10702, n102, n10701, 
        n10668, n10700, n10669, n10699, n10670, n10698, n10671, 
        n10697, n10672, n10696, n10673, n10695, n10674, n10694, 
        n10675, n10693, n10676, n10692, n10677, n10691, n10678, 
        n10690, n10679, n10689, n10680, n10688, n10681, n10687, 
        n10682, n10686, n10683, n10685, n68, n10684, n10076, n10667, 
        n10077, n10666, n10078, n10665, n10079, n10664, n10080, 
        n10663, n10081, n10662, n10082, n10661, n10083, n10660, 
        n10084, n10659, n10085, n10658, n10086, n10657, n10087, 
        n10656, n10088, n10655, n10089, n10654, n10090, n10653, 
        n10091, n10652, n10092, n10651, n10093, n10650, n10094, 
        n10649, n10095, n10648, n10096, n10647, n10097, n10646, 
        n10098, n10645, n10099, n10644, n10100, n10643, n10101, 
        n10642, n10102, n10641, n10103, n10640, n10104, n10639, 
        n10105, n10638, n10106, n10637, n10107, n10636, n10572, 
        n10573, n128_adj_164, n10574, n10575, n10576, n125, n10577, 
        n10578, n10579, n122_adj_165, n10580, n10581, n10582, n119, 
        n10583, n10584, n10585, n116_adj_166, n10586, n10587, n10588, 
        n10589, n10590, n10591, n10592, n10593, n10594, n10595, 
        n10596, n10597, n1503, n1504, n1505, n1506, n1507, n1508, 
        n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
        n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
        n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
        n1533, n1534, n1536, n10598, n10599, n10600, n10601, n10602, 
        n10603, n10604, n113, n10605, n10606, n10607, n110_adj_167, 
        n10608, n10609, n10610, n107, n10611, n10612, n10613, 
        n104_adj_168, n10614, n10615, n10616, n101, n10617, n10618, 
        n10619, n9970, n10620, n9969, n10621, n9968, n10622, n9967, 
        n10623, n9966, n10624, n9965, n10625, n9964, n10626, n9963, 
        n10627, n9962, n10628, n9961, n10629, n9960, n10630, n9959, 
        n10631, n9958, n10632, n9957, n10633, n9956, n10634, n9955, 
        n10635, n9753, n9752, n9751, n9750, n9749, n9748, n9747, 
        n9746, n9745, n9744, n9743, n9742, n9741, n9740, n9739, 
        n9738, n10059, n10058, n10057, n10056, n10055, n10054, 
        n10053, n10052, n10051, n10050, n10049, n10048, n10047, 
        n10046, n10045, n10044, n9737, n9736, n9735, n9734, n9733, 
        n9732, n9731, n9730, n9729, n9728, n9727, n9726, n9725, 
        n9724, n9723, n9722, n9721, n9720, n9719, n9718, n9717, 
        n9716, n9715, n9714, n9713, n9712, n9711, n9710, n9709, 
        n9708, n9707, n9706, n10508, n10571, n10509, n10570, n10510, 
        n10569, n10511, n10568, n10512, n10567, n10513, n10566, 
        n10514, n10565, n10515, n10564, n10516, n10563, n10517, 
        n10562, n10518, n10561, n10130, n10131, n10132, n10133, 
        n10134, n10135, n10136, n10137, n10138, n10139, n9954, 
        n10412, n9953, n10413, n9952, n10414, n9951, n10415, n9950, 
        n10416, n9949, n10417, n9948, n10418, n9947, n10419, n9946, 
        n10420, n9945, n10421, n9944, n10422, n9943, n10423, n9942, 
        n10424, n9941, n10425, n9940, n10426, n9939, n10427, n10428, 
        n10429, n10430, n10431, n10432, n10433, n10434, n10435, 
        n10436, n10437, n10438, n10439, n10440, n10441, n10442, 
        n10443, n9938, n10444, n9937, n10445, n9936, n10227, n10446, 
        n9935, n10507, n10506, n10505, n10504, n10503, n10502, 
        n10501, n10500, n10499, n10498, n10497, n10496, n10495, 
        n10494, n10493, n10492, n10491, n10490, n10489, n10488, 
        n10487, n10486, n10485, n10484, n10483, n10482, n10481, 
        n10480, n10479, n2039, n2040, n2041, n2042, n2043, n2044, 
        n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
        n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
        n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
        n2069, n2070, n2072, n10478, n10477, n10476, n10447, n9934, 
        n10448, n9933, n10449, n9932, n10450, n9931, n10451, n9930, 
        n10452, n9929, n10453, n9928, n10454, n9927, n10455, n9926, 
        n10456, n9925, n10457, n9924, n10458, n9923, n10459, n9922, 
        n10460, n9921, n10461, n2139, n9920, n10462, n9919, n10316, 
        n10317, n10318, n10319, n10320, n10321, n10322, n10323, 
        n10324, n10325, n10326, n10327, n10328, n10329, n10330, 
        n10331, n10332, n10333, n10334, n10335, n10336, n10337, 
        n10338, n10339, n10340, n10341, n10342, n10343, n10344, 
        n10345, n10346, n10347, n10463, n9918, n10464, n9917, 
        n10465, n9916, n10466, n9915, n10467, n9914, n10468, n9913, 
        n10469, n9912, n10470, n9911, n10471, n9910, n10472, n9909, 
        n10473, n9908, n10474, n9907, n10475, n9705, n9704, n9703, 
        n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
        n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
        n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, 
        n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, 
        n2273, n9702, n9701, n9700, n9699, n9698, n9697, n9696, 
        n9695, n9694, n9693, n9692, n9691, n9690, n9689, n9688, 
        n9687, n9686, n9685, n9684, n9683, n9682, n9681, n9680, 
        n9679, n9678, n9677, n9676, n9675, n9674, n9673, n9672, 
        n9671, n9670, n9669, n9668, n9667, n9666, n9665, n9664, 
        n9663, n9662, n9661, n9660, n9659, n9658, n10043, n10042, 
        n10041, n10040, n10039, n10038, n10037, n10036, n10035, 
        n10034, n10033, n10032, n10031, n10030, n10029, n10028, 
        n9657, n9656, n9655, n9654, n9653, n9652, n9651, n9650, 
        n9649, n9648, n9647, n9646, n9645, n9644, n9643, n9642, 
        n9641, n9640, n9639, n9638, n9637, n9636, n9635, n9634, 
        n9633, n9632, n9631, n9630, n9629, n9628, n9627, n9626, 
        n98, n10411, n10410, n10409, n95, n10408, n10407, n10406, 
        n92, n10405, n10404, n10403, n89, n10402, n10401, n10400, 
        n86, n10399, n10398, n10397, n83, n10396, n10395, n10394, 
        n80, n10393, n10392, n10391, n77, n10390, n10389, n10388, 
        n74, n10016, n10015, n10014, n10013, n10012, n71, n68_adj_169, 
        n10225, n10387, n10386, n10385, n10384, n10383, n10382, 
        n10381, n10380, n10140, n10141, n10142, n10143, n10144, 
        n10145, n10146, n10147, n10148, n10149, n10150, n10151, 
        n10152, n10153, n10154, n10155, n10156, n10157, n10158, 
        n10159, n10160, n10161, n10162, n10163, n10164, n10165, 
        n10166, n10167, n10168, n10169, n10170, n10171, n9906, 
        n10252, n9905, n10253, n9904, n10254, n9903, n10255, n9902, 
        n10256, n9901, n10257, n9900, n10258, n9899, n10259, n10238, 
        n9898, n102_adj_170, n10260, n130_adj_171, n10251, n3044, 
        n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
        n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, 
        n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
        n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3077, 
        n128_adj_172, n10250, n126_adj_173, n10249, n124_adj_174, 
        n10248, n122_adj_175, n10247, n120_adj_176, n10246, n118_adj_177, 
        n10245, n116_adj_178, n10244, n114_adj_179, n10243, n112_adj_180, 
        n10242, n110_adj_181, n10241, n108_adj_182, n10240, n106_adj_183, 
        n10239, n104_adj_184, n3111, n3112, n3113, n3114, n3115, 
        n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
        n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
        n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
        n3140, n3141, n3142, n13004, n9897, n10231, n10261, n10210, 
        n9896, n10230, n10262, n10211, n9895, n10229, n10263, 
        n10212, n10209, n9894, n10236, n10264, n10205, n9893, 
        n10206, n10265, n10234, n9892, n10207, n10266, n10233, 
        n9891, n10208, n10267, n10232, n10268, n10204, n10269, 
        n9890, n10235, n10270, n10271, n10224, n10272, n10217, 
        n10273, n10223, n10274, n10218, n10275, n10222, n10276, 
        n10219, n10277, n10221, n10278, n68_adj_185, n10279, n10220, 
        n10280, n10203, n10281, n10202, n10282, n10201, n10283, 
        n10200, n9889, n10199, n10284, n10198, n9888, n10197, 
        n10285, n10196, n9887, n10195, n10286, n10194, n9886, 
        n10193, n10287, n10192, n9885, n10191, n10288, n10190, 
        n9884, n10189, n10289, n10188, n9883, n10187, n10290, 
        n10186, n9882, n10185, n10291, n10184, n9881, n10183, 
        n10292, n10182, n9880, n10181, n10293, n10180, n9879, 
        n10179, n10294, n10178, n9878, n10177, n10295, n10176, 
        n9877, n10175, n10296, n10174, n9876, n10173, n10297, 
        n10172, n9875, n10298, n9874, n10299, n9873, n10300, n9872, 
        n10301, n9871, n10302, n9870, n10303, n9869, n10304, n9868, 
        n10305, n9867, n10306, n9866, n10307, n9865, n10308, n9864, 
        n10309, n9863, n10310, n9862, n10311, n9861, n10312, n9860, 
        n9859, n10771, n9858, n10770, n9857, n10769, n9856, n10768, 
        n9855, n10767, n9854, n10766, n9853, n10765, n9852, n10764, 
        n9851, n10763, n9850, n10762, n9849, n10761, n9848, n10760, 
        n9847, n10759, n9846, n10758, n9845, n10757, n9844, n9843, 
        n9842, n9841, n9840, n9839, n9838, n9837, n9836, n9835, 
        n9834, n9833, n9832, n9831, n9830, n9829, n9828, n10724, 
        n9827, n10723, n9826, n10722, n9825, n10721, n9824, n10720, 
        n9823, n10719, n9822, n10718, n9821, n10717, n9820, n10716, 
        n9819, n9818, n10780, n10781, n10782, n10783, n10784, 
        n10785, n10786, n10787, n10788, n10789, n10790, n10791, 
        n10792, n10793, n10794, n10795, n10796, n10797, n10798, 
        n10799, n10800, n10801, n10802, n10803, n10804, n10805, 
        n10806, n10807, n10808, n10809, n10810, n10811, n10812, 
        n10813, n10814, n10815, n10816, n10817, n10818, n10819, 
        n10820, n10821, n10822, n10823, n10824, n10825, n10826, 
        n10827, n10828, n10829, n10830, n10831, n10832, n10833, 
        n10834, n10835, n10836, n10837, n10838, n10839, n10840, 
        n10841, n10842, n10843, n10844, n10845, n10846, n10847, 
        n10848, n10849, n10850, n10851, n10852, n10853, n10854, 
        n10855, n10856, n10857, n10858, n10859, n10860, n10861, 
        n10862, n10863, n10864, n10865, n10866, n10867, n10868, 
        n10869, n10870, n10871, n10872, n10873, n10874, n10875, 
        n10876, n10877, n10878, n10879, n10880, n10881, n10882, 
        n10883, n10884, n10885, n10886, n10887, n10888, n10889, 
        n10890, n10891, n10892, n10893, n10894, n10895, n10896, 
        n10897, n10898, n10899, n10900, n10901, n10902, n10903, 
        n10904, n10905, n10906, n10907, n10908, n10909, n10910, 
        n10911, n10912, n10913, n10914, n10915, n10916, n10917, 
        n10918, n10919, n10920, n10921, n10922, n10923, n10924, 
        n10925, n10926, n10927, n10928, n10929, n10930, n10931, 
        n10932, n10933, n10934, n10935, n10936, n10937, n10938, 
        n10939, n10940, n10941, n10942, n10943, n10944, n10945, 
        n10946, n10947, n10948, n10949, n10950, n10951, n10952, 
        n10953, n10954, n10955, n10956, n10957, n10958, n10959, 
        n10960, n10961, n10962, n10963, n10964, n10965, n10966, 
        n10967, n10968, n10969, n10970, n10971, n10972, n10973, 
        n10974, n10975, n10976, n10977, n10978, n10979, n10980, 
        n10981, n10982, n10983, n10984, n10985, n10986, n10987, 
        n10988, n10989, n10990, n10991, n10992, n10993, n10994, 
        n10995, n10996, n10997, n10998, n10999, n11000, n11001, 
        n11002, n11003, n11004, n11005, n11006, n11007, n11008, 
        n11009, n11010, n11011, n11012, n11013, n11014, n11015, 
        n11016, n11017, n11018, n11019, n11020, n11021, n11022, 
        n11023, n11024, n11025, n11026, n11027, n11028, n11029, 
        n11030, n11031, n11032, n11033, n11034, n11035, n11036, 
        n11037, n11038, n11039, n11040, n11041, n11042, n11043, 
        n11044, n11045, n11046, n11047, n11048, n11049, n11050, 
        n11051, n11052, n11053, n11054, n11055, n11056, n11057, 
        n11058, n11059, n11060, n11061, n11062, n11063, n11064, 
        n11065, n11066, n11067, n11068, n11069, n11070, n11071, 
        n11072, n11073, n11074, n11075, n11076, n11077, n11078, 
        n11079, n11080, n11081, n11082, n11083, n11084, n11085, 
        n11086, n11087, n11088, n11089, n11090, n11091, n11092, 
        n11093, n11094, n11095, n11096, n11097, n11098, n11099, 
        n11100, n11101, n131, n134, n137, n140, n143, n146, 
        n149, n152, n155, n158, n161, n68_adj_186, n71_adj_187, 
        n74_adj_188, n77_adj_189, n80_adj_190, n83_adj_191, n86_adj_192, 
        n89_adj_193, n92_adj_194, n95_adj_195, n98_adj_196, n101_adj_197, 
        n104_adj_198, n107_adj_199, n110_adj_200, n113_adj_201, n116_adj_202, 
        n119_adj_203, n122_adj_204, n125_adj_205, n128_adj_206, n131_adj_207, 
        n134_adj_208, n137_adj_209, n140_adj_210, n143_adj_211, n146_adj_212, 
        n149_adj_213, n152_adj_214, n155_adj_215, n158_adj_216, n161_adj_217, 
        n68_adj_218, n71_adj_219, n74_adj_220, n77_adj_221, n80_adj_222, 
        n83_adj_223, n86_adj_224, n89_adj_225, n92_adj_226, n95_adj_227, 
        n98_adj_228, n101_adj_229, n104_adj_230, n107_adj_231, n110_adj_232, 
        n113_adj_233, n116_adj_234, n119_adj_235, n122_adj_236, n125_adj_237, 
        n128_adj_238, n131_adj_239, n134_adj_240, n137_adj_241, n140_adj_242, 
        n143_adj_243, n146_adj_244, n149_adj_245, n152_adj_246, n155_adj_247, 
        n158_adj_248, n161_adj_249, n68_adj_250, n71_adj_251, n74_adj_252, 
        n77_adj_253, n80_adj_254, n83_adj_255, n86_adj_256, n89_adj_257, 
        n92_adj_258, n95_adj_259, n98_adj_260, n101_adj_261, n104_adj_262, 
        n107_adj_263, n110_adj_264, n113_adj_265, n116_adj_266, n119_adj_267, 
        n122_adj_268, n125_adj_269, n128_adj_270, n131_adj_271, n134_adj_272, 
        n137_adj_273, n140_adj_274, n143_adj_275, n146_adj_276, n149_adj_277, 
        n152_adj_278, n155_adj_279, n158_adj_280, n161_adj_281, n68_adj_282, 
        n71_adj_283, n74_adj_284, n77_adj_285, n80_adj_286, n83_adj_287, 
        n86_adj_288, n89_adj_289, n92_adj_290, n95_adj_291, n98_adj_292, 
        n101_adj_293, n104_adj_294, n107_adj_295, n110_adj_296, n113_adj_297, 
        n116_adj_298, n119_adj_299, n122_adj_300, n125_adj_301, n128_adj_302, 
        n131_adj_303, n134_adj_304, n137_adj_305, n140_adj_306, n143_adj_307, 
        n146_adj_308, n149_adj_309, n152_adj_310, n155_adj_311, n158_adj_312, 
        n161_adj_313, n71_adj_314, n74_adj_315, n77_adj_316, n80_adj_317, 
        n83_adj_318, n86_adj_319, n89_adj_320, n92_adj_321, n95_adj_322, 
        n98_adj_323, n101_adj_324, n104_adj_325, n107_adj_326, n110_adj_327, 
        n113_adj_328, n116_adj_329, n119_adj_330, n122_adj_331, n125_adj_332, 
        n128_adj_333, n131_adj_334, n134_adj_335, n137_adj_336, n140_adj_337, 
        n143_adj_338, n146_adj_339, n149_adj_340, n152_adj_341, n155_adj_342, 
        n158_adj_343, n161_adj_344, n68_adj_345, n71_adj_346, n74_adj_347, 
        n77_adj_348, n80_adj_349, n83_adj_350, n86_adj_351, n89_adj_352, 
        n92_adj_353, n95_adj_354, n98_adj_355, n101_adj_356, n104_adj_357, 
        n107_adj_358, n110_adj_359, n113_adj_360, n116_adj_361, n119_adj_362, 
        n122_adj_363, n125_adj_364, n128_adj_365, n131_adj_366, n134_adj_367, 
        n137_adj_368, n140_adj_369, n143_adj_370, n146_adj_371, n149_adj_372, 
        n152_adj_373, n155_adj_374, n158_adj_375, n161_adj_376, n68_adj_377, 
        n71_adj_378, n74_adj_379, n77_adj_380, n80_adj_381, n83_adj_382, 
        n86_adj_383, n89_adj_384, n92_adj_385, n95_adj_386, n98_adj_387, 
        n101_adj_388, n104_adj_389, n107_adj_390, n110_adj_391, n113_adj_392, 
        n116_adj_393, n119_adj_394, n122_adj_395, n125_adj_396, n128_adj_397, 
        n131_adj_398, n134_adj_399, n137_adj_400, n140_adj_401, n143_adj_402, 
        n146_adj_403, n149_adj_404, n152_adj_405, n155_adj_406, n158_adj_407, 
        n161_adj_408, n71_adj_409, n74_adj_410, n77_adj_411, n80_adj_412, 
        n83_adj_413, n86_adj_414, n89_adj_415, n92_adj_416, n95_adj_417, 
        n98_adj_418, n101_adj_419, n104_adj_420, n107_adj_421, n110_adj_422, 
        n113_adj_423, n116_adj_424, n119_adj_425, n122_adj_426, n125_adj_427, 
        n128_adj_428, n131_adj_429, n134_adj_430, n137_adj_431, n140_adj_432, 
        n143_adj_433, n146_adj_434, n149_adj_435, n152_adj_436, n155_adj_437, 
        n158_adj_438, n161_adj_439, n68_adj_440, n71_adj_441, n74_adj_442, 
        n77_adj_443, n80_adj_444, n83_adj_445, n86_adj_446, n89_adj_447, 
        n92_adj_448, n95_adj_449, n98_adj_450, n101_adj_451, n104_adj_452, 
        n107_adj_453, n110_adj_454, n113_adj_455, n116_adj_456, n119_adj_457, 
        n122_adj_458, n125_adj_459, n128_adj_460, n131_adj_461, n134_adj_462, 
        n137_adj_463, n140_adj_464, n143_adj_465, n146_adj_466, n149_adj_467, 
        n152_adj_468, n155_adj_469, n158_adj_470, n161_adj_471, n68_adj_472, 
        n71_adj_473, n74_adj_474, n77_adj_475, n80_adj_476, n83_adj_477, 
        n86_adj_478, n89_adj_479, n92_adj_480, n95_adj_481, n98_adj_482, 
        n101_adj_483, n104_adj_484, n107_adj_485, n110_adj_486, n113_adj_487, 
        n116_adj_488, n119_adj_489, n122_adj_490, n125_adj_491, n128_adj_492, 
        n131_adj_493, n134_adj_494, n137_adj_495, n140_adj_496, n143_adj_497, 
        n146_adj_498, n149_adj_499, n152_adj_500, n155_adj_501, n158_adj_502, 
        n161_adj_503, n68_adj_504, n71_adj_505, n74_adj_506, n77_adj_507, 
        n80_adj_508, n83_adj_509, n86_adj_510, n89_adj_511, n92_adj_512, 
        n95_adj_513, n98_adj_514, n101_adj_515, n104_adj_516, n107_adj_517, 
        n110_adj_518, n113_adj_519, n116_adj_520, n119_adj_521, n122_adj_522, 
        n125_adj_523, n128_adj_524, n131_adj_525, n134_adj_526, n137_adj_527, 
        n140_adj_528, n143_adj_529, n146_adj_530, n149_adj_531, n152_adj_532, 
        n155_adj_533, n158_adj_534, n161_adj_535, n68_adj_536, n71_adj_537, 
        n74_adj_538, n77_adj_539, n80_adj_540, n83_adj_541, n86_adj_542, 
        n89_adj_543, n92_adj_544, n95_adj_545, n98_adj_546, n101_adj_547, 
        n104_adj_548, n107_adj_549, n110_adj_550, n113_adj_551, n116_adj_552, 
        n119_adj_553, n122_adj_554, n125_adj_555, n128_adj_556, n131_adj_557, 
        n134_adj_558, n137_adj_559, n140_adj_560, n143_adj_561, n146_adj_562, 
        n149_adj_563, n152_adj_564, n155_adj_565, n158_adj_566, n161_adj_567, 
        n68_adj_568, n71_adj_569, n74_adj_570, n77_adj_571, n80_adj_572, 
        n83_adj_573, n86_adj_574, n89_adj_575, n92_adj_576, n95_adj_577, 
        n98_adj_578, n101_adj_579, n104_adj_580, n107_adj_581, n110_adj_582, 
        n113_adj_583, n116_adj_584, n119_adj_585, n122_adj_586, n125_adj_587, 
        n128_adj_588, n131_adj_589, n134_adj_590, n137_adj_591, n140_adj_592, 
        n143_adj_593, n146_adj_594, n149_adj_595, n152_adj_596, n155_adj_597, 
        n158_adj_598, n161_adj_599, n68_adj_600, n71_adj_601, n74_adj_602, 
        n77_adj_603, n80_adj_604, n83_adj_605, n86_adj_606, n89_adj_607, 
        n92_adj_608, n95_adj_609, n98_adj_610, n101_adj_611, n104_adj_612, 
        n107_adj_613, n110_adj_614, n113_adj_615, n116_adj_616, n119_adj_617, 
        n122_adj_618, n125_adj_619, n128_adj_620, n131_adj_621, n134_adj_622, 
        n137_adj_623, n140_adj_624, n143_adj_625, n146_adj_626, n149_adj_627, 
        n152_adj_628, n155_adj_629, n158_adj_630, n161_adj_631, n68_adj_632, 
        n71_adj_633, n74_adj_634, n77_adj_635, n80_adj_636, n83_adj_637, 
        n86_adj_638, n89_adj_639, n92_adj_640, n95_adj_641, n98_adj_642, 
        n101_adj_643, n104_adj_644, n107_adj_645, n110_adj_646, n113_adj_647, 
        n116_adj_648, n119_adj_649, n122_adj_650, n125_adj_651, n128_adj_652, 
        n131_adj_653, n134_adj_654, n137_adj_655, n140_adj_656, n143_adj_657, 
        n146_adj_658, n149_adj_659, n152_adj_660, n155_adj_661, n158_adj_662, 
        n161_adj_663, n68_adj_664, n71_adj_665, n74_adj_666, n77_adj_667, 
        n80_adj_668, n83_adj_669, n86_adj_670, n89_adj_671, n92_adj_672, 
        n95_adj_673, n98_adj_674, n101_adj_675, n104_adj_676, n107_adj_677, 
        n110_adj_678, n113_adj_679, n116_adj_680, n119_adj_681, n122_adj_682, 
        n125_adj_683, n128_adj_684, n131_adj_685, n134_adj_686, n137_adj_687, 
        n140_adj_688, n143_adj_689, n146_adj_690, n149_adj_691, n152_adj_692, 
        n155_adj_693, n158_adj_694, n161_adj_695, n68_adj_696, n71_adj_697, 
        n74_adj_698, n77_adj_699, n80_adj_700, n83_adj_701, n86_adj_702, 
        n89_adj_703, n92_adj_704, n95_adj_705, n98_adj_706, n101_adj_707, 
        n104_adj_708, n107_adj_709, n110_adj_710, n113_adj_711, n116_adj_712, 
        n119_adj_713, n122_adj_714, n125_adj_715, n128_adj_716, n131_adj_717, 
        n134_adj_718, n137_adj_719, n140_adj_720, n143_adj_721, n146_adj_722, 
        n149_adj_723, n152_adj_724, n155_adj_725, n158_adj_726, n161_adj_727, 
        n68_adj_728, n71_adj_729, n74_adj_730, n77_adj_731, n80_adj_732, 
        n83_adj_733, n86_adj_734, n89_adj_735, n92_adj_736, n95_adj_737, 
        n98_adj_738, n101_adj_739, n104_adj_740, n107_adj_741, n110_adj_742, 
        n113_adj_743, n116_adj_744, n119_adj_745, n122_adj_746, n125_adj_747, 
        n128_adj_748, n131_adj_749, n134_adj_750, n137_adj_751, n140_adj_752, 
        n143_adj_753, n146_adj_754, n149_adj_755, n152_adj_756, n155_adj_757, 
        n158_adj_758, n161_adj_759, n68_adj_760, n71_adj_761, n74_adj_762, 
        n77_adj_763, n80_adj_764, n83_adj_765, n86_adj_766, n89_adj_767, 
        n92_adj_768, n95_adj_769, n98_adj_770, n101_adj_771, n104_adj_772, 
        n107_adj_773, n110_adj_774, n113_adj_775, n116_adj_776, n119_adj_777, 
        n122_adj_778, n125_adj_779, n128_adj_780, n131_adj_781, n134_adj_782, 
        n137_adj_783, n140_adj_784, n143_adj_785, n146_adj_786, n149_adj_787, 
        n152_adj_788, n155_adj_789, n158_adj_790, n161_adj_791, n68_adj_792, 
        n71_adj_793, n74_adj_794, n77_adj_795, n80_adj_796, n83_adj_797, 
        n86_adj_798, n89_adj_799, n92_adj_800, n95_adj_801, n98_adj_802, 
        n101_adj_803, n104_adj_804, n107_adj_805, n110_adj_806, n113_adj_807, 
        n116_adj_808, n119_adj_809, n122_adj_810, n125_adj_811, n128_adj_812, 
        n131_adj_813, n134_adj_814, n137_adj_815, n140_adj_816, n143_adj_817, 
        n146_adj_818, n149_adj_819, n152_adj_820, n155_adj_821, n158_adj_822, 
        n71_adj_823, n74_adj_824, n77_adj_825, n80_adj_826, n83_adj_827, 
        n86_adj_828, n89_adj_829, n92_adj_830, n95_adj_831, n98_adj_832, 
        n101_adj_833, n104_adj_834, n107_adj_835, n110_adj_836, n113_adj_837, 
        n116_adj_838, n119_adj_839, n122_adj_840, n125_adj_841, n128_adj_842, 
        n131_adj_843, n134_adj_844, n137_adj_845, n140_adj_846, n143_adj_847, 
        n146_adj_848, n149_adj_849, n152_adj_850, n155_adj_851, n158_adj_852, 
        n161_adj_853, n68_adj_854, n71_adj_855, n74_adj_856, n77_adj_857, 
        n80_adj_858, n83_adj_859, n86_adj_860, n89_adj_861, n92_adj_862, 
        n95_adj_863, n98_adj_864, n101_adj_865, n104_adj_866, n107_adj_867, 
        n110_adj_868, n113_adj_869, n116_adj_870, n119_adj_871, n122_adj_872, 
        n125_adj_873, n128_adj_874, n131_adj_875, n134_adj_876, n137_adj_877, 
        n140_adj_878, n143_adj_879, n146_adj_880, n149_adj_881, n152_adj_882, 
        n155_adj_883, n158_adj_884, n161_adj_885, n68_adj_886, n71_adj_887, 
        n74_adj_888, n77_adj_889, n80_adj_890, n83_adj_891, n86_adj_892, 
        n89_adj_893, n92_adj_894, n95_adj_895, n98_adj_896, n101_adj_897, 
        n104_adj_898, n107_adj_899, n110_adj_900, n113_adj_901, n116_adj_902, 
        n119_adj_903, n122_adj_904, n125_adj_905, n128_adj_906, n131_adj_907, 
        n134_adj_908, n137_adj_909, n140_adj_910, n143_adj_911, n146_adj_912, 
        n149_adj_913, n152_adj_914, n155_adj_915, n158_adj_916, n161_adj_917, 
        n68_adj_918, n71_adj_919, n74_adj_920, n77_adj_921, n80_adj_922, 
        n83_adj_923, n86_adj_924, n89_adj_925, n92_adj_926, n95_adj_927, 
        n98_adj_928, n101_adj_929, n104_adj_930, n107_adj_931, n110_adj_932, 
        n113_adj_933, n116_adj_934, n119_adj_935, n122_adj_936, n125_adj_937, 
        n128_adj_938, n131_adj_939, n134_adj_940, n137_adj_941, n140_adj_942, 
        n143_adj_943, n146_adj_944, n149_adj_945, n152_adj_946, n155_adj_947, 
        n158_adj_948, n161_adj_949, n68_adj_950, n71_adj_951, n74_adj_952, 
        n77_adj_953, n80_adj_954, n83_adj_955, n86_adj_956, n89_adj_957, 
        n92_adj_958, n95_adj_959, n98_adj_960, n101_adj_961, n104_adj_962, 
        n107_adj_963, n110_adj_964, n113_adj_965, n116_adj_966, n119_adj_967, 
        n122_adj_968, n125_adj_969, n128_adj_970, n131_adj_971, n134_adj_972, 
        n137_adj_973, n140_adj_974, n143_adj_975, n146_adj_976, n149_adj_977, 
        n152_adj_978, n155_adj_979, n158_adj_980, n161_adj_981, n68_adj_982, 
        n71_adj_983, n74_adj_984, n77_adj_985, n80_adj_986, n83_adj_987, 
        n86_adj_988, n89_adj_989, n92_adj_990, n95_adj_991, n98_adj_992, 
        n101_adj_993, n104_adj_994, n107_adj_995, n110_adj_996, n113_adj_997, 
        n116_adj_998, n119_adj_999, n122_adj_1000, n125_adj_1001, n128_adj_1002, 
        n131_adj_1003, n134_adj_1004, n137_adj_1005, n140_adj_1006, 
        n143_adj_1007, n146_adj_1008, n149_adj_1009, n152_adj_1010, 
        n155_adj_1011, n158_adj_1012, n161_adj_1013, n68_adj_1014, n71_adj_1015, 
        n74_adj_1016, n77_adj_1017, n80_adj_1018, n83_adj_1019, n86_adj_1020, 
        n89_adj_1021, n92_adj_1022, n95_adj_1023, n98_adj_1024, n101_adj_1025, 
        n104_adj_1026, n107_adj_1027, n110_adj_1028, n113_adj_1029, 
        n116_adj_1030, n119_adj_1031, n122_adj_1032, n125_adj_1033, 
        n128_adj_1034, n131_adj_1035, n134_adj_1036, n137_adj_1037, 
        n140_adj_1038, n143_adj_1039, n146_adj_1040, n149_adj_1041, 
        n152_adj_1042, n155_adj_1043, n158_adj_1044, n161_adj_1045, 
        n68_adj_1046, n71_adj_1047, n74_adj_1048, n77_adj_1049, n80_adj_1050, 
        n83_adj_1051, n86_adj_1052, n89_adj_1053, n92_adj_1054, n95_adj_1055, 
        n98_adj_1056, n101_adj_1057, n104_adj_1058, n107_adj_1059, n110_adj_1060, 
        n113_adj_1061, n116_adj_1062, n119_adj_1063, n122_adj_1064, 
        n125_adj_1065, n128_adj_1066, n131_adj_1067, n134_adj_1068, 
        n137_adj_1069, n140_adj_1070, n143_adj_1071, n146_adj_1072, 
        n149_adj_1073, n152_adj_1074, n155_adj_1075, n158_adj_1076, 
        n161_adj_1077, n68_adj_1078, n71_adj_1079, n74_adj_1080, n77_adj_1081, 
        n80_adj_1082, n83_adj_1083, n86_adj_1084, n89_adj_1085, n92_adj_1086, 
        n95_adj_1087, n98_adj_1088, n101_adj_1089, n104_adj_1090, n107_adj_1091, 
        n110_adj_1092, n113_adj_1093, n116_adj_1094, n119_adj_1095, 
        n122_adj_1096, n125_adj_1097, n128_adj_1098, n131_adj_1099, 
        n134_adj_1100, n137_adj_1101, n140_adj_1102, n143_adj_1103, 
        n146_adj_1104, n149_adj_1105, n152_adj_1106, n155_adj_1107, 
        n158_adj_1108, n161_adj_1109, n68_adj_1110, n71_adj_1111, n74_adj_1112, 
        n77_adj_1113, n80_adj_1114, n83_adj_1115, n86_adj_1116, n89_adj_1117, 
        n92_adj_1118, n95_adj_1119, n98_adj_1120, n101_adj_1121, n104_adj_1122, 
        n107_adj_1123, n110_adj_1124, n113_adj_1125, n116_adj_1126, 
        n119_adj_1127, n122_adj_1128, n125_adj_1129, n128_adj_1130, 
        n131_adj_1131, n134_adj_1132, n137_adj_1133, n140_adj_1134, 
        n143_adj_1135, n146_adj_1136, n149_adj_1137, n152_adj_1138, 
        n155_adj_1139, n158_adj_1140, n161_adj_1141, n68_adj_1142, n68_adj_1143, 
        n71_adj_1144, n74_adj_1145, n77_adj_1146, n80_adj_1147, n83_adj_1148, 
        n86_adj_1149, n89_adj_1150, n92_adj_1151, n95_adj_1152, n98_adj_1153, 
        n101_adj_1154, n104_adj_1155, n107_adj_1156, n110_adj_1157, 
        n113_adj_1158, n116_adj_1159, n119_adj_1160, n122_adj_1161, 
        n125_adj_1162, n128_adj_1163, n131_adj_1164, n134_adj_1165, 
        n137_adj_1166, n140_adj_1167, n143_adj_1168, n146_adj_1169, 
        n149_adj_1170, n152_adj_1171, n155_adj_1172, n158_adj_1173, 
        n161_adj_1174, n68_adj_1175, n71_adj_1176, n74_adj_1177, n77_adj_1178, 
        n80_adj_1179, n83_adj_1180, n86_adj_1181, n89_adj_1182, n92_adj_1183, 
        n95_adj_1184, n98_adj_1185, n101_adj_1186, n104_adj_1187, n107_adj_1188, 
        n110_adj_1189, n113_adj_1190, n116_adj_1191, n119_adj_1192, 
        n122_adj_1193, n125_adj_1194, n128_adj_1195, n131_adj_1196, 
        n134_adj_1197, n137_adj_1198, n140_adj_1199, n143_adj_1200, 
        n146_adj_1201, n149_adj_1202, n152_adj_1203, n155_adj_1204, 
        n158_adj_1205, n71_adj_1206, n74_adj_1207, n77_adj_1208, n80_adj_1209, 
        n83_adj_1210, n86_adj_1211, n89_adj_1212, n92_adj_1213, n95_adj_1214, 
        n98_adj_1215, n101_adj_1216, n104_adj_1217, n107_adj_1218, n110_adj_1219, 
        n113_adj_1220, n116_adj_1221, n119_adj_1222, n122_adj_1223, 
        n125_adj_1224, n128_adj_1225, n131_adj_1226, n134_adj_1227, 
        n137_adj_1228, n140_adj_1229, n143_adj_1230, n146_adj_1231, 
        n149_adj_1232, n152_adj_1233, n155_adj_1234, n158_adj_1235, 
        n161_adj_1236, n68_adj_1237, n71_adj_1238, n74_adj_1239, n77_adj_1240, 
        n80_adj_1241, n83_adj_1242, n86_adj_1243, n89_adj_1244, n92_adj_1245, 
        n95_adj_1246, n98_adj_1247, n101_adj_1248, n104_adj_1249, n107_adj_1250, 
        n110_adj_1251, n113_adj_1252, n116_adj_1253, n119_adj_1254, 
        n122_adj_1255, n125_adj_1256, n128_adj_1257, n131_adj_1258, 
        n134_adj_1259, n137_adj_1260, n140_adj_1261, n143_adj_1262, 
        n146_adj_1263, n149_adj_1264, n152_adj_1265, n155_adj_1266, 
        n158_adj_1267, n68_adj_1268, n71_adj_1269, n74_adj_1270, n77_adj_1271, 
        n80_adj_1272, n83_adj_1273, n86_adj_1274, n89_adj_1275, n92_adj_1276, 
        n95_adj_1277, n98_adj_1278, n101_adj_1279, n104_adj_1280, n107_adj_1281, 
        n110_adj_1282, n113_adj_1283, n116_adj_1284, n119_adj_1285, 
        n122_adj_1286, n125_adj_1287, n128_adj_1288, n131_adj_1289, 
        n134_adj_1290, n137_adj_1291, n140_adj_1292, n143_adj_1293, 
        n146_adj_1294, n149_adj_1295, n152_adj_1296, n155_adj_1297, 
        n158_adj_1298, n68_adj_1299, n71_adj_1300, n74_adj_1301, n77_adj_1302, 
        n80_adj_1303, n83_adj_1304, n86_adj_1305, n89_adj_1306, n92_adj_1307, 
        n95_adj_1308, n98_adj_1309, n101_adj_1310, n104_adj_1311, n107_adj_1312, 
        n110_adj_1313, n113_adj_1314, n116_adj_1315, n119_adj_1316, 
        n122_adj_1317, n125_adj_1318, n128_adj_1319, n131_adj_1320, 
        n134_adj_1321, n137_adj_1322, n140_adj_1323, n143_adj_1324, 
        n146_adj_1325, n149_adj_1326, n152_adj_1327, n155_adj_1328, 
        n158_adj_1329, n68_adj_1330, n71_adj_1331, n74_adj_1332, n77_adj_1333, 
        n80_adj_1334, n83_adj_1335, n86_adj_1336, n89_adj_1337, n92_adj_1338, 
        n95_adj_1339, n98_adj_1340, n101_adj_1341, n104_adj_1342, n107_adj_1343, 
        n110_adj_1344, n113_adj_1345, n116_adj_1346, n119_adj_1347, 
        n122_adj_1348, n125_adj_1349, n128_adj_1350, n131_adj_1351, 
        n134_adj_1352, n137_adj_1353, n140_adj_1354, n143_adj_1355, 
        n146_adj_1356, n149_adj_1357, n152_adj_1358, n155_adj_1359, 
        n158_adj_1360, n161_adj_1361, n68_adj_1362, n71_adj_1363, n74_adj_1364, 
        n77_adj_1365, n80_adj_1366, n83_adj_1367, n86_adj_1368, n89_adj_1369, 
        n92_adj_1370, n95_adj_1371, n98_adj_1372, n101_adj_1373, n104_adj_1374, 
        n107_adj_1375, n110_adj_1376, n113_adj_1377, n116_adj_1378, 
        n119_adj_1379, n122_adj_1380, n125_adj_1381, n128_adj_1382, 
        n131_adj_1383, n134_adj_1384, n137_adj_1385, n140_adj_1386, 
        n143_adj_1387, n146_adj_1388, n149_adj_1389, n152_adj_1390, 
        n155_adj_1391, n158_adj_1392, n161_adj_1393, n68_adj_1394, n71_adj_1395, 
        n74_adj_1396, n77_adj_1397, n80_adj_1398, n83_adj_1399, n86_adj_1400, 
        n89_adj_1401, n92_adj_1402, n95_adj_1403, n98_adj_1404, n101_adj_1405, 
        n104_adj_1406, n107_adj_1407, n110_adj_1408, n113_adj_1409, 
        n116_adj_1410, n119_adj_1411, n122_adj_1412, n125_adj_1413, 
        n128_adj_1414, n131_adj_1415, n134_adj_1416, n137_adj_1417, 
        n140_adj_1418, n143_adj_1419, n146_adj_1420, n149_adj_1421, 
        n152_adj_1422, n155_adj_1423, n158_adj_1424, n161_adj_1425, 
        n68_adj_1426, n71_adj_1427, n74_adj_1428, n77_adj_1429, n80_adj_1430, 
        n83_adj_1431, n86_adj_1432, n89_adj_1433, n92_adj_1434, n95_adj_1435, 
        n98_adj_1436, n101_adj_1437, n104_adj_1438, n107_adj_1439, n110_adj_1440, 
        n113_adj_1441, n116_adj_1442, n119_adj_1443, n122_adj_1444, 
        n125_adj_1445, n128_adj_1446, n131_adj_1447, n134_adj_1448, 
        n137_adj_1449, n140_adj_1450, n143_adj_1451, n146_adj_1452, 
        n149_adj_1453, n152_adj_1454, n155_adj_1455, n158_adj_1456, 
        n161_adj_1457, n68_adj_1458, n71_adj_1459, n74_adj_1460, n77_adj_1461, 
        n80_adj_1462, n83_adj_1463, n86_adj_1464, n89_adj_1465, n92_adj_1466, 
        n95_adj_1467, n98_adj_1468, n101_adj_1469, n104_adj_1470, n107_adj_1471, 
        n110_adj_1472, n113_adj_1473, n116_adj_1474, n119_adj_1475, 
        n122_adj_1476, n125_adj_1477, n128_adj_1478, n131_adj_1479, 
        n134_adj_1480, n137_adj_1481, n140_adj_1482, n143_adj_1483, 
        n146_adj_1484, n149_adj_1485, n152_adj_1486, n155_adj_1487, 
        n158_adj_1488, n161_adj_1489, n68_adj_1490, n71_adj_1491, n74_adj_1492, 
        n77_adj_1493, n80_adj_1494, n83_adj_1495, n86_adj_1496, n89_adj_1497, 
        n92_adj_1498, n95_adj_1499, n98_adj_1500, n101_adj_1501, n104_adj_1502, 
        n107_adj_1503, n110_adj_1504, n113_adj_1505, n116_adj_1506, 
        n119_adj_1507, n122_adj_1508, n125_adj_1509, n128_adj_1510, 
        n131_adj_1511, n134_adj_1512, n137_adj_1513, n140_adj_1514, 
        n143_adj_1515, n146_adj_1516, n149_adj_1517, n152_adj_1518, 
        n155_adj_1519, n158_adj_1520, n161_adj_1521, n68_adj_1522, n71_adj_1523, 
        n74_adj_1524, n77_adj_1525, n80_adj_1526, n83_adj_1527, n86_adj_1528, 
        n89_adj_1529, n92_adj_1530, n95_adj_1531, n98_adj_1532, n101_adj_1533, 
        n104_adj_1534, n107_adj_1535, n110_adj_1536, n113_adj_1537, 
        n116_adj_1538, n119_adj_1539, n122_adj_1540, n125_adj_1541, 
        n128_adj_1542, n131_adj_1543, n134_adj_1544, n137_adj_1545, 
        n140_adj_1546, n143_adj_1547, n146_adj_1548, n149_adj_1549, 
        n152_adj_1550, n155_adj_1551, n158_adj_1552, n161_adj_1553, 
        n68_adj_1554, n71_adj_1555, n74_adj_1556, n77_adj_1557, n80_adj_1558, 
        n83_adj_1559, n86_adj_1560, n89_adj_1561, n92_adj_1562, n95_adj_1563, 
        n98_adj_1564, n101_adj_1565, n104_adj_1566, n107_adj_1567, n110_adj_1568, 
        n113_adj_1569, n116_adj_1570, n119_adj_1571, n122_adj_1572, 
        n125_adj_1573, n128_adj_1574, n131_adj_1575, n134_adj_1576, 
        n137_adj_1577, n140_adj_1578, n143_adj_1579, n146_adj_1580, 
        n149_adj_1581, n152_adj_1582, n155_adj_1583, n158_adj_1584, 
        n161_adj_1585, n71_adj_1586, n74_adj_1587, n77_adj_1588, n80_adj_1589, 
        n83_adj_1590, n86_adj_1591, n89_adj_1592, n92_adj_1593, n95_adj_1594, 
        n98_adj_1595, n101_adj_1596, n104_adj_1597, n107_adj_1598, n110_adj_1599, 
        n113_adj_1600, n116_adj_1601, n119_adj_1602, n122_adj_1603, 
        n125_adj_1604, n128_adj_1605, n131_adj_1606, n134_adj_1607, 
        n137_adj_1608, n140_adj_1609, n143_adj_1610, n146_adj_1611, 
        n149_adj_1612, n152_adj_1613, n155_adj_1614, n158_adj_1615, 
        n161_adj_1616, n68_adj_1617, n71_adj_1618, n74_adj_1619, n77_adj_1620, 
        n80_adj_1621, n83_adj_1622, n86_adj_1623, n89_adj_1624, n92_adj_1625, 
        n95_adj_1626, n98_adj_1627, n101_adj_1628, n104_adj_1629, n107_adj_1630, 
        n110_adj_1631, n113_adj_1632, n116_adj_1633, n119_adj_1634, 
        n122_adj_1635, n125_adj_1636, n128_adj_1637, n131_adj_1638, 
        n134_adj_1639, n137_adj_1640, n140_adj_1641, n143_adj_1642, 
        n146_adj_1643, n149_adj_1644, n152_adj_1645, n155_adj_1646, 
        n158_adj_1647, n161_adj_1648, n68_adj_1649, n71_adj_1650, n74_adj_1651, 
        n77_adj_1652, n80_adj_1653, n83_adj_1654, n86_adj_1655, n89_adj_1656, 
        n92_adj_1657, n95_adj_1658, n98_adj_1659, n101_adj_1660, n104_adj_1661, 
        n107_adj_1662, n110_adj_1663, n113_adj_1664, n116_adj_1665, 
        n119_adj_1666, n122_adj_1667, n125_adj_1668, n128_adj_1669, 
        n131_adj_1670, n134_adj_1671, n137_adj_1672, n140_adj_1673, 
        n143_adj_1674, n146_adj_1675, n149_adj_1676, n152_adj_1677, 
        n155_adj_1678, n158_adj_1679, n161_adj_1680, n68_adj_1681, n71_adj_1682, 
        n74_adj_1683, n77_adj_1684, n80_adj_1685, n83_adj_1686, n86_adj_1687, 
        n89_adj_1688, n92_adj_1689, n95_adj_1690, n98_adj_1691, n101_adj_1692, 
        n104_adj_1693, n107_adj_1694, n110_adj_1695, n113_adj_1696, 
        n116_adj_1697, n119_adj_1698, n122_adj_1699, n125_adj_1700, 
        n128_adj_1701, n131_adj_1702, n134_adj_1703, n137_adj_1704, 
        n140_adj_1705, n143_adj_1706, n146_adj_1707, n149_adj_1708, 
        n152_adj_1709, n155_adj_1710, n158_adj_1711, n161_adj_1712, 
        n68_adj_1713, n71_adj_1714, n74_adj_1715, n77_adj_1716, n80_adj_1717, 
        n83_adj_1718, n86_adj_1719, n89_adj_1720, n92_adj_1721, n95_adj_1722, 
        n98_adj_1723, n101_adj_1724, n104_adj_1725, n107_adj_1726, n110_adj_1727, 
        n113_adj_1728, n116_adj_1729, n119_adj_1730, n122_adj_1731, 
        n125_adj_1732, n128_adj_1733, n131_adj_1734, n134_adj_1735, 
        n137_adj_1736, n140_adj_1737, n143_adj_1738, n146_adj_1739, 
        n149_adj_1740, n152_adj_1741, n155_adj_1742, n158_adj_1743, 
        n161_adj_1744, n12806, n12805, n12804, n12803, n12802, n12801, 
        n12800, n12799, n12798, n12797, n12796, n12795, n12794, 
        n12793, n12792, n12791, n12790, n12789, n12788, n12787, 
        n12786, n12785, n12784, n12783, n12782, n12781, n12780, 
        n12779, n12778, n12777, n12776, n12775, n12774, n12773, 
        n12772, n12771, n12770, n12769, n12768, n12767, n12766, 
        n12765, n12764, n12763, n12762, n12761, n12760, n12759, 
        n12758, n68_adj_1745, n12757, n71_adj_1746, n12756, n74_adj_1747, 
        n12755, n77_adj_1748, n12754, n80_adj_1749, n12753, n83_adj_1750, 
        n12752, n86_adj_1751, n12751, n89_adj_1752, n12750, n92_adj_1753, 
        n12749, n95_adj_1754, n12748, n98_adj_1755, n12747, n101_adj_1756, 
        n12746, n104_adj_1757, n12745, n107_adj_1758, n12744, n110_adj_1759, 
        n12743, n113_adj_1760, n116_adj_1761, n12741, n119_adj_1762, 
        n12740, n122_adj_1763, n12739, n125_adj_1764, n12738, n128_adj_1765, 
        n12737, n131_adj_1766, n12736, n134_adj_1767, n12735, n137_adj_1768, 
        n12734, n140_adj_1769, n12733, n143_adj_1770, n12732, n146_adj_1771, 
        n12731, n149_adj_1772, n12730, n152_adj_1773, n12729, n155_adj_1774, 
        n12728, n158_adj_1775, n12727, n161_adj_1776, n12726, n12725, 
        n12724, n12723, n12722, n12721, n12720, n12719, n12718, 
        n12717, n12716, n12715, n12714, n12713, n12712, n12711, 
        n12710, n12709, n12708, n12707, n12706, n12705, n12704, 
        n12703, n12702, n12701, n12700, n12699, n12698, n12697, 
        n12696, n12695, n12694, n12693, n12692, n12691, n12690, 
        n12689, n12688, n12687, n12686, n12685, n12684, n12683, 
        n12682, n12681, n12680, n12679, n12678, n12677, n12676, 
        n12675, n12674, n12673, n12672, n12671, n12670, n12669, 
        n12668, n12667, n12666, n12665, n12664, n12663, n12662, 
        n12661, n68_adj_1777, n12660, n12659, n12658, n12657, n12656, 
        n12655, n12654, n12653, n12652, n12651, n12650, n12649, 
        n12648, n12647, n12646, n12645, n12644, n12643, n12642, 
        n12641, n12640, n12639, n12638, n12637, n12636, n12635, 
        n12634, n12633, n12632, n12631, n12630, n12629, n12628, 
        n12627, n12626, n12625, n12624, n12623, n12622, n12621, 
        n12620, n12619, n12618, n12617, n12616, n12615, n12614, 
        n12613, n12612, n12611, n12610, n12609, n12608, n12607, 
        n12606, n12604, n12603, n12602, n12601, n12600, n12599, 
        n12598, n12597, n12596, n12595, n12594, n12593, n12592, 
        n12591, n12590, n12589, n12588, n12587, n12586, n12585, 
        n12584, n12583, n12582, n12581, n12580, n12579, n12578, 
        n12577, n12576, n12575, n12574, n12573, n12572, n12571, 
        n12570, n12569, n12568, n12567, n12566, n12565, n12564, 
        n12563, n12562, n12561, n12560, n12559, n12558, n12557, 
        n12556, n12555, n12554, n12553, n12552, n12551, n12550, 
        n12549, n12548, n12547, n12546, n12545, n12544, n12543, 
        n12542, n12541, n12540, n12539, n12538, n12537, n12536, 
        n12535, n12534, n12533, n12532, n12531, n12530, n12529, 
        n12528, n12527, n12526, n12525, n12524, n12523, n12522, 
        n12521, n12520, n12519, n12518, n12517, n12516, n12515, 
        n12514, n12513, n12512, n12511, n12510, n12508, n12507, 
        n12506, n12505, n12504, n12503, n12502, n68_adj_1778, n12501, 
        n71_adj_1779, n12500, n74_adj_1780, n12499, n77_adj_1781, 
        n12498, n80_adj_1782, n12497, n83_adj_1783, n12496, n86_adj_1784, 
        n12495, n89_adj_1785, n12494, n92_adj_1786, n12493, n95_adj_1787, 
        n98_adj_1788, n101_adj_1789, n12489, n104_adj_1790, n12488, 
        n107_adj_1791, n12487, n110_adj_1792, n12486, n113_adj_1793, 
        n12485, n116_adj_1794, n12484, n119_adj_1795, n12483, n122_adj_1796, 
        n12482, n125_adj_1797, n12481, n128_adj_1798, n12480, n131_adj_1799, 
        n12479, n134_adj_1800, n12478, n137_adj_1801, n12477, n140_adj_1802, 
        n12476, n143_adj_1803, n12475, n146_adj_1804, n12474, n149_adj_1805, 
        n12473, n152_adj_1806, n12472, n155_adj_1807, n12471, n158_adj_1808, 
        n12470, n161_adj_1809, n12469, n12468, n12467, n12466, n12465, 
        n12464, n12463, n12462, n12461, n12460, n12459, n12458, 
        n12457, n12456, n12455, n12454, n12453, n12452, n12451, 
        n12450, n12449, n12448, n12447, n12446, n12445, n12444, 
        n12443, n12442, n12441, n12440, n12439, n12438, n12437, 
        n12436, n12435, n12434, n12433, n12432, n12431, n12430, 
        n12429, n12428, n12427, n12426, n12425, n12424, n12423, 
        n12422, n12421, n12420, n12419, n12418, n12417, n12416, 
        n12415, n12414, n12413, n12412, n12411, n12410, n12409, 
        n12408, n12407, n12406, n12405, n12404, n68_adj_1810, n12403, 
        n71_adj_1811, n12402, n74_adj_1812, n12401, n77_adj_1813, 
        n12400, n80_adj_1814, n12399, n83_adj_1815, n12398, n86_adj_1816, 
        n12397, n89_adj_1817, n12396, n92_adj_1818, n12395, n95_adj_1819, 
        n12394, n98_adj_1820, n12393, n101_adj_1821, n12392, n104_adj_1822, 
        n12391, n107_adj_1823, n12390, n110_adj_1824, n12389, n113_adj_1825, 
        n12388, n116_adj_1826, n12387, n119_adj_1827, n12386, n122_adj_1828, 
        n12385, n125_adj_1829, n12384, n128_adj_1830, n12383, n131_adj_1831, 
        n12382, n134_adj_1832, n12381, n137_adj_1833, n12380, n140_adj_1834, 
        n12379, n143_adj_1835, n12378, n146_adj_1836, n12377, n149_adj_1837, 
        n12376, n152_adj_1838, n12375, n155_adj_1839, n12374, n158_adj_1840, 
        n12373, n161_adj_1841, n12372, n12371, n12370, n12369, n12368, 
        n12367, n12366, n12365, n12364, n12363, n12362, n12361, 
        n12360, n12359, n12358, n12357, n12356, n12355, n12354, 
        n12353, n12352, n12351, n12350, n12349, n12348, n12347, 
        n12346, n12344, n12343, n12342, n12341, n12340, n12339, 
        n12338, n12337, n12336, n12335, n12334, n12333, n12332, 
        n12331, n12330, n12327, n12326, n12325, n12324, n12323, 
        n12322, n12321, n12320, n12319, n12318, n12317, n12316, 
        n12315, n12314, n12313, n12310, n12309, n12308, n12307, 
        n12306, n12305, n68_adj_1842, n12304, n71_adj_1843, n12303, 
        n74_adj_1844, n12302, n77_adj_1845, n12301, n80_adj_1846, 
        n12300, n83_adj_1847, n12299, n86_adj_1848, n12298, n89_adj_1849, 
        n12297, n92_adj_1850, n12296, n95_adj_1851, n98_adj_1852, 
        n12293, n101_adj_1853, n12292, n104_adj_1854, n12291, n107_adj_1855, 
        n12290, n110_adj_1856, n12289, n113_adj_1857, n12288, n116_adj_1858, 
        n12287, n119_adj_1859, n12286, n122_adj_1860, n12285, n125_adj_1861, 
        n12284, n128_adj_1862, n12283, n131_adj_1863, n12282, n134_adj_1864, 
        n12281, n137_adj_1865, n12280, n140_adj_1866, n12279, n143_adj_1867, 
        n12278, n146_adj_1868, n149_adj_1869, n152_adj_1870, n155_adj_1871, 
        n12273, n158_adj_1872, n12272, n161_adj_1873, n12271, n12270, 
        n12269, n12268, n12267, n12266, n12265, n12264, n12263, 
        n12262, n12261, n12260, n12259, n12256, n12255, n12254, 
        n12253, n12252, n12251, n12250, n12249, n12248, n12247, 
        n12246, n12245, n12244, n12243, n12242, n12239, n12238, 
        n12237, n12236, n12235, n12234, n12233, n12232, n12231, 
        n12230, n12229, n12228, n12227, n12226, n12225, n12224, 
        n12223, n12222, n12221, n12220, n12219, n12218, n12217, 
        n12216, n12215, n12214, n12213, n12212, n12211, n12210, 
        n12209, n12208, n12207, n12206, n12205, n68_adj_1874, n12204, 
        n71_adj_1875, n12203, n74_adj_1876, n12202, n77_adj_1877, 
        n12201, n80_adj_1878, n12200, n83_adj_1879, n12199, n86_adj_1880, 
        n12198, n89_adj_1881, n12197, n92_adj_1882, n12196, n95_adj_1883, 
        n12195, n98_adj_1884, n12194, n101_adj_1885, n12193, n104_adj_1886, 
        n107_adj_1887, n12191, n110_adj_1888, n12190, n113_adj_1889, 
        n12189, n116_adj_1890, n12188, n119_adj_1891, n12187, n122_adj_1892, 
        n12186, n125_adj_1893, n12185, n128_adj_1894, n12184, n131_adj_1895, 
        n12183, n134_adj_1896, n12182, n137_adj_1897, n12181, n140_adj_1898, 
        n12180, n143_adj_1899, n12179, n146_adj_1900, n12178, n149_adj_1901, 
        n12177, n152_adj_1902, n12176, n155_adj_1903, n12175, n158_adj_1904, 
        n12174, n161_adj_1905, n12173, n12172, n12171, n12170, n12169, 
        n12168, n12167, n12166, n12165, n12164, n12163, n12162, 
        n12161, n12160, n12159, n12158, n12157, n12156, n12155, 
        n12154, n12153, n12152, n12151, n12150, n12149, n12148, 
        n12147, n12146, n12145, n12144, n12143, n12142, n12141, 
        n12140, n12139, n12138, n12137, n12136, n12135, n12134, 
        n12133, n12132, n12131, n12130, n12129, n12128, n12127, 
        n12126, n12125, n12124, n12123, n12122, n12121, n12120, 
        n12119, n12118, n12117, n12116, n12115, n12114, n12113, 
        n12112, n12111, n12110, n12109, n12108, n68_adj_1906, n12107, 
        n71_adj_1907, n12106, n74_adj_1908, n12105, n77_adj_1909, 
        n12104, n80_adj_1910, n12103, n83_adj_1911, n12102, n86_adj_1912, 
        n12101, n89_adj_1913, n12100, n92_adj_1914, n12099, n95_adj_1915, 
        n12098, n98_adj_1916, n12097, n101_adj_1917, n12096, n104_adj_1918, 
        n12095, n107_adj_1919, n12094, n110_adj_1920, n12093, n113_adj_1921, 
        n12092, n116_adj_1922, n12091, n119_adj_1923, n12090, n122_adj_1924, 
        n12089, n125_adj_1925, n12088, n128_adj_1926, n12087, n131_adj_1927, 
        n12086, n134_adj_1928, n12085, n137_adj_1929, n12084, n140_adj_1930, 
        n12083, n143_adj_1931, n12082, n146_adj_1932, n12081, n149_adj_1933, 
        n12080, n152_adj_1934, n12079, n155_adj_1935, n12078, n158_adj_1936, 
        n12077, n161_adj_1937, n12076, n12075, n12074, n12073, n12072, 
        n12070, n12069, n12068, n12067, n12066, n12065, n12064, 
        n12063, n12062, n12061, n12060, n12059, n12058, n12057, 
        n12056, n12055, n12050, n12049, n12048, n12047, n12046, 
        n12045, n12044, n12043, n12042, n12041, n12040, n12039, 
        n12038, n12037, n12036, n12033, n12032, n12031, n12030, 
        n12029, n12028, n12027, n12026, n12025, n12024, n12023, 
        n12022, n12021, n12020, n12019, n12017, n12016, n12015, 
        n12014, n12013, n12012, n12011, n12010, n12009, n12008, 
        n68_adj_1938, n12007, n71_adj_1939, n12006, n74_adj_1940, 
        n12005, n77_adj_1941, n12004, n80_adj_1942, n12003, n83_adj_1943, 
        n12002, n86_adj_1944, n12001, n89_adj_1945, n12000, n92_adj_1946, 
        n11999, n95_adj_1947, n11998, n98_adj_1948, n11997, n101_adj_1949, 
        n11996, n104_adj_1950, n11995, n107_adj_1951, n11994, n110_adj_1952, 
        n11993, n113_adj_1953, n11992, n116_adj_1954, n11991, n119_adj_1955, 
        n11990, n122_adj_1956, n11989, n125_adj_1957, n11988, n128_adj_1958, 
        n11987, n131_adj_1959, n11986, n134_adj_1960, n11985, n137_adj_1961, 
        n11984, n140_adj_1962, n11983, n143_adj_1963, n11982, n146_adj_1964, 
        n11981, n149_adj_1965, n11980, n152_adj_1966, n11979, n155_adj_1967, 
        n11978, n158_adj_1968, n11977, n161_adj_1969, n11976, n11975, 
        n11974, n11973, n11972, n11971, n11970, n11969, n11968, 
        n11967, n11966, n11965, n11964, n11963, n11962, n11961, 
        n11960, n11959, n11958, n11957, n11956, n11955, n11954, 
        n11953, n11952, n11951, n11950, n11949, n11948, n11947, 
        n11946, n11945, n11944, n11943, n11942, n11941, n11940, 
        n11939, n11938, n11937, n11936, n11935, n11934, n11933, 
        n11932, n11931, n11930, n11929, n11928, n11927, n11926, 
        n11925, n11924, n11923, n11922, n11921, n11920, n11919, 
        n11918, n11917, n11916, n11915, n11914, n11913, n11912, 
        n11911, n68_adj_1970, n11910, n71_adj_1971, n11909, n74_adj_1972, 
        n11908, n77_adj_1973, n11907, n80_adj_1974, n11906, n83_adj_1975, 
        n86_adj_1976, n11904, n89_adj_1977, n11903, n92_adj_1978, 
        n11902, n95_adj_1979, n11901, n98_adj_1980, n11900, n101_adj_1981, 
        n11899, n104_adj_1982, n11898, n107_adj_1983, n11897, n110_adj_1984, 
        n11896, n113_adj_1985, n11895, n116_adj_1986, n11894, n119_adj_1987, 
        n11893, n122_adj_1988, n11892, n125_adj_1989, n11891, n128_adj_1990, 
        n11890, n131_adj_1991, n11889, n134_adj_1992, n137_adj_1993, 
        n140_adj_1994, n11885, n143_adj_1995, n11884, n146_adj_1996, 
        n11883, n149_adj_1997, n11882, n152_adj_1998, n11881, n155_adj_1999, 
        n11880, n158_adj_2000, n11879, n161_adj_2001, n11878, n11877, 
        n11876, n11875, n11874, n11873, n11872, n11871, n11870, 
        n11869, n11868, n11867, n11866, n11865, n11864, n11863, 
        n11862, n11861, n11860, n11859, n11858, n11857, n11856, 
        n11855, n11854, n11853, n11852, n11851, n11850, n11849, 
        n11848, n11847, n11846, n11845, n11844, n11843, n11842, 
        n11841, n11840, n11839, n11838, n11836, n11835, n11834, 
        n11833, n11832, n11831, n11830, n11829, n11828, n11827, 
        n11826, n11825, n11824, n11823, n11822, n11821, n11817, 
        n11816, n11815, n11814, n11813, n11812, n11811, n11810, 
        n11809, n11808, n11807, n11806, n11805, n11804, n11803, 
        n11802, n11801, n11800, n11799, n11798, n11797, n11796, 
        n11795, n11794, n11793, n11792, n11791, n11790, n11789, 
        n11788, n11787, n11786, n11785, n11784, n11783, n11782, 
        n11781, n11780, n11779, n11778, n11777, n11776, n11775, 
        n11774, n11773, n11772, n11771, n11770, n11768, n11767, 
        n11766, n11765, n11764, n11763, n11762, n11761, n11760, 
        n11759, n11758, n11757, n11756, n11755, n11754, n11753, 
        n11749, n11748, n11747, n11746, n11745, n11744, n11743, 
        n11742, n11741, n11740, n11739, n11738, n11737, n11736, 
        n11735, n11734, n11733, n11732, n11731, n11730, n11729, 
        n11728, n11727, n11726, n11725, n11724, n11723, n11722, 
        n11721, n11720, n11719, n11718, n11717, n11716, n11715, 
        n11714, n11713, n11712, n68_adj_2002, n11711, n71_adj_2003, 
        n11710, n74_adj_2004, n11709, n77_adj_2005, n11708, n80_adj_2006, 
        n11707, n83_adj_2007, n11706, n86_adj_2008, n11705, n89_adj_2009, 
        n11704, n92_adj_2010, n11703, n95_adj_2011, n11702, n98_adj_2012, 
        n11701, n101_adj_2013, n11700, n104_adj_2014, n11699, n107_adj_2015, 
        n11698, n110_adj_2016, n11697, n113_adj_2017, n11696, n116_adj_2018, 
        n11695, n119_adj_2019, n11694, n122_adj_2020, n11693, n125_adj_2021, 
        n11692, n128_adj_2022, n11691, n131_adj_2023, n11690, n134_adj_2024, 
        n11689, n137_adj_2025, n11688, n140_adj_2026, n11687, n143_adj_2027, 
        n11686, n146_adj_2028, n149_adj_2029, n152_adj_2030, n155_adj_2031, 
        n158_adj_2032, n161_adj_2033, n68_adj_2034, n71_adj_2035, n74_adj_2036, 
        n77_adj_2037, n80_adj_2038, n83_adj_2039, n86_adj_2040, n89_adj_2041, 
        n92_adj_2042, n95_adj_2043, n98_adj_2044, n101_adj_2045, n104_adj_2046, 
        n107_adj_2047, n110_adj_2048, n113_adj_2049, n116_adj_2050, 
        n119_adj_2051, n122_adj_2052, n125_adj_2053, n128_adj_2054, 
        n131_adj_2055, n134_adj_2056, n137_adj_2057, n140_adj_2058, 
        n143_adj_2059, n146_adj_2060, n149_adj_2061, n152_adj_2062, 
        n155_adj_2063, n158_adj_2064, n161_adj_2065, n68_adj_2066, n71_adj_2067, 
        n74_adj_2068, n77_adj_2069, n80_adj_2070, n83_adj_2071, n86_adj_2072, 
        n89_adj_2073, n92_adj_2074, n95_adj_2075, n98_adj_2076, n101_adj_2077, 
        n104_adj_2078, n107_adj_2079, n110_adj_2080, n113_adj_2081, 
        n116_adj_2082, n119_adj_2083, n122_adj_2084, n125_adj_2085, 
        n128_adj_2086, n131_adj_2087, n134_adj_2088, n137_adj_2089, 
        n140_adj_2090, n143_adj_2091, n146_adj_2092, n149_adj_2093, 
        n152_adj_2094, n155_adj_2095, n158_adj_2096, n161_adj_2097, 
        n68_adj_2098, n71_adj_2099, n74_adj_2100, n77_adj_2101, n80_adj_2102, 
        n83_adj_2103, n86_adj_2104, n89_adj_2105, n92_adj_2106, n95_adj_2107, 
        n98_adj_2108, n101_adj_2109, n104_adj_2110, n107_adj_2111, n110_adj_2112, 
        n113_adj_2113, n116_adj_2114, n119_adj_2115, n122_adj_2116, 
        n125_adj_2117, n13028, n128_adj_2118, n13027, n131_adj_2119, 
        n134_adj_2120, n13026, n137_adj_2121, n140_adj_2122, n13025, 
        n143_adj_2123, n146_adj_2124, n13024, n149_adj_2125, n152_adj_2126, 
        n13023, n155_adj_2127, n13022, n158_adj_2128, n161_adj_2129, 
        n13021, n13020, n13019, n13018, n13017, n13016, n13015, 
        n13014, n13013, n13012, n11172, n13011, n13010, n13009, 
        n13008, n13007, n13006, n13005;
    
    VHI i2 (.Z(VCC_net));
    LUT4 mux_315_i1_3_lut_rep_68 (.A(n68_adj_377), .B(n68_adj_345), .C(n2273), 
         .Z(n13004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_315_i1_3_lut_rep_68.init = 16'hcaca;
    OB d_inv_pad_14 (.I(d_inv_c_14), .O(d_inv[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_15 (.I(d_inv_c_15), .O(d_inv[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB c_inv_pad_0 (.I(c_inv_c_0), .O(c_inv[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_1 (.I(c_inv_c_1), .O(c_inv[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_2 (.I(c_inv_c_2), .O(c_inv[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_3 (.I(c_inv_c_3), .O(c_inv[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_4 (.I(c_inv_c_4), .O(c_inv[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_5 (.I(c_inv_c_5), .O(c_inv[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_6 (.I(c_inv_c_6), .O(c_inv[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    FD1S3AX det_q4_28_res1_i0 (.D(det_q4_28_31__N_1[0]), .CK(clk_c), .Q(det_q4_28[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i0.GSR = "ENABLED";
    OB c_inv_pad_7 (.I(c_inv_c_7), .O(c_inv[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_8 (.I(c_inv_c_8), .O(c_inv[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_9 (.I(c_inv_c_9), .O(c_inv[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_10 (.I(c_inv_c_10), .O(c_inv[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_11 (.I(c_inv_c_11), .O(c_inv[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_12 (.I(c_inv_c_12), .O(c_inv[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_13 (.I(c_inv_c_13), .O(c_inv[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_14 (.I(c_inv_c_14), .O(c_inv[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    OB c_inv_pad_15 (.I(c_inv_c_15), .O(c_inv[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[40:45])
    FD1S3AX d_reg_15__I_0_e2__i1 (.D(d_c_0), .CK(clk_c), .Q(n130_adj_171));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i1.GSR = "ENABLED";
    CCU2C _add_1_612_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13015), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11870), .S1(n161));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_612_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_1.INJECT1_1 = "NO";
    OB b_inv_pad_0 (.I(b_inv_c_0), .O(b_inv[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_1 (.I(b_inv_c_1), .O(b_inv[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_2 (.I(b_inv_c_2), .O(b_inv[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_3 (.I(b_inv_c_3), .O(b_inv[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_4 (.I(b_inv_c_4), .O(b_inv[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    CCU2C _add_1_609_add_4_33 (.A0(n1067), .B0(n3077), .C0(n71_adj_283), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11869), .S0(n68_adj_186));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_609_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_609_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_33.INJECT1_1 = "NO";
    OB b_inv_pad_5 (.I(b_inv_c_5), .O(b_inv[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_6 (.I(b_inv_c_6), .O(b_inv[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_7 (.I(b_inv_c_7), .O(b_inv[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_8 (.I(b_inv_c_8), .O(b_inv[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_9 (.I(b_inv_c_9), .O(b_inv[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    CCU2C _add_1_609_add_4_31 (.A0(n77_adj_285), .B0(n3077), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_284), .B1(n3077), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11868), .COUT(n11869), .S0(n74_adj_188), 
          .S1(n71_adj_187));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_31.INJECT1_1 = "NO";
    OB b_inv_pad_10 (.I(b_inv_c_10), .O(b_inv[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    OB b_inv_pad_11 (.I(b_inv_c_11), .O(b_inv[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    IB a_pad_11 (.I(a[11]), .O(a_c_11));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_8 (.I(a[8]), .O(a_c_8));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    OB b_inv_pad_12 (.I(b_inv_c_12), .O(b_inv[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    IB a_pad_7 (.I(a[7]), .O(a_c_7));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB b_pad_13 (.I(b[13]), .O(b_c_13));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    OB b_inv_pad_13 (.I(b_inv_c_13), .O(b_inv[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    CCU2C _add_1_609_add_4_29 (.A0(n83_adj_287), .B0(n3077), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_286), .B1(n3077), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11867), .COUT(n11868), .S0(n80_adj_190), 
          .S1(n77_adj_189));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_29.INJECT1_1 = "NO";
    OB b_inv_pad_14 (.I(b_inv_c_14), .O(b_inv[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    CCU2C _add_1_609_add_4_27 (.A0(n89_adj_289), .B0(n3077), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_288), .B1(n3077), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11866), .COUT(n11867), .S0(n86_adj_192), 
          .S1(n83_adj_191));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_25 (.A0(n95_adj_291), .B0(n3077), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_290), .B1(n3077), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11865), .COUT(n11866), .S0(n92_adj_194), 
          .S1(n89_adj_193));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_25.INJECT1_1 = "NO";
    OB b_inv_pad_15 (.I(b_inv_c_15), .O(b_inv[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[33:38])
    FD1S3AX det_q4_28_res1_i8 (.D(det_q4_28_31__N_1[8]), .CK(clk_c), .Q(det_q4_28[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i8.GSR = "ENABLED";
    OB a_inv_pad_0 (.I(a_inv_c_0), .O(a_inv[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_1 (.I(a_inv_c_1), .O(a_inv[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_2 (.I(a_inv_c_2), .O(a_inv[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_3 (.I(a_inv_c_3), .O(a_inv[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_4 (.I(a_inv_c_4), .O(a_inv[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_5 (.I(a_inv_c_5), .O(a_inv[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_6 (.I(a_inv_c_6), .O(a_inv[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_7 (.I(a_inv_c_7), .O(a_inv[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_8 (.I(a_inv_c_8), .O(a_inv[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_9 (.I(a_inv_c_9), .O(a_inv[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_10 (.I(a_inv_c_10), .O(a_inv[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_11 (.I(a_inv_c_11), .O(a_inv[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_12 (.I(a_inv_c_12), .O(a_inv[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_13 (.I(a_inv_c_13), .O(a_inv[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    OB a_inv_pad_14 (.I(a_inv_c_14), .O(a_inv[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    FD1S3AX a_reg_15__I_0_e2__i1 (.D(a_c_0), .CK(clk_c), .Q(n130));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i1.GSR = "ENABLED";
    MULT18X18D mult_3 (.A17(d_c_15), .A16(d_c_15), .A15(d_c_15), .A14(d_c_14), 
            .A13(d_c_13), .A12(d_c_12), .A11(d_c_11), .A10(d_c_10), 
            .A9(d_c_9), .A8(d_c_8), .A7(d_c_7), .A6(d_c_6), .A5(d_c_5), 
            .A4(d_c_4), .A3(d_c_3), .A2(d_c_2), .A1(d_c_1), .A0(d_c_0), 
            .B17(a_c_15), .B16(a_c_15), .B15(a_c_15), .B14(a_c_14), 
            .B13(a_c_13), .B12(a_c_12), .B11(a_c_11), .B10(a_c_10), 
            .B9(a_c_9), .B8(a_c_8), .B7(a_c_7), .B6(a_c_6), .B5(a_c_5), 
            .B4(a_c_4), .B3(a_c_3), .B2(a_c_2), .B1(a_c_1), .B0(a_c_0), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P31(det_q4_28_31__N_33[31]), 
            .P30(det_q4_28_31__N_33[30]), .P29(det_q4_28_31__N_33[29]), 
            .P28(det_q4_28_31__N_33[28]), .P27(det_q4_28_31__N_33[27]), 
            .P26(det_q4_28_31__N_33[26]), .P25(det_q4_28_31__N_33[25]), 
            .P24(det_q4_28_31__N_33[24]), .P23(det_q4_28_31__N_33[23]), 
            .P22(det_q4_28_31__N_33[22]), .P21(det_q4_28_31__N_33[21]), 
            .P20(det_q4_28_31__N_33[20]), .P19(det_q4_28_31__N_33[19]), 
            .P18(det_q4_28_31__N_33[18]), .P17(det_q4_28_31__N_33[17]), 
            .P16(det_q4_28_31__N_33[16]), .P15(det_q4_28_31__N_33[15]), 
            .P14(det_q4_28_31__N_33[14]), .P13(det_q4_28_31__N_33[13]), 
            .P12(det_q4_28_31__N_33[12]), .P11(det_q4_28_31__N_33[11]), 
            .P10(det_q4_28_31__N_33[10]), .P9(det_q4_28_31__N_33[9]), .P8(det_q4_28_31__N_33[8]), 
            .P7(det_q4_28_31__N_33[7]), .P6(det_q4_28_31__N_33[6]), .P5(det_q4_28_31__N_33[5]), 
            .P4(det_q4_28_31__N_33[4]), .P3(det_q4_28_31__N_33[3]), .P2(det_q4_28_31__N_33[2]), 
            .P1(det_q4_28_31__N_33[1]), .P0(det_q4_28_31__N_33[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:33])
    defparam mult_3.REG_INPUTA_CLK = "NONE";
    defparam mult_3.REG_INPUTA_CE = "CE0";
    defparam mult_3.REG_INPUTA_RST = "RST0";
    defparam mult_3.REG_INPUTB_CLK = "NONE";
    defparam mult_3.REG_INPUTB_CE = "CE0";
    defparam mult_3.REG_INPUTB_RST = "RST0";
    defparam mult_3.REG_INPUTC_CLK = "NONE";
    defparam mult_3.REG_INPUTC_CE = "CE0";
    defparam mult_3.REG_INPUTC_RST = "RST0";
    defparam mult_3.REG_PIPELINE_CLK = "NONE";
    defparam mult_3.REG_PIPELINE_CE = "CE0";
    defparam mult_3.REG_PIPELINE_RST = "RST0";
    defparam mult_3.REG_OUTPUT_CLK = "NONE";
    defparam mult_3.REG_OUTPUT_CE = "CE0";
    defparam mult_3.REG_OUTPUT_RST = "RST0";
    defparam mult_3.CLK0_DIV = "ENABLED";
    defparam mult_3.CLK1_DIV = "ENABLED";
    defparam mult_3.CLK2_DIV = "ENABLED";
    defparam mult_3.CLK3_DIV = "ENABLED";
    defparam mult_3.HIGHSPEED_CLK = "NONE";
    defparam mult_3.GSR = "DISABLED";
    defparam mult_3.CAS_MATCH_REG = "FALSE";
    defparam mult_3.SOURCEB_MODE = "B_SHIFT";
    defparam mult_3.MULT_BYPASS = "DISABLED";
    defparam mult_3.RESETMODE = "SYNC";
    MULT18X18D mult_4 (.A17(c_c_15), .A16(c_c_15), .A15(c_c_15), .A14(c_c_14), 
            .A13(c_c_13), .A12(c_c_12), .A11(c_c_11), .A10(c_c_10), 
            .A9(c_c_9), .A8(c_c_8), .A7(c_c_7), .A6(c_c_6), .A5(c_c_5), 
            .A4(c_c_4), .A3(c_c_3), .A2(c_c_2), .A1(c_c_1), .A0(c_c_0), 
            .B17(b_c_15), .B16(b_c_15), .B15(b_c_15), .B14(b_c_14), 
            .B13(b_c_13), .B12(b_c_12), .B11(b_c_11), .B10(b_c_10), 
            .B9(b_c_9), .B8(b_c_8), .B7(b_c_7), .B6(b_c_6), .B5(b_c_5), 
            .B4(b_c_4), .B3(b_c_3), .B2(b_c_2), .B1(b_c_1), .B0(b_c_0), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P31(det_q4_28_31__N_65[31]), 
            .P30(det_q4_28_31__N_65[30]), .P29(det_q4_28_31__N_65[29]), 
            .P28(det_q4_28_31__N_65[28]), .P27(det_q4_28_31__N_65[27]), 
            .P26(det_q4_28_31__N_65[26]), .P25(det_q4_28_31__N_65[25]), 
            .P24(det_q4_28_31__N_65[24]), .P23(det_q4_28_31__N_65[23]), 
            .P22(det_q4_28_31__N_65[22]), .P21(det_q4_28_31__N_65[21]), 
            .P20(det_q4_28_31__N_65[20]), .P19(det_q4_28_31__N_65[19]), 
            .P18(det_q4_28_31__N_65[18]), .P17(det_q4_28_31__N_65[17]), 
            .P16(det_q4_28_31__N_65[16]), .P15(det_q4_28_31__N_65[15]), 
            .P14(det_q4_28_31__N_65[14]), .P13(det_q4_28_31__N_65[13]), 
            .P12(det_q4_28_31__N_65[12]), .P11(det_q4_28_31__N_65[11]), 
            .P10(det_q4_28_31__N_65[10]), .P9(det_q4_28_31__N_65[9]), .P8(det_q4_28_31__N_65[8]), 
            .P7(det_q4_28_31__N_65[7]), .P6(det_q4_28_31__N_65[6]), .P5(det_q4_28_31__N_65[5]), 
            .P4(det_q4_28_31__N_65[4]), .P3(det_q4_28_31__N_65[3]), .P2(det_q4_28_31__N_65[2]), 
            .P1(det_q4_28_31__N_65[1]), .P0(det_q4_28_31__N_65[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[36:43])
    defparam mult_4.REG_INPUTA_CLK = "NONE";
    defparam mult_4.REG_INPUTA_CE = "CE0";
    defparam mult_4.REG_INPUTA_RST = "RST0";
    defparam mult_4.REG_INPUTB_CLK = "NONE";
    defparam mult_4.REG_INPUTB_CE = "CE0";
    defparam mult_4.REG_INPUTB_RST = "RST0";
    defparam mult_4.REG_INPUTC_CLK = "NONE";
    defparam mult_4.REG_INPUTC_CE = "CE0";
    defparam mult_4.REG_INPUTC_RST = "RST0";
    defparam mult_4.REG_PIPELINE_CLK = "NONE";
    defparam mult_4.REG_PIPELINE_CE = "CE0";
    defparam mult_4.REG_PIPELINE_RST = "RST0";
    defparam mult_4.REG_OUTPUT_CLK = "NONE";
    defparam mult_4.REG_OUTPUT_CE = "CE0";
    defparam mult_4.REG_OUTPUT_RST = "RST0";
    defparam mult_4.CLK0_DIV = "ENABLED";
    defparam mult_4.CLK1_DIV = "ENABLED";
    defparam mult_4.CLK2_DIV = "ENABLED";
    defparam mult_4.CLK3_DIV = "ENABLED";
    defparam mult_4.HIGHSPEED_CLK = "NONE";
    defparam mult_4.GSR = "DISABLED";
    defparam mult_4.CAS_MATCH_REG = "FALSE";
    defparam mult_4.SOURCEB_MODE = "B_SHIFT";
    defparam mult_4.MULT_BYPASS = "DISABLED";
    defparam mult_4.RESETMODE = "SYNC";
    ALU54B lat_alu_19 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10955), .SIGNEDIB(n11028), .SIGNEDCIN(n11101), .A35(n10954), 
           .A34(n10953), .A33(n10952), .A32(n10951), .A31(n10950), .A30(n10949), 
           .A29(n10948), .A28(n10947), .A27(n10946), .A26(n10945), .A25(n10944), 
           .A24(n10943), .A23(n10942), .A22(n10941), .A21(n10940), .A20(n10939), 
           .A19(n10938), .A18(n10937), .A17(n10936), .A16(n10935), .A15(n10934), 
           .A14(n10933), .A13(n10932), .A12(n10931), .A11(n10930), .A10(n10929), 
           .A9(n10928), .A8(n10927), .A7(n10926), .A6(n10925), .A5(n10924), 
           .A4(n10923), .A3(n10922), .A2(n10921), .A1(n10920), .A0(n10919), 
           .B35(n11027), .B34(n11026), .B33(n11025), .B32(n11024), .B31(n11023), 
           .B30(n11022), .B29(n11021), .B28(n11020), .B27(n11019), .B26(n11018), 
           .B25(n11017), .B24(n11016), .B23(n11015), .B22(n11014), .B21(n11013), 
           .B20(n11012), .B19(n11011), .B18(n11010), .B17(n11009), .B16(n11008), 
           .B15(n11007), .B14(n11006), .B13(n11005), .B12(n11004), .B11(n11003), 
           .B10(n11002), .B9(n11001), .B8(n11000), .B7(n10999), .B6(n10998), 
           .B5(n10997), .B4(n10996), .B3(n10995), .B2(n10994), .B1(n10993), 
           .B0(n10992), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10991), .MA34(n10990), .MA33(n10989), .MA32(n10988), 
           .MA31(n10987), .MA30(n10986), .MA29(n10985), .MA28(n10984), 
           .MA27(n10983), .MA26(n10982), .MA25(n10981), .MA24(n10980), 
           .MA23(n10979), .MA22(n10978), .MA21(n10977), .MA20(n10976), 
           .MA19(n10975), .MA18(n10974), .MA17(n10973), .MA16(n10972), 
           .MA15(n10971), .MA14(n10970), .MA13(n10969), .MA12(n10968), 
           .MA11(n10967), .MA10(n10966), .MA9(n10965), .MA8(n10964), 
           .MA7(n10963), .MA6(n10962), .MA5(n10961), .MA4(n10960), .MA3(n10959), 
           .MA2(n10958), .MA1(n10957), .MA0(n10956), .MB35(n11064), 
           .MB34(n11063), .MB33(n11062), .MB32(n11061), .MB31(n11060), 
           .MB30(n11059), .MB29(n11058), .MB28(n11057), .MB27(n11056), 
           .MB26(n11055), .MB25(n11054), .MB24(n11053), .MB23(n11052), 
           .MB22(n11051), .MB21(n11050), .MB20(n11049), .MB19(n11048), 
           .MB18(n11047), .MB17(n11046), .MB16(n11045), .MB15(n11044), 
           .MB14(n11043), .MB13(n11042), .MB12(n11041), .MB11(n11040), 
           .MB10(n11039), .MB9(n11038), .MB8(n11037), .MB7(n11036), 
           .MB6(n11035), .MB5(n11034), .MB4(n11033), .MB3(n11032), .MB2(n11031), 
           .MB1(n11030), .MB0(n11029), .CIN53(n11100), .CIN52(n11099), 
           .CIN51(n11098), .CIN50(n11097), .CIN49(n11096), .CIN48(n11095), 
           .CIN47(n11094), .CIN46(n11093), .CIN45(n11092), .CIN44(n11091), 
           .CIN43(n11090), .CIN42(n11089), .CIN41(n11088), .CIN40(n11087), 
           .CIN39(n11086), .CIN38(n11085), .CIN37(n11084), .CIN36(n11083), 
           .CIN35(n11082), .CIN34(n11081), .CIN33(n11080), .CIN32(n11079), 
           .CIN31(n11078), .CIN30(n11077), .CIN29(n11076), .CIN28(n11075), 
           .CIN27(n11074), .CIN26(n11073), .CIN25(n11072), .CIN24(n11071), 
           .CIN23(n11070), .CIN22(n11069), .CIN21(n11068), .CIN20(n11067), 
           .CIN19(n11066), .CIN18(n11065), .CIN17(d_inv_c_1), .CIN16(d_inv_c_0), 
           .CIN15(n10757), .CIN14(n10758), .CIN13(n10759), .CIN12(n10760), 
           .CIN11(n10761), .CIN10(n10762), .CIN9(n10763), .CIN8(n10764), 
           .CIN7(n10765), .CIN6(n10766), .CIN5(n10767), .CIN4(n10768), 
           .CIN3(n10769), .CIN2(n10770), .CIN1(n10771), .CIN0(n10772), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R13(prod_d[31]), 
           .R12(prod_d[30]), .R11(prod_d[29]), .R10(d_inv_c_12), .R9(d_inv_c_11), 
           .R8(d_inv_c_10), .R7(d_inv_c_9), .R6(d_inv_c_8), .R5(d_inv_c_7), 
           .R4(d_inv_c_6), .R3(d_inv_c_5), .R2(d_inv_c_4), .R1(d_inv_c_3), 
           .R0(d_inv_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam lat_alu_19.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_19.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_19.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_19.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_19.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_19.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_19.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_19.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_19.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_19.REG_FLAG_CLK = "NONE";
    defparam lat_alu_19.REG_FLAG_CE = "CE0";
    defparam lat_alu_19.REG_FLAG_RST = "RST0";
    defparam lat_alu_19.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_19.MASK01 = "0x00000000000000";
    defparam lat_alu_19.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_19.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_19.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_19.CLK0_DIV = "ENABLED";
    defparam lat_alu_19.CLK1_DIV = "ENABLED";
    defparam lat_alu_19.CLK2_DIV = "ENABLED";
    defparam lat_alu_19.CLK3_DIV = "ENABLED";
    defparam lat_alu_19.MCPAT = "0x00000000000000";
    defparam lat_alu_19.MASKPAT = "0x00000000000000";
    defparam lat_alu_19.RNDPAT = "0x00000000000000";
    defparam lat_alu_19.GSR = "DISABLED";
    defparam lat_alu_19.RESETMODE = "SYNC";
    defparam lat_alu_19.MULT9_MODE = "DISABLED";
    defparam lat_alu_19.LEGACY = "DISABLED";
    ALU54B lat_alu_18 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10809), .SIGNEDIB(n10882), .SIGNEDCIN(GND_net), 
           .A35(n10808), .A34(n10807), .A33(n10806), .A32(n10805), .A31(n10804), 
           .A30(n10803), .A29(n10802), .A28(n10801), .A27(n10800), .A26(n10799), 
           .A25(n10798), .A24(n10797), .A23(n10796), .A22(n10795), .A21(n10794), 
           .A20(n10793), .A19(n10792), .A18(n10791), .A17(n10790), .A16(n10789), 
           .A15(n10788), .A14(n10787), .A13(n10786), .A12(n10785), .A11(n10784), 
           .A10(n10783), .A9(n10782), .A8(n10781), .A7(n10780), .A6(n10779), 
           .A5(n10778), .A4(n10777), .A3(n10776), .A2(n10775), .A1(n10774), 
           .A0(n10773), .B35(n10881), .B34(n10880), .B33(n10879), .B32(n10878), 
           .B31(n10877), .B30(n10876), .B29(n10875), .B28(n10874), .B27(n10873), 
           .B26(n10872), .B25(n10871), .B24(n10870), .B23(n10869), .B22(n10868), 
           .B21(n10867), .B20(n10866), .B19(n10865), .B18(n10864), .B17(n10863), 
           .B16(n10862), .B15(n10861), .B14(n10860), .B13(n10859), .B12(n10858), 
           .B11(n10857), .B10(n10856), .B9(n10855), .B8(n10854), .B7(n10853), 
           .B6(n10852), .B5(n10851), .B4(n10850), .B3(n10849), .B2(n10848), 
           .B1(n10847), .B0(n10846), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10845), .MA34(n10844), .MA33(n10843), .MA32(n10842), 
           .MA31(n10841), .MA30(n10840), .MA29(n10839), .MA28(n10838), 
           .MA27(n10837), .MA26(n10836), .MA25(n10835), .MA24(n10834), 
           .MA23(n10833), .MA22(n10832), .MA21(n10831), .MA20(n10830), 
           .MA19(n10829), .MA18(n10828), .MA17(n10827), .MA16(n10826), 
           .MA15(n10825), .MA14(n10824), .MA13(n10823), .MA12(n10822), 
           .MA11(n10821), .MA10(n10820), .MA9(n10819), .MA8(n10818), 
           .MA7(n10817), .MA6(n10816), .MA5(n10815), .MA4(n10814), .MA3(n10813), 
           .MA2(n10812), .MA1(n10811), .MA0(n10810), .MB35(n10918), 
           .MB34(n10917), .MB33(n10916), .MB32(n10915), .MB31(n10914), 
           .MB30(n10913), .MB29(n10912), .MB28(n10911), .MB27(n10910), 
           .MB26(n10909), .MB25(n10908), .MB24(n10907), .MB23(n10906), 
           .MB22(n10905), .MB21(n10904), .MB20(n10903), .MB19(n10902), 
           .MB18(n10901), .MB17(n10900), .MB16(n10899), .MB15(n10898), 
           .MB14(n10897), .MB13(n10896), .MB12(n10895), .MB11(n10894), 
           .MB10(n10893), .MB9(n10892), .MB8(n10891), .MB7(n10890), 
           .MB6(n10889), .MB5(n10888), .MB4(n10887), .MB3(n10886), .MB2(n10885), 
           .MB1(n10884), .MB0(n10883), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n11100), 
           .R52(n11099), .R51(n11098), .R50(n11097), .R49(n11096), .R48(n11095), 
           .R47(n11094), .R46(n11093), .R45(n11092), .R44(n11091), .R43(n11090), 
           .R42(n11089), .R41(n11088), .R40(n11087), .R39(n11086), .R38(n11085), 
           .R37(n11084), .R36(n11083), .R35(n11082), .R34(n11081), .R33(n11080), 
           .R32(n11079), .R31(n11078), .R30(n11077), .R29(n11076), .R28(n11075), 
           .R27(n11074), .R26(n11073), .R25(n11072), .R24(n11071), .R23(n11070), 
           .R22(n11069), .R21(n11068), .R20(n11067), .R19(n11066), .R18(n11065), 
           .R17(d_inv_c_1), .R16(d_inv_c_0), .R15(n10757), .R14(n10758), 
           .R13(n10759), .R12(n10760), .R11(n10761), .R10(n10762), .R9(n10763), 
           .R8(n10764), .R7(n10765), .R6(n10766), .R5(n10767), .R4(n10768), 
           .R3(n10769), .R2(n10770), .R1(n10771), .R0(n10772), .SIGNEDR(n11101));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam lat_alu_18.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_18.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_18.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_18.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_18.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_18.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_18.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_18.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_18.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_18.REG_FLAG_CLK = "NONE";
    defparam lat_alu_18.REG_FLAG_CE = "CE0";
    defparam lat_alu_18.REG_FLAG_RST = "RST0";
    defparam lat_alu_18.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_18.MASK01 = "0x00000000000000";
    defparam lat_alu_18.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_18.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_18.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_18.CLK0_DIV = "ENABLED";
    defparam lat_alu_18.CLK1_DIV = "ENABLED";
    defparam lat_alu_18.CLK2_DIV = "ENABLED";
    defparam lat_alu_18.CLK3_DIV = "ENABLED";
    defparam lat_alu_18.MCPAT = "0x00000000000000";
    defparam lat_alu_18.MASKPAT = "0x00000000000000";
    defparam lat_alu_18.RNDPAT = "0x00000000000000";
    defparam lat_alu_18.GSR = "DISABLED";
    defparam lat_alu_18.RESETMODE = "SYNC";
    defparam lat_alu_18.MULT9_MODE = "DISABLED";
    defparam lat_alu_18.LEGACY = "DISABLED";
    FD1S3AX c_reg_i15 (.D(c_c_15), .CK(clk_c), .Q(c_reg[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i15.GSR = "ENABLED";
    MULT18X18D lat_mult_17 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68), .B16(n68), .B15(n68), 
            .B14(n68), .B13(n68), .B12(n68), .B11(n68), .B10(n68), 
            .B9(n68), .B8(n68), .B7(n68), .B6(n68), .B5(n68), .B4(n68), 
            .B3(n68), .B2(n68), .B1(n68), .B0(n68), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n11009), .ROA16(n11008), .ROA15(n11007), 
            .ROA14(n11006), .ROA13(n11005), .ROA12(n11004), .ROA11(n11003), 
            .ROA10(n11002), .ROA9(n11001), .ROA8(n11000), .ROA7(n10999), 
            .ROA6(n10998), .ROA5(n10997), .ROA4(n10996), .ROA3(n10995), 
            .ROA2(n10994), .ROA1(n10993), .ROA0(n10992), .ROB17(n11027), 
            .ROB16(n11026), .ROB15(n11025), .ROB14(n11024), .ROB13(n11023), 
            .ROB12(n11022), .ROB11(n11021), .ROB10(n11020), .ROB9(n11019), 
            .ROB8(n11018), .ROB7(n11017), .ROB6(n11016), .ROB5(n11015), 
            .ROB4(n11014), .ROB3(n11013), .ROB2(n11012), .ROB1(n11011), 
            .ROB0(n11010), .P35(n11064), .P34(n11063), .P33(n11062), 
            .P32(n11061), .P31(n11060), .P30(n11059), .P29(n11058), 
            .P28(n11057), .P27(n11056), .P26(n11055), .P25(n11054), 
            .P24(n11053), .P23(n11052), .P22(n11051), .P21(n11050), 
            .P20(n11049), .P19(n11048), .P18(n11047), .P17(n11046), 
            .P16(n11045), .P15(n11044), .P14(n11043), .P13(n11042), 
            .P12(n11041), .P11(n11040), .P10(n11039), .P9(n11038), .P8(n11037), 
            .P7(n11036), .P6(n11035), .P5(n11034), .P4(n11033), .P3(n11032), 
            .P2(n11031), .P1(n11030), .P0(n11029), .SIGNEDP(n11028));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam lat_mult_17.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_17.REG_INPUTA_CE = "CE3";
    defparam lat_mult_17.REG_INPUTA_RST = "RST3";
    defparam lat_mult_17.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTB_CE = "CE0";
    defparam lat_mult_17.REG_INPUTB_RST = "RST0";
    defparam lat_mult_17.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_17.REG_INPUTC_CE = "CE0";
    defparam lat_mult_17.REG_INPUTC_RST = "RST0";
    defparam lat_mult_17.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_17.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_17.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_17.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_17.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_17.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_17.CLK0_DIV = "ENABLED";
    defparam lat_mult_17.CLK1_DIV = "ENABLED";
    defparam lat_mult_17.CLK2_DIV = "ENABLED";
    defparam lat_mult_17.CLK3_DIV = "ENABLED";
    defparam lat_mult_17.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_17.GSR = "DISABLED";
    defparam lat_mult_17.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_17.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_17.MULT_BYPASS = "DISABLED";
    defparam lat_mult_17.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_16 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(n68), .B16(n68), .B15(n68), 
            .B14(n68), .B13(n68), .B12(n68), .B11(n68), .B10(n68), 
            .B9(n68), .B8(n68), .B7(n68), .B6(n68), .B5(n68), .B4(n68), 
            .B3(n68), .B2(n68), .B1(n68), .B0(n68), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .ROA17(n10936), .ROA16(n10935), .ROA15(n10934), 
            .ROA14(n10933), .ROA13(n10932), .ROA12(n10931), .ROA11(n10930), 
            .ROA10(n10929), .ROA9(n10928), .ROA8(n10927), .ROA7(n10926), 
            .ROA6(n10925), .ROA5(n10924), .ROA4(n10923), .ROA3(n10922), 
            .ROA2(n10921), .ROA1(n10920), .ROA0(n10919), .ROB17(n10954), 
            .ROB16(n10953), .ROB15(n10952), .ROB14(n10951), .ROB13(n10950), 
            .ROB12(n10949), .ROB11(n10948), .ROB10(n10947), .ROB9(n10946), 
            .ROB8(n10945), .ROB7(n10944), .ROB6(n10943), .ROB5(n10942), 
            .ROB4(n10941), .ROB3(n10940), .ROB2(n10939), .ROB1(n10938), 
            .ROB0(n10937), .P35(n10991), .P34(n10990), .P33(n10989), 
            .P32(n10988), .P31(n10987), .P30(n10986), .P29(n10985), 
            .P28(n10984), .P27(n10983), .P26(n10982), .P25(n10981), 
            .P24(n10980), .P23(n10979), .P22(n10978), .P21(n10977), 
            .P20(n10976), .P19(n10975), .P18(n10974), .P17(n10973), 
            .P16(n10972), .P15(n10971), .P14(n10970), .P13(n10969), 
            .P12(n10968), .P11(n10967), .P10(n10966), .P9(n10965), .P8(n10964), 
            .P7(n10963), .P6(n10962), .P5(n10961), .P4(n10960), .P3(n10959), 
            .P2(n10958), .P1(n10957), .P0(n10956), .SIGNEDP(n10955));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam lat_mult_16.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_16.REG_INPUTA_CE = "CE3";
    defparam lat_mult_16.REG_INPUTA_RST = "RST3";
    defparam lat_mult_16.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTB_CE = "CE0";
    defparam lat_mult_16.REG_INPUTB_RST = "RST0";
    defparam lat_mult_16.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_16.REG_INPUTC_CE = "CE0";
    defparam lat_mult_16.REG_INPUTC_RST = "RST0";
    defparam lat_mult_16.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_16.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_16.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_16.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_16.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_16.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_16.CLK0_DIV = "ENABLED";
    defparam lat_mult_16.CLK1_DIV = "ENABLED";
    defparam lat_mult_16.CLK2_DIV = "ENABLED";
    defparam lat_mult_16.CLK3_DIV = "ENABLED";
    defparam lat_mult_16.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_16.GSR = "DISABLED";
    defparam lat_mult_16.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_16.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_16.MULT_BYPASS = "DISABLED";
    defparam lat_mult_16.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_15 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68), .B16(n68), .B15(n68), 
            .B14(n102), .B13(n104), .B12(n106), .B11(n108), .B10(n110), 
            .B9(n112), .B8(n114), .B7(n116), .B6(n118), .B5(n120), 
            .B4(n122), .B3(n124), .B2(n126), .B1(n128), .B0(n130), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10863), .ROA16(n10862), 
            .ROA15(n10861), .ROA14(n10860), .ROA13(n10859), .ROA12(n10858), 
            .ROA11(n10857), .ROA10(n10856), .ROA9(n10855), .ROA8(n10854), 
            .ROA7(n10853), .ROA6(n10852), .ROA5(n10851), .ROA4(n10850), 
            .ROA3(n10849), .ROA2(n10848), .ROA1(n10847), .ROA0(n10846), 
            .ROB17(n10881), .ROB16(n10880), .ROB15(n10879), .ROB14(n10878), 
            .ROB13(n10877), .ROB12(n10876), .ROB11(n10875), .ROB10(n10874), 
            .ROB9(n10873), .ROB8(n10872), .ROB7(n10871), .ROB6(n10870), 
            .ROB5(n10869), .ROB4(n10868), .ROB3(n10867), .ROB2(n10866), 
            .ROB1(n10865), .ROB0(n10864), .P35(n10918), .P34(n10917), 
            .P33(n10916), .P32(n10915), .P31(n10914), .P30(n10913), 
            .P29(n10912), .P28(n10911), .P27(n10910), .P26(n10909), 
            .P25(n10908), .P24(n10907), .P23(n10906), .P22(n10905), 
            .P21(n10904), .P20(n10903), .P19(n10902), .P18(n10901), 
            .P17(n10900), .P16(n10899), .P15(n10898), .P14(n10897), 
            .P13(n10896), .P12(n10895), .P11(n10894), .P10(n10893), 
            .P9(n10892), .P8(n10891), .P7(n10890), .P6(n10889), .P5(n10888), 
            .P4(n10887), .P3(n10886), .P2(n10885), .P1(n10884), .P0(n10883), 
            .SIGNEDP(n10882));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam lat_mult_15.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_15.REG_INPUTA_CE = "CE3";
    defparam lat_mult_15.REG_INPUTA_RST = "RST3";
    defparam lat_mult_15.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTB_CE = "CE0";
    defparam lat_mult_15.REG_INPUTB_RST = "RST0";
    defparam lat_mult_15.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_15.REG_INPUTC_CE = "CE0";
    defparam lat_mult_15.REG_INPUTC_RST = "RST0";
    defparam lat_mult_15.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_15.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_15.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_15.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_15.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_15.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_15.CLK0_DIV = "ENABLED";
    defparam lat_mult_15.CLK1_DIV = "ENABLED";
    defparam lat_mult_15.CLK2_DIV = "ENABLED";
    defparam lat_mult_15.CLK3_DIV = "ENABLED";
    defparam lat_mult_15.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_15.GSR = "DISABLED";
    defparam lat_mult_15.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_15.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_15.MULT_BYPASS = "DISABLED";
    defparam lat_mult_15.RESETMODE = "ASYNC";
    LUT4 i327_2_lut (.A(prod_d[30]), .B(prod_d[29]), .Z(d_inv_c_14)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i327_2_lut.init = 16'h6666;
    MULT18X18D a_reg_15__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), 
            .A14(n50), .A13(n51), .A12(n52), .A11(n53), .A10(n54), 
            .A9(n55), .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), 
            .A3(n61), .A2(n62), .A1(n63), .A0(n64), .B17(n68), .B16(n68), 
            .B15(n68), .B14(n102), .B13(n104), .B12(n106), .B11(n108), 
            .B10(n110), .B9(n112), .B8(n114), .B7(n116), .B6(n118), 
            .B5(n120), .B4(n122), .B3(n124), .B2(n126), .B1(n128), 
            .B0(n130), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10790), 
            .ROA16(n10789), .ROA15(n10788), .ROA14(n10787), .ROA13(n10786), 
            .ROA12(n10785), .ROA11(n10784), .ROA10(n10783), .ROA9(n10782), 
            .ROA8(n10781), .ROA7(n10780), .ROA6(n10779), .ROA5(n10778), 
            .ROA4(n10777), .ROA3(n10776), .ROA2(n10775), .ROA1(n10774), 
            .ROA0(n10773), .ROB17(n10808), .ROB16(n10807), .ROB15(n10806), 
            .ROB14(n10805), .ROB13(n10804), .ROB12(n10803), .ROB11(n10802), 
            .ROB10(n10801), .ROB9(n10800), .ROB8(n10799), .ROB7(n10798), 
            .ROB6(n10797), .ROB5(n10796), .ROB4(n10795), .ROB3(n10794), 
            .ROB2(n10793), .ROB1(n10792), .ROB0(n10791), .P35(n10845), 
            .P34(n10844), .P33(n10843), .P32(n10842), .P31(n10841), 
            .P30(n10840), .P29(n10839), .P28(n10838), .P27(n10837), 
            .P26(n10836), .P25(n10835), .P24(n10834), .P23(n10833), 
            .P22(n10832), .P21(n10831), .P20(n10830), .P19(n10829), 
            .P18(n10828), .P17(n10827), .P16(n10826), .P15(n10825), 
            .P14(n10824), .P13(n10823), .P12(n10822), .P11(n10821), 
            .P10(n10820), .P9(n10819), .P8(n10818), .P7(n10817), .P6(n10816), 
            .P5(n10815), .P4(n10814), .P3(n10813), .P2(n10812), .P1(n10811), 
            .P0(n10810), .SIGNEDP(n10809));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam a_reg_15__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam a_reg_15__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam a_reg_15__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam a_reg_15__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam a_reg_15__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam a_reg_15__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam a_reg_15__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam a_reg_15__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam a_reg_15__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam a_reg_15__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam a_reg_15__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam a_reg_15__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam a_reg_15__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam a_reg_15__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam a_reg_15__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam a_reg_15__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam a_reg_15__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam a_reg_15__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam a_reg_15__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam a_reg_15__I_0_mult_2.GSR = "DISABLED";
    defparam a_reg_15__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam a_reg_15__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam a_reg_15__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam a_reg_15__I_0_mult_2.RESETMODE = "ASYNC";
    ALU54B lat_alu_14 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10578), .SIGNEDIB(n10651), .SIGNEDCIN(n10724), .A35(n10577), 
           .A34(n10576), .A33(n10575), .A32(n10574), .A31(n10573), .A30(n10572), 
           .A29(n10571), .A28(n10570), .A27(n10569), .A26(n10568), .A25(n10567), 
           .A24(n10566), .A23(n10565), .A22(n10564), .A21(n10563), .A20(n10562), 
           .A19(n10561), .A18(n10560), .A17(n10559), .A16(n10558), .A15(n10557), 
           .A14(n10556), .A13(n10555), .A12(n10554), .A11(n10553), .A10(n10552), 
           .A9(n10551), .A8(n10550), .A7(n10549), .A6(n10548), .A5(n10547), 
           .A4(n10546), .A3(n10545), .A2(n10544), .A1(n10543), .A0(n10542), 
           .B35(n10650), .B34(n10649), .B33(n10648), .B32(n10647), .B31(n10646), 
           .B30(n10645), .B29(n10644), .B28(n10643), .B27(n10642), .B26(n10641), 
           .B25(n10640), .B24(n10639), .B23(n10638), .B22(n10637), .B21(n10636), 
           .B20(n10635), .B19(n10634), .B18(n10633), .B17(n10632), .B16(n10631), 
           .B15(n10630), .B14(n10629), .B13(n10628), .B12(n10627), .B11(n10626), 
           .B10(n10625), .B9(n10624), .B8(n10623), .B7(n10622), .B6(n10621), 
           .B5(n10620), .B4(n10619), .B3(n10618), .B2(n10617), .B1(n10616), 
           .B0(n10615), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10614), .MA34(n10613), .MA33(n10612), .MA32(n10611), 
           .MA31(n10610), .MA30(n10609), .MA29(n10608), .MA28(n10607), 
           .MA27(n10606), .MA26(n10605), .MA25(n10604), .MA24(n10603), 
           .MA23(n10602), .MA22(n10601), .MA21(n10600), .MA20(n10599), 
           .MA19(n10598), .MA18(n10597), .MA17(n10596), .MA16(n10595), 
           .MA15(n10594), .MA14(n10593), .MA13(n10592), .MA12(n10591), 
           .MA11(n10590), .MA10(n10589), .MA9(n10588), .MA8(n10587), 
           .MA7(n10586), .MA6(n10585), .MA5(n10584), .MA4(n10583), .MA3(n10582), 
           .MA2(n10581), .MA1(n10580), .MA0(n10579), .MB35(n10687), 
           .MB34(n10686), .MB33(n10685), .MB32(n10684), .MB31(n10683), 
           .MB30(n10682), .MB29(n10681), .MB28(n10680), .MB27(n10679), 
           .MB26(n10678), .MB25(n10677), .MB24(n10676), .MB23(n10675), 
           .MB22(n10674), .MB21(n10673), .MB20(n10672), .MB19(n10671), 
           .MB18(n10670), .MB17(n10669), .MB16(n10668), .MB15(n10667), 
           .MB14(n10666), .MB13(n10665), .MB12(n10664), .MB11(n10663), 
           .MB10(n10662), .MB9(n10661), .MB8(n10660), .MB7(n10659), 
           .MB6(n10658), .MB5(n10657), .MB4(n10656), .MB3(n10655), .MB2(n10654), 
           .MB1(n10653), .MB0(n10652), .CIN53(n10723), .CIN52(n10722), 
           .CIN51(n10721), .CIN50(n10720), .CIN49(n10719), .CIN48(n10718), 
           .CIN47(n10717), .CIN46(n10716), .CIN45(n10715), .CIN44(n10714), 
           .CIN43(n10713), .CIN42(n10712), .CIN41(n10711), .CIN40(n10710), 
           .CIN39(n10709), .CIN38(n10708), .CIN37(n10707), .CIN36(n10706), 
           .CIN35(n10705), .CIN34(n10704), .CIN33(n10703), .CIN32(n10702), 
           .CIN31(n10701), .CIN30(n10700), .CIN29(n10699), .CIN28(n10698), 
           .CIN27(n10697), .CIN26(n10696), .CIN25(n10695), .CIN24(n10694), 
           .CIN23(n10693), .CIN22(n10692), .CIN21(n10691), .CIN20(n10690), 
           .CIN19(n10689), .CIN18(n10688), .CIN17(c_inv_c_1), .CIN16(c_inv_c_0), 
           .CIN15(n10380), .CIN14(n10381), .CIN13(n10382), .CIN12(n10383), 
           .CIN11(n10384), .CIN10(n10385), .CIN9(n10386), .CIN8(n10387), 
           .CIN7(n10388), .CIN6(n10389), .CIN5(n10390), .CIN4(n10391), 
           .CIN3(n10392), .CIN2(n10393), .CIN1(n10394), .CIN0(n10395), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R13(prod_c[31]), 
           .R12(prod_c[30]), .R11(prod_c[29]), .R10(c_inv_c_12), .R9(c_inv_c_11), 
           .R8(c_inv_c_10), .R7(c_inv_c_9), .R6(c_inv_c_8), .R5(c_inv_c_7), 
           .R4(c_inv_c_6), .R3(c_inv_c_5), .R2(c_inv_c_4), .R1(c_inv_c_3), 
           .R0(c_inv_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[44:57])
    defparam lat_alu_14.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_14.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_14.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_14.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_14.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_14.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_14.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_14.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_14.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_14.REG_FLAG_CLK = "NONE";
    defparam lat_alu_14.REG_FLAG_CE = "CE0";
    defparam lat_alu_14.REG_FLAG_RST = "RST0";
    defparam lat_alu_14.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_14.MASK01 = "0x00000000000000";
    defparam lat_alu_14.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_14.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_14.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_14.CLK0_DIV = "ENABLED";
    defparam lat_alu_14.CLK1_DIV = "ENABLED";
    defparam lat_alu_14.CLK2_DIV = "ENABLED";
    defparam lat_alu_14.CLK3_DIV = "ENABLED";
    defparam lat_alu_14.MCPAT = "0x00000000000000";
    defparam lat_alu_14.MASKPAT = "0x00000000000000";
    defparam lat_alu_14.RNDPAT = "0x00000000000000";
    defparam lat_alu_14.GSR = "DISABLED";
    defparam lat_alu_14.RESETMODE = "SYNC";
    defparam lat_alu_14.MULT9_MODE = "DISABLED";
    defparam lat_alu_14.LEGACY = "DISABLED";
    ALU54B lat_alu_13 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10432), .SIGNEDIB(n10505), .SIGNEDCIN(GND_net), 
           .A35(n10431), .A34(n10430), .A33(n10429), .A32(n10428), .A31(n10427), 
           .A30(n10426), .A29(n10425), .A28(n10424), .A27(n10423), .A26(n10422), 
           .A25(n10421), .A24(n10420), .A23(n10419), .A22(n10418), .A21(n10417), 
           .A20(n10416), .A19(n10415), .A18(n10414), .A17(n10413), .A16(n10412), 
           .A15(n10411), .A14(n10410), .A13(n10409), .A12(n10408), .A11(n10407), 
           .A10(n10406), .A9(n10405), .A8(n10404), .A7(n10403), .A6(n10402), 
           .A5(n10401), .A4(n10400), .A3(n10399), .A2(n10398), .A1(n10397), 
           .A0(n10396), .B35(n10504), .B34(n10503), .B33(n10502), .B32(n10501), 
           .B31(n10500), .B30(n10499), .B29(n10498), .B28(n10497), .B27(n10496), 
           .B26(n10495), .B25(n10494), .B24(n10493), .B23(n10492), .B22(n10491), 
           .B21(n10490), .B20(n10489), .B19(n10488), .B18(n10487), .B17(n10486), 
           .B16(n10485), .B15(n10484), .B14(n10483), .B13(n10482), .B12(n10481), 
           .B11(n10480), .B10(n10479), .B9(n10478), .B8(n10477), .B7(n10476), 
           .B6(n10475), .B5(n10474), .B4(n10473), .B3(n10472), .B2(n10471), 
           .B1(n10470), .B0(n10469), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10468), .MA34(n10467), .MA33(n10466), .MA32(n10465), 
           .MA31(n10464), .MA30(n10463), .MA29(n10462), .MA28(n10461), 
           .MA27(n10460), .MA26(n10459), .MA25(n10458), .MA24(n10457), 
           .MA23(n10456), .MA22(n10455), .MA21(n10454), .MA20(n10453), 
           .MA19(n10452), .MA18(n10451), .MA17(n10450), .MA16(n10449), 
           .MA15(n10448), .MA14(n10447), .MA13(n10446), .MA12(n10445), 
           .MA11(n10444), .MA10(n10443), .MA9(n10442), .MA8(n10441), 
           .MA7(n10440), .MA6(n10439), .MA5(n10438), .MA4(n10437), .MA3(n10436), 
           .MA2(n10435), .MA1(n10434), .MA0(n10433), .MB35(n10541), 
           .MB34(n10540), .MB33(n10539), .MB32(n10538), .MB31(n10537), 
           .MB30(n10536), .MB29(n10535), .MB28(n10534), .MB27(n10533), 
           .MB26(n10532), .MB25(n10531), .MB24(n10530), .MB23(n10529), 
           .MB22(n10528), .MB21(n10527), .MB20(n10526), .MB19(n10525), 
           .MB18(n10524), .MB17(n10523), .MB16(n10522), .MB15(n10521), 
           .MB14(n10520), .MB13(n10519), .MB12(n10518), .MB11(n10517), 
           .MB10(n10516), .MB9(n10515), .MB8(n10514), .MB7(n10513), 
           .MB6(n10512), .MB5(n10511), .MB4(n10510), .MB3(n10509), .MB2(n10508), 
           .MB1(n10507), .MB0(n10506), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n10723), 
           .R52(n10722), .R51(n10721), .R50(n10720), .R49(n10719), .R48(n10718), 
           .R47(n10717), .R46(n10716), .R45(n10715), .R44(n10714), .R43(n10713), 
           .R42(n10712), .R41(n10711), .R40(n10710), .R39(n10709), .R38(n10708), 
           .R37(n10707), .R36(n10706), .R35(n10705), .R34(n10704), .R33(n10703), 
           .R32(n10702), .R31(n10701), .R30(n10700), .R29(n10699), .R28(n10698), 
           .R27(n10697), .R26(n10696), .R25(n10695), .R24(n10694), .R23(n10693), 
           .R22(n10692), .R21(n10691), .R20(n10690), .R19(n10689), .R18(n10688), 
           .R17(c_inv_c_1), .R16(c_inv_c_0), .R15(n10380), .R14(n10381), 
           .R13(n10382), .R12(n10383), .R11(n10384), .R10(n10385), .R9(n10386), 
           .R8(n10387), .R7(n10388), .R6(n10389), .R5(n10390), .R4(n10391), 
           .R3(n10392), .R2(n10393), .R1(n10394), .R0(n10395), .SIGNEDR(n10724));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[44:57])
    defparam lat_alu_13.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_13.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_13.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_13.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_13.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_13.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_13.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_13.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_13.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_13.REG_FLAG_CLK = "NONE";
    defparam lat_alu_13.REG_FLAG_CE = "CE0";
    defparam lat_alu_13.REG_FLAG_RST = "RST0";
    defparam lat_alu_13.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_13.MASK01 = "0x00000000000000";
    defparam lat_alu_13.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_13.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_13.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_13.CLK0_DIV = "ENABLED";
    defparam lat_alu_13.CLK1_DIV = "ENABLED";
    defparam lat_alu_13.CLK2_DIV = "ENABLED";
    defparam lat_alu_13.CLK3_DIV = "ENABLED";
    defparam lat_alu_13.MCPAT = "0x00000000000000";
    defparam lat_alu_13.MASKPAT = "0x00000000000000";
    defparam lat_alu_13.RNDPAT = "0x00000000000000";
    defparam lat_alu_13.GSR = "DISABLED";
    defparam lat_alu_13.RESETMODE = "SYNC";
    defparam lat_alu_13.MULT9_MODE = "DISABLED";
    defparam lat_alu_13.LEGACY = "DISABLED";
    MULT18X18D lat_mult_12 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[16]), .B14(c_s[16]), .B13(c_s[16]), .B12(c_s[16]), 
            .B11(c_s[16]), .B10(c_s[16]), .B9(c_s[16]), .B8(c_s[16]), 
            .B7(c_s[16]), .B6(c_s[16]), .B5(c_s[16]), .B4(c_s[16]), 
            .B3(c_s[16]), .B2(c_s[16]), .B1(c_s[16]), .B0(c_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10632), .ROA16(n10631), 
            .ROA15(n10630), .ROA14(n10629), .ROA13(n10628), .ROA12(n10627), 
            .ROA11(n10626), .ROA10(n10625), .ROA9(n10624), .ROA8(n10623), 
            .ROA7(n10622), .ROA6(n10621), .ROA5(n10620), .ROA4(n10619), 
            .ROA3(n10618), .ROA2(n10617), .ROA1(n10616), .ROA0(n10615), 
            .ROB17(n10650), .ROB16(n10649), .ROB15(n10648), .ROB14(n10647), 
            .ROB13(n10646), .ROB12(n10645), .ROB11(n10644), .ROB10(n10643), 
            .ROB9(n10642), .ROB8(n10641), .ROB7(n10640), .ROB6(n10639), 
            .ROB5(n10638), .ROB4(n10637), .ROB3(n10636), .ROB2(n10635), 
            .ROB1(n10634), .ROB0(n10633), .P35(n10687), .P34(n10686), 
            .P33(n10685), .P32(n10684), .P31(n10683), .P30(n10682), 
            .P29(n10681), .P28(n10680), .P27(n10679), .P26(n10678), 
            .P25(n10677), .P24(n10676), .P23(n10675), .P22(n10674), 
            .P21(n10673), .P20(n10672), .P19(n10671), .P18(n10670), 
            .P17(n10669), .P16(n10668), .P15(n10667), .P14(n10666), 
            .P13(n10665), .P12(n10664), .P11(n10663), .P10(n10662), 
            .P9(n10661), .P8(n10660), .P7(n10659), .P6(n10658), .P5(n10657), 
            .P4(n10656), .P3(n10655), .P2(n10654), .P1(n10653), .P0(n10652), 
            .SIGNEDP(n10651));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[44:57])
    defparam lat_mult_12.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_12.REG_INPUTA_CE = "CE3";
    defparam lat_mult_12.REG_INPUTA_RST = "RST3";
    defparam lat_mult_12.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTB_CE = "CE0";
    defparam lat_mult_12.REG_INPUTB_RST = "RST0";
    defparam lat_mult_12.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_12.REG_INPUTC_CE = "CE0";
    defparam lat_mult_12.REG_INPUTC_RST = "RST0";
    defparam lat_mult_12.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_12.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_12.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_12.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_12.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_12.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_12.CLK0_DIV = "ENABLED";
    defparam lat_mult_12.CLK1_DIV = "ENABLED";
    defparam lat_mult_12.CLK2_DIV = "ENABLED";
    defparam lat_mult_12.CLK3_DIV = "ENABLED";
    defparam lat_mult_12.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_12.GSR = "DISABLED";
    defparam lat_mult_12.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_12.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_12.MULT_BYPASS = "DISABLED";
    defparam lat_mult_12.RESETMODE = "ASYNC";
    LUT4 i1446_2_lut_4_lut (.A(n68_adj_377), .B(n68_adj_345), .C(n2273), 
         .D(det_zero), .Z(n61)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1446_2_lut_4_lut.init = 16'h0035;
    MULT18X18D lat_mult_11 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[16]), .B14(c_s[16]), .B13(c_s[16]), .B12(c_s[16]), 
            .B11(c_s[16]), .B10(c_s[16]), .B9(c_s[16]), .B8(c_s[16]), 
            .B7(c_s[16]), .B6(c_s[16]), .B5(c_s[16]), .B4(c_s[16]), 
            .B3(c_s[16]), .B2(c_s[16]), .B1(c_s[16]), .B0(c_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10559), .ROA16(n10558), 
            .ROA15(n10557), .ROA14(n10556), .ROA13(n10555), .ROA12(n10554), 
            .ROA11(n10553), .ROA10(n10552), .ROA9(n10551), .ROA8(n10550), 
            .ROA7(n10549), .ROA6(n10548), .ROA5(n10547), .ROA4(n10546), 
            .ROA3(n10545), .ROA2(n10544), .ROA1(n10543), .ROA0(n10542), 
            .ROB17(n10577), .ROB16(n10576), .ROB15(n10575), .ROB14(n10574), 
            .ROB13(n10573), .ROB12(n10572), .ROB11(n10571), .ROB10(n10570), 
            .ROB9(n10569), .ROB8(n10568), .ROB7(n10567), .ROB6(n10566), 
            .ROB5(n10565), .ROB4(n10564), .ROB3(n10563), .ROB2(n10562), 
            .ROB1(n10561), .ROB0(n10560), .P35(n10614), .P34(n10613), 
            .P33(n10612), .P32(n10611), .P31(n10610), .P30(n10609), 
            .P29(n10608), .P28(n10607), .P27(n10606), .P26(n10605), 
            .P25(n10604), .P24(n10603), .P23(n10602), .P22(n10601), 
            .P21(n10600), .P20(n10599), .P19(n10598), .P18(n10597), 
            .P17(n10596), .P16(n10595), .P15(n10594), .P14(n10593), 
            .P13(n10592), .P12(n10591), .P11(n10590), .P10(n10589), 
            .P9(n10588), .P8(n10587), .P7(n10586), .P6(n10585), .P5(n10584), 
            .P4(n10583), .P3(n10582), .P2(n10581), .P1(n10580), .P0(n10579), 
            .SIGNEDP(n10578));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[44:57])
    defparam lat_mult_11.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_11.REG_INPUTA_CE = "CE3";
    defparam lat_mult_11.REG_INPUTA_RST = "RST3";
    defparam lat_mult_11.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTB_CE = "CE0";
    defparam lat_mult_11.REG_INPUTB_RST = "RST0";
    defparam lat_mult_11.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_11.REG_INPUTC_CE = "CE0";
    defparam lat_mult_11.REG_INPUTC_RST = "RST0";
    defparam lat_mult_11.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_11.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_11.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_11.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_11.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_11.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_11.CLK0_DIV = "ENABLED";
    defparam lat_mult_11.CLK1_DIV = "ENABLED";
    defparam lat_mult_11.CLK2_DIV = "ENABLED";
    defparam lat_mult_11.CLK3_DIV = "ENABLED";
    defparam lat_mult_11.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_11.GSR = "DISABLED";
    defparam lat_mult_11.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_11.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_11.MULT_BYPASS = "DISABLED";
    defparam lat_mult_11.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_10 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[15]), .B14(c_s[14]), .B13(c_s[13]), .B12(c_s[12]), 
            .B11(c_s[11]), .B10(c_s[10]), .B9(c_s[9]), .B8(c_s[8]), 
            .B7(c_s[7]), .B6(c_s[6]), .B5(c_s[5]), .B4(c_s[4]), .B3(c_s[3]), 
            .B2(c_s[2]), .B1(c_s[1]), .B0(c_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10486), .ROA16(n10485), .ROA15(n10484), .ROA14(n10483), 
            .ROA13(n10482), .ROA12(n10481), .ROA11(n10480), .ROA10(n10479), 
            .ROA9(n10478), .ROA8(n10477), .ROA7(n10476), .ROA6(n10475), 
            .ROA5(n10474), .ROA4(n10473), .ROA3(n10472), .ROA2(n10471), 
            .ROA1(n10470), .ROA0(n10469), .ROB17(n10504), .ROB16(n10503), 
            .ROB15(n10502), .ROB14(n10501), .ROB13(n10500), .ROB12(n10499), 
            .ROB11(n10498), .ROB10(n10497), .ROB9(n10496), .ROB8(n10495), 
            .ROB7(n10494), .ROB6(n10493), .ROB5(n10492), .ROB4(n10491), 
            .ROB3(n10490), .ROB2(n10489), .ROB1(n10488), .ROB0(n10487), 
            .P35(n10541), .P34(n10540), .P33(n10539), .P32(n10538), 
            .P31(n10537), .P30(n10536), .P29(n10535), .P28(n10534), 
            .P27(n10533), .P26(n10532), .P25(n10531), .P24(n10530), 
            .P23(n10529), .P22(n10528), .P21(n10527), .P20(n10526), 
            .P19(n10525), .P18(n10524), .P17(n10523), .P16(n10522), 
            .P15(n10521), .P14(n10520), .P13(n10519), .P12(n10518), 
            .P11(n10517), .P10(n10516), .P9(n10515), .P8(n10514), .P7(n10513), 
            .P6(n10512), .P5(n10511), .P4(n10510), .P3(n10509), .P2(n10508), 
            .P1(n10507), .P0(n10506), .SIGNEDP(n10505));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[44:57])
    defparam lat_mult_10.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_10.REG_INPUTA_CE = "CE3";
    defparam lat_mult_10.REG_INPUTA_RST = "RST3";
    defparam lat_mult_10.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTB_CE = "CE0";
    defparam lat_mult_10.REG_INPUTB_RST = "RST0";
    defparam lat_mult_10.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_10.REG_INPUTC_CE = "CE0";
    defparam lat_mult_10.REG_INPUTC_RST = "RST0";
    defparam lat_mult_10.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_10.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_10.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_10.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_10.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_10.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_10.CLK0_DIV = "ENABLED";
    defparam lat_mult_10.CLK1_DIV = "ENABLED";
    defparam lat_mult_10.CLK2_DIV = "ENABLED";
    defparam lat_mult_10.CLK3_DIV = "ENABLED";
    defparam lat_mult_10.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_10.GSR = "DISABLED";
    defparam lat_mult_10.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_10.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_10.MULT_BYPASS = "DISABLED";
    defparam lat_mult_10.RESETMODE = "ASYNC";
    MULT18X18D c_s_31__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(c_s[16]), .B16(c_s[16]), 
            .B15(c_s[15]), .B14(c_s[14]), .B13(c_s[13]), .B12(c_s[12]), 
            .B11(c_s[11]), .B10(c_s[10]), .B9(c_s[9]), .B8(c_s[8]), 
            .B7(c_s[7]), .B6(c_s[6]), .B5(c_s[5]), .B4(c_s[4]), .B3(c_s[3]), 
            .B2(c_s[2]), .B1(c_s[1]), .B0(c_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10413), .ROA16(n10412), .ROA15(n10411), .ROA14(n10410), 
            .ROA13(n10409), .ROA12(n10408), .ROA11(n10407), .ROA10(n10406), 
            .ROA9(n10405), .ROA8(n10404), .ROA7(n10403), .ROA6(n10402), 
            .ROA5(n10401), .ROA4(n10400), .ROA3(n10399), .ROA2(n10398), 
            .ROA1(n10397), .ROA0(n10396), .ROB17(n10431), .ROB16(n10430), 
            .ROB15(n10429), .ROB14(n10428), .ROB13(n10427), .ROB12(n10426), 
            .ROB11(n10425), .ROB10(n10424), .ROB9(n10423), .ROB8(n10422), 
            .ROB7(n10421), .ROB6(n10420), .ROB5(n10419), .ROB4(n10418), 
            .ROB3(n10417), .ROB2(n10416), .ROB1(n10415), .ROB0(n10414), 
            .P35(n10468), .P34(n10467), .P33(n10466), .P32(n10465), 
            .P31(n10464), .P30(n10463), .P29(n10462), .P28(n10461), 
            .P27(n10460), .P26(n10459), .P25(n10458), .P24(n10457), 
            .P23(n10456), .P22(n10455), .P21(n10454), .P20(n10453), 
            .P19(n10452), .P18(n10451), .P17(n10450), .P16(n10449), 
            .P15(n10448), .P14(n10447), .P13(n10446), .P12(n10445), 
            .P11(n10444), .P10(n10443), .P9(n10442), .P8(n10441), .P7(n10440), 
            .P6(n10439), .P5(n10438), .P4(n10437), .P3(n10436), .P2(n10435), 
            .P1(n10434), .P0(n10433), .SIGNEDP(n10432));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(86[44:57])
    defparam c_s_31__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam c_s_31__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam c_s_31__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam c_s_31__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam c_s_31__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam c_s_31__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam c_s_31__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam c_s_31__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam c_s_31__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam c_s_31__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam c_s_31__I_0_mult_2.GSR = "DISABLED";
    defparam c_s_31__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam c_s_31__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam c_s_31__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam c_s_31__I_0_mult_2.RESETMODE = "ASYNC";
    ALU54B lat_alu_9 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10201), .SIGNEDIB(n10274), .SIGNEDCIN(n10347), .A35(n10200), 
           .A34(n10199), .A33(n10198), .A32(n10197), .A31(n10196), .A30(n10195), 
           .A29(n10194), .A28(n10193), .A27(n10192), .A26(n10191), .A25(n10190), 
           .A24(n10189), .A23(n10188), .A22(n10187), .A21(n10186), .A20(n10185), 
           .A19(n10184), .A18(n10183), .A17(n10182), .A16(n10181), .A15(n10180), 
           .A14(n10179), .A13(n10178), .A12(n10177), .A11(n10176), .A10(n10175), 
           .A9(n10174), .A8(n10173), .A7(n10172), .A6(n10171), .A5(n10170), 
           .A4(n10169), .A3(n10168), .A2(n10167), .A1(n10166), .A0(n10165), 
           .B35(n10273), .B34(n10272), .B33(n10271), .B32(n10270), .B31(n10269), 
           .B30(n10268), .B29(n10267), .B28(n10266), .B27(n10265), .B26(n10264), 
           .B25(n10263), .B24(n10262), .B23(n10261), .B22(n10260), .B21(n10259), 
           .B20(n10258), .B19(n10257), .B18(n10256), .B17(n10255), .B16(n10254), 
           .B15(n10253), .B14(n10252), .B13(n10251), .B12(n10250), .B11(n10249), 
           .B10(n10248), .B9(n10247), .B8(n10246), .B7(n10245), .B6(n10244), 
           .B5(n10243), .B4(n10242), .B3(n10241), .B2(n10240), .B1(n10239), 
           .B0(n10238), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10237), .MA34(n10236), .MA33(n10235), .MA32(n10234), 
           .MA31(n10233), .MA30(n10232), .MA29(n10231), .MA28(n10230), 
           .MA27(n10229), .MA26(n10228), .MA25(n10227), .MA24(n10226), 
           .MA23(n10225), .MA22(n10224), .MA21(n10223), .MA20(n10222), 
           .MA19(n10221), .MA18(n10220), .MA17(n10219), .MA16(n10218), 
           .MA15(n10217), .MA14(n10216), .MA13(n10215), .MA12(n10214), 
           .MA11(n10213), .MA10(n10212), .MA9(n10211), .MA8(n10210), 
           .MA7(n10209), .MA6(n10208), .MA5(n10207), .MA4(n10206), .MA3(n10205), 
           .MA2(n10204), .MA1(n10203), .MA0(n10202), .MB35(n10310), 
           .MB34(n10309), .MB33(n10308), .MB32(n10307), .MB31(n10306), 
           .MB30(n10305), .MB29(n10304), .MB28(n10303), .MB27(n10302), 
           .MB26(n10301), .MB25(n10300), .MB24(n10299), .MB23(n10298), 
           .MB22(n10297), .MB21(n10296), .MB20(n10295), .MB19(n10294), 
           .MB18(n10293), .MB17(n10292), .MB16(n10291), .MB15(n10290), 
           .MB14(n10289), .MB13(n10288), .MB12(n10287), .MB11(n10286), 
           .MB10(n10285), .MB9(n10284), .MB8(n10283), .MB7(n10282), 
           .MB6(n10281), .MB5(n10280), .MB4(n10279), .MB3(n10278), .MB2(n10277), 
           .MB1(n10276), .MB0(n10275), .CIN53(n10346), .CIN52(n10345), 
           .CIN51(n10344), .CIN50(n10343), .CIN49(n10342), .CIN48(n10341), 
           .CIN47(n10340), .CIN46(n10339), .CIN45(n10338), .CIN44(n10337), 
           .CIN43(n10336), .CIN42(n10335), .CIN41(n10334), .CIN40(n10333), 
           .CIN39(n10332), .CIN38(n10331), .CIN37(n10330), .CIN36(n10329), 
           .CIN35(n10328), .CIN34(n10327), .CIN33(n10326), .CIN32(n10325), 
           .CIN31(n10324), .CIN30(n10323), .CIN29(n10322), .CIN28(n10321), 
           .CIN27(n10320), .CIN26(n10319), .CIN25(n10318), .CIN24(n10317), 
           .CIN23(n10316), .CIN22(n10315), .CIN21(n10314), .CIN20(n10313), 
           .CIN19(n10312), .CIN18(n10311), .CIN17(b_inv_c_1), .CIN16(b_inv_c_0), 
           .CIN15(n10003), .CIN14(n10004), .CIN13(n10005), .CIN12(n10006), 
           .CIN11(n10007), .CIN10(n10008), .CIN9(n10009), .CIN8(n10010), 
           .CIN7(n10011), .CIN6(n10012), .CIN5(n10013), .CIN4(n10014), 
           .CIN3(n10015), .CIN2(n10016), .CIN1(n10017), .CIN0(n10018), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R13(prod_b[31]), 
           .R12(prod_b[30]), .R11(prod_b[29]), .R10(b_inv_c_12), .R9(b_inv_c_11), 
           .R8(b_inv_c_10), .R7(b_inv_c_9), .R6(b_inv_c_8), .R5(b_inv_c_7), 
           .R4(b_inv_c_6), .R3(b_inv_c_5), .R2(b_inv_c_4), .R1(b_inv_c_3), 
           .R0(b_inv_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[44:57])
    defparam lat_alu_9.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_9.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_9.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_9.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_9.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_9.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_9.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_9.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_9.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_9.REG_FLAG_CLK = "NONE";
    defparam lat_alu_9.REG_FLAG_CE = "CE0";
    defparam lat_alu_9.REG_FLAG_RST = "RST0";
    defparam lat_alu_9.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_9.MASK01 = "0x00000000000000";
    defparam lat_alu_9.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_9.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_9.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_9.CLK0_DIV = "ENABLED";
    defparam lat_alu_9.CLK1_DIV = "ENABLED";
    defparam lat_alu_9.CLK2_DIV = "ENABLED";
    defparam lat_alu_9.CLK3_DIV = "ENABLED";
    defparam lat_alu_9.MCPAT = "0x00000000000000";
    defparam lat_alu_9.MASKPAT = "0x00000000000000";
    defparam lat_alu_9.RNDPAT = "0x00000000000000";
    defparam lat_alu_9.GSR = "DISABLED";
    defparam lat_alu_9.RESETMODE = "SYNC";
    defparam lat_alu_9.MULT9_MODE = "DISABLED";
    defparam lat_alu_9.LEGACY = "DISABLED";
    LUT4 i334_3_lut (.A(prod_d[31]), .B(prod_d[30]), .C(prod_d[29]), .Z(d_inv_c_15)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i334_3_lut.init = 16'h6a6a;
    ALU54B lat_alu_8 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n10055), .SIGNEDIB(n10128), .SIGNEDCIN(GND_net), 
           .A35(n10054), .A34(n10053), .A33(n10052), .A32(n10051), .A31(n10050), 
           .A30(n10049), .A29(n10048), .A28(n10047), .A27(n10046), .A26(n10045), 
           .A25(n10044), .A24(n10043), .A23(n10042), .A22(n10041), .A21(n10040), 
           .A20(n10039), .A19(n10038), .A18(n10037), .A17(n10036), .A16(n10035), 
           .A15(n10034), .A14(n10033), .A13(n10032), .A12(n10031), .A11(n10030), 
           .A10(n10029), .A9(n10028), .A8(n10027), .A7(n10026), .A6(n10025), 
           .A5(n10024), .A4(n10023), .A3(n10022), .A2(n10021), .A1(n10020), 
           .A0(n10019), .B35(n10127), .B34(n10126), .B33(n10125), .B32(n10124), 
           .B31(n10123), .B30(n10122), .B29(n10121), .B28(n10120), .B27(n10119), 
           .B26(n10118), .B25(n10117), .B24(n10116), .B23(n10115), .B22(n10114), 
           .B21(n10113), .B20(n10112), .B19(n10111), .B18(n10110), .B17(n10109), 
           .B16(n10108), .B15(n10107), .B14(n10106), .B13(n10105), .B12(n10104), 
           .B11(n10103), .B10(n10102), .B9(n10101), .B8(n10100), .B7(n10099), 
           .B6(n10098), .B5(n10097), .B4(n10096), .B3(n10095), .B2(n10094), 
           .B1(n10093), .B0(n10092), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n10091), .MA34(n10090), .MA33(n10089), .MA32(n10088), 
           .MA31(n10087), .MA30(n10086), .MA29(n10085), .MA28(n10084), 
           .MA27(n10083), .MA26(n10082), .MA25(n10081), .MA24(n10080), 
           .MA23(n10079), .MA22(n10078), .MA21(n10077), .MA20(n10076), 
           .MA19(n10075), .MA18(n10074), .MA17(n10073), .MA16(n10072), 
           .MA15(n10071), .MA14(n10070), .MA13(n10069), .MA12(n10068), 
           .MA11(n10067), .MA10(n10066), .MA9(n10065), .MA8(n10064), 
           .MA7(n10063), .MA6(n10062), .MA5(n10061), .MA4(n10060), .MA3(n10059), 
           .MA2(n10058), .MA1(n10057), .MA0(n10056), .MB35(n10164), 
           .MB34(n10163), .MB33(n10162), .MB32(n10161), .MB31(n10160), 
           .MB30(n10159), .MB29(n10158), .MB28(n10157), .MB27(n10156), 
           .MB26(n10155), .MB25(n10154), .MB24(n10153), .MB23(n10152), 
           .MB22(n10151), .MB21(n10150), .MB20(n10149), .MB19(n10148), 
           .MB18(n10147), .MB17(n10146), .MB16(n10145), .MB15(n10144), 
           .MB14(n10143), .MB13(n10142), .MB12(n10141), .MB11(n10140), 
           .MB10(n10139), .MB9(n10138), .MB8(n10137), .MB7(n10136), 
           .MB6(n10135), .MB5(n10134), .MB4(n10133), .MB3(n10132), .MB2(n10131), 
           .MB1(n10130), .MB0(n10129), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n10346), 
           .R52(n10345), .R51(n10344), .R50(n10343), .R49(n10342), .R48(n10341), 
           .R47(n10340), .R46(n10339), .R45(n10338), .R44(n10337), .R43(n10336), 
           .R42(n10335), .R41(n10334), .R40(n10333), .R39(n10332), .R38(n10331), 
           .R37(n10330), .R36(n10329), .R35(n10328), .R34(n10327), .R33(n10326), 
           .R32(n10325), .R31(n10324), .R30(n10323), .R29(n10322), .R28(n10321), 
           .R27(n10320), .R26(n10319), .R25(n10318), .R24(n10317), .R23(n10316), 
           .R22(n10315), .R21(n10314), .R20(n10313), .R19(n10312), .R18(n10311), 
           .R17(b_inv_c_1), .R16(b_inv_c_0), .R15(n10003), .R14(n10004), 
           .R13(n10005), .R12(n10006), .R11(n10007), .R10(n10008), .R9(n10009), 
           .R8(n10010), .R7(n10011), .R6(n10012), .R5(n10013), .R4(n10014), 
           .R3(n10015), .R2(n10016), .R1(n10017), .R0(n10018), .SIGNEDR(n10347));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[44:57])
    defparam lat_alu_8.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_8.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_8.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_8.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_8.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_8.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_8.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_8.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_8.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_8.REG_FLAG_CLK = "NONE";
    defparam lat_alu_8.REG_FLAG_CE = "CE0";
    defparam lat_alu_8.REG_FLAG_RST = "RST0";
    defparam lat_alu_8.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_8.MASK01 = "0x00000000000000";
    defparam lat_alu_8.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_8.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_8.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_8.CLK0_DIV = "ENABLED";
    defparam lat_alu_8.CLK1_DIV = "ENABLED";
    defparam lat_alu_8.CLK2_DIV = "ENABLED";
    defparam lat_alu_8.CLK3_DIV = "ENABLED";
    defparam lat_alu_8.MCPAT = "0x00000000000000";
    defparam lat_alu_8.MASKPAT = "0x00000000000000";
    defparam lat_alu_8.RNDPAT = "0x00000000000000";
    defparam lat_alu_8.GSR = "DISABLED";
    defparam lat_alu_8.RESETMODE = "SYNC";
    defparam lat_alu_8.MULT9_MODE = "DISABLED";
    defparam lat_alu_8.LEGACY = "DISABLED";
    MULT18X18D lat_mult_7 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[16]), .B14(b_s[16]), .B13(b_s[16]), .B12(b_s[16]), 
            .B11(b_s[16]), .B10(b_s[16]), .B9(b_s[16]), .B8(b_s[16]), 
            .B7(b_s[16]), .B6(b_s[16]), .B5(b_s[16]), .B4(b_s[16]), 
            .B3(b_s[16]), .B2(b_s[16]), .B1(b_s[16]), .B0(b_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10255), .ROA16(n10254), 
            .ROA15(n10253), .ROA14(n10252), .ROA13(n10251), .ROA12(n10250), 
            .ROA11(n10249), .ROA10(n10248), .ROA9(n10247), .ROA8(n10246), 
            .ROA7(n10245), .ROA6(n10244), .ROA5(n10243), .ROA4(n10242), 
            .ROA3(n10241), .ROA2(n10240), .ROA1(n10239), .ROA0(n10238), 
            .ROB17(n10273), .ROB16(n10272), .ROB15(n10271), .ROB14(n10270), 
            .ROB13(n10269), .ROB12(n10268), .ROB11(n10267), .ROB10(n10266), 
            .ROB9(n10265), .ROB8(n10264), .ROB7(n10263), .ROB6(n10262), 
            .ROB5(n10261), .ROB4(n10260), .ROB3(n10259), .ROB2(n10258), 
            .ROB1(n10257), .ROB0(n10256), .P35(n10310), .P34(n10309), 
            .P33(n10308), .P32(n10307), .P31(n10306), .P30(n10305), 
            .P29(n10304), .P28(n10303), .P27(n10302), .P26(n10301), 
            .P25(n10300), .P24(n10299), .P23(n10298), .P22(n10297), 
            .P21(n10296), .P20(n10295), .P19(n10294), .P18(n10293), 
            .P17(n10292), .P16(n10291), .P15(n10290), .P14(n10289), 
            .P13(n10288), .P12(n10287), .P11(n10286), .P10(n10285), 
            .P9(n10284), .P8(n10283), .P7(n10282), .P6(n10281), .P5(n10280), 
            .P4(n10279), .P3(n10278), .P2(n10277), .P1(n10276), .P0(n10275), 
            .SIGNEDP(n10274));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[44:57])
    defparam lat_mult_7.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_7.REG_INPUTA_CE = "CE3";
    defparam lat_mult_7.REG_INPUTA_RST = "RST3";
    defparam lat_mult_7.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTB_CE = "CE0";
    defparam lat_mult_7.REG_INPUTB_RST = "RST0";
    defparam lat_mult_7.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_7.REG_INPUTC_CE = "CE0";
    defparam lat_mult_7.REG_INPUTC_RST = "RST0";
    defparam lat_mult_7.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_7.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_7.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_7.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_7.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_7.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_7.CLK0_DIV = "ENABLED";
    defparam lat_mult_7.CLK1_DIV = "ENABLED";
    defparam lat_mult_7.CLK2_DIV = "ENABLED";
    defparam lat_mult_7.CLK3_DIV = "ENABLED";
    defparam lat_mult_7.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_7.GSR = "DISABLED";
    defparam lat_mult_7.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_7.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_7.MULT_BYPASS = "DISABLED";
    defparam lat_mult_7.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_6 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[16]), .B14(b_s[16]), .B13(b_s[16]), .B12(b_s[16]), 
            .B11(b_s[16]), .B10(b_s[16]), .B9(b_s[16]), .B8(b_s[16]), 
            .B7(b_s[16]), .B6(b_s[16]), .B5(b_s[16]), .B4(b_s[16]), 
            .B3(b_s[16]), .B2(b_s[16]), .B1(b_s[16]), .B0(b_s[16]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n10182), .ROA16(n10181), 
            .ROA15(n10180), .ROA14(n10179), .ROA13(n10178), .ROA12(n10177), 
            .ROA11(n10176), .ROA10(n10175), .ROA9(n10174), .ROA8(n10173), 
            .ROA7(n10172), .ROA6(n10171), .ROA5(n10170), .ROA4(n10169), 
            .ROA3(n10168), .ROA2(n10167), .ROA1(n10166), .ROA0(n10165), 
            .ROB17(n10200), .ROB16(n10199), .ROB15(n10198), .ROB14(n10197), 
            .ROB13(n10196), .ROB12(n10195), .ROB11(n10194), .ROB10(n10193), 
            .ROB9(n10192), .ROB8(n10191), .ROB7(n10190), .ROB6(n10189), 
            .ROB5(n10188), .ROB4(n10187), .ROB3(n10186), .ROB2(n10185), 
            .ROB1(n10184), .ROB0(n10183), .P35(n10237), .P34(n10236), 
            .P33(n10235), .P32(n10234), .P31(n10233), .P30(n10232), 
            .P29(n10231), .P28(n10230), .P27(n10229), .P26(n10228), 
            .P25(n10227), .P24(n10226), .P23(n10225), .P22(n10224), 
            .P21(n10223), .P20(n10222), .P19(n10221), .P18(n10220), 
            .P17(n10219), .P16(n10218), .P15(n10217), .P14(n10216), 
            .P13(n10215), .P12(n10214), .P11(n10213), .P10(n10212), 
            .P9(n10211), .P8(n10210), .P7(n10209), .P6(n10208), .P5(n10207), 
            .P4(n10206), .P3(n10205), .P2(n10204), .P1(n10203), .P0(n10202), 
            .SIGNEDP(n10201));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[44:57])
    defparam lat_mult_6.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_6.REG_INPUTA_CE = "CE3";
    defparam lat_mult_6.REG_INPUTA_RST = "RST3";
    defparam lat_mult_6.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTB_CE = "CE0";
    defparam lat_mult_6.REG_INPUTB_RST = "RST0";
    defparam lat_mult_6.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_6.REG_INPUTC_CE = "CE0";
    defparam lat_mult_6.REG_INPUTC_RST = "RST0";
    defparam lat_mult_6.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_6.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_6.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_6.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_6.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_6.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_6.CLK0_DIV = "ENABLED";
    defparam lat_mult_6.CLK1_DIV = "ENABLED";
    defparam lat_mult_6.CLK2_DIV = "ENABLED";
    defparam lat_mult_6.CLK3_DIV = "ENABLED";
    defparam lat_mult_6.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_6.GSR = "DISABLED";
    defparam lat_mult_6.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_6.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_6.MULT_BYPASS = "DISABLED";
    defparam lat_mult_6.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_5 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[15]), .B14(b_s[14]), .B13(b_s[13]), .B12(b_s[12]), 
            .B11(b_s[11]), .B10(b_s[10]), .B9(b_s[9]), .B8(b_s[8]), 
            .B7(b_s[7]), .B6(b_s[6]), .B5(b_s[5]), .B4(b_s[4]), .B3(b_s[3]), 
            .B2(b_s[2]), .B1(b_s[1]), .B0(b_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10109), .ROA16(n10108), .ROA15(n10107), .ROA14(n10106), 
            .ROA13(n10105), .ROA12(n10104), .ROA11(n10103), .ROA10(n10102), 
            .ROA9(n10101), .ROA8(n10100), .ROA7(n10099), .ROA6(n10098), 
            .ROA5(n10097), .ROA4(n10096), .ROA3(n10095), .ROA2(n10094), 
            .ROA1(n10093), .ROA0(n10092), .ROB17(n10127), .ROB16(n10126), 
            .ROB15(n10125), .ROB14(n10124), .ROB13(n10123), .ROB12(n10122), 
            .ROB11(n10121), .ROB10(n10120), .ROB9(n10119), .ROB8(n10118), 
            .ROB7(n10117), .ROB6(n10116), .ROB5(n10115), .ROB4(n10114), 
            .ROB3(n10113), .ROB2(n10112), .ROB1(n10111), .ROB0(n10110), 
            .P35(n10164), .P34(n10163), .P33(n10162), .P32(n10161), 
            .P31(n10160), .P30(n10159), .P29(n10158), .P28(n10157), 
            .P27(n10156), .P26(n10155), .P25(n10154), .P24(n10153), 
            .P23(n10152), .P22(n10151), .P21(n10150), .P20(n10149), 
            .P19(n10148), .P18(n10147), .P17(n10146), .P16(n10145), 
            .P15(n10144), .P14(n10143), .P13(n10142), .P12(n10141), 
            .P11(n10140), .P10(n10139), .P9(n10138), .P8(n10137), .P7(n10136), 
            .P6(n10135), .P5(n10134), .P4(n10133), .P3(n10132), .P2(n10131), 
            .P1(n10130), .P0(n10129), .SIGNEDP(n10128));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[44:57])
    defparam lat_mult_5.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_5.REG_INPUTA_CE = "CE3";
    defparam lat_mult_5.REG_INPUTA_RST = "RST3";
    defparam lat_mult_5.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTB_CE = "CE0";
    defparam lat_mult_5.REG_INPUTB_RST = "RST0";
    defparam lat_mult_5.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_5.REG_INPUTC_CE = "CE0";
    defparam lat_mult_5.REG_INPUTC_RST = "RST0";
    defparam lat_mult_5.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_5.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_5.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_5.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_5.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_5.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_5.CLK0_DIV = "ENABLED";
    defparam lat_mult_5.CLK1_DIV = "ENABLED";
    defparam lat_mult_5.CLK2_DIV = "ENABLED";
    defparam lat_mult_5.CLK3_DIV = "ENABLED";
    defparam lat_mult_5.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_5.GSR = "DISABLED";
    defparam lat_mult_5.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_5.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_5.MULT_BYPASS = "DISABLED";
    defparam lat_mult_5.RESETMODE = "ASYNC";
    MULT18X18D b_s_31__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(b_s[16]), .B16(b_s[16]), 
            .B15(b_s[15]), .B14(b_s[14]), .B13(b_s[13]), .B12(b_s[12]), 
            .B11(b_s[11]), .B10(b_s[10]), .B9(b_s[9]), .B8(b_s[8]), 
            .B7(b_s[7]), .B6(b_s[6]), .B5(b_s[5]), .B4(b_s[4]), .B3(b_s[3]), 
            .B2(b_s[2]), .B1(b_s[1]), .B0(b_s[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n10036), .ROA16(n10035), .ROA15(n10034), .ROA14(n10033), 
            .ROA13(n10032), .ROA12(n10031), .ROA11(n10030), .ROA10(n10029), 
            .ROA9(n10028), .ROA8(n10027), .ROA7(n10026), .ROA6(n10025), 
            .ROA5(n10024), .ROA4(n10023), .ROA3(n10022), .ROA2(n10021), 
            .ROA1(n10020), .ROA0(n10019), .ROB17(n10054), .ROB16(n10053), 
            .ROB15(n10052), .ROB14(n10051), .ROB13(n10050), .ROB12(n10049), 
            .ROB11(n10048), .ROB10(n10047), .ROB9(n10046), .ROB8(n10045), 
            .ROB7(n10044), .ROB6(n10043), .ROB5(n10042), .ROB4(n10041), 
            .ROB3(n10040), .ROB2(n10039), .ROB1(n10038), .ROB0(n10037), 
            .P35(n10091), .P34(n10090), .P33(n10089), .P32(n10088), 
            .P31(n10087), .P30(n10086), .P29(n10085), .P28(n10084), 
            .P27(n10083), .P26(n10082), .P25(n10081), .P24(n10080), 
            .P23(n10079), .P22(n10078), .P21(n10077), .P20(n10076), 
            .P19(n10075), .P18(n10074), .P17(n10073), .P16(n10072), 
            .P15(n10071), .P14(n10070), .P13(n10069), .P12(n10068), 
            .P11(n10067), .P10(n10066), .P9(n10065), .P8(n10064), .P7(n10063), 
            .P6(n10062), .P5(n10061), .P4(n10060), .P3(n10059), .P2(n10058), 
            .P1(n10057), .P0(n10056), .SIGNEDP(n10055));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(85[44:57])
    defparam b_s_31__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam b_s_31__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam b_s_31__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam b_s_31__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam b_s_31__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam b_s_31__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam b_s_31__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam b_s_31__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam b_s_31__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam b_s_31__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam b_s_31__I_0_mult_2.GSR = "DISABLED";
    defparam b_s_31__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam b_s_31__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam b_s_31__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam b_s_31__I_0_mult_2.RESETMODE = "ASYNC";
    LUT4 i391_1_lut (.A(prod_c[29]), .Z(c_inv_c_13)) /* synthesis lut_function=(!(A)) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i391_1_lut.init = 16'h5555;
    ALU54B lat_alu_4 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n9824), .SIGNEDIB(n9897), .SIGNEDCIN(n9970), .A35(n9823), 
           .A34(n9822), .A33(n9821), .A32(n9820), .A31(n9819), .A30(n9818), 
           .A29(n9817), .A28(n9816), .A27(n9815), .A26(n9814), .A25(n9813), 
           .A24(n9812), .A23(n9811), .A22(n9810), .A21(n9809), .A20(n9808), 
           .A19(n9807), .A18(n9806), .A17(n9805), .A16(n9804), .A15(n9803), 
           .A14(n9802), .A13(n9801), .A12(n9800), .A11(n9799), .A10(n9798), 
           .A9(n9797), .A8(n9796), .A7(n9795), .A6(n9794), .A5(n9793), 
           .A4(n9792), .A3(n9791), .A2(n9790), .A1(n9789), .A0(n9788), 
           .B35(n9896), .B34(n9895), .B33(n9894), .B32(n9893), .B31(n9892), 
           .B30(n9891), .B29(n9890), .B28(n9889), .B27(n9888), .B26(n9887), 
           .B25(n9886), .B24(n9885), .B23(n9884), .B22(n9883), .B21(n9882), 
           .B20(n9881), .B19(n9880), .B18(n9879), .B17(n9878), .B16(n9877), 
           .B15(n9876), .B14(n9875), .B13(n9874), .B12(n9873), .B11(n9872), 
           .B10(n9871), .B9(n9870), .B8(n9869), .B7(n9868), .B6(n9867), 
           .B5(n9866), .B4(n9865), .B3(n9864), .B2(n9863), .B1(n9862), 
           .B0(n9861), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n9860), .MA34(n9859), .MA33(n9858), .MA32(n9857), .MA31(n9856), 
           .MA30(n9855), .MA29(n9854), .MA28(n9853), .MA27(n9852), .MA26(n9851), 
           .MA25(n9850), .MA24(n9849), .MA23(n9848), .MA22(n9847), .MA21(n9846), 
           .MA20(n9845), .MA19(n9844), .MA18(n9843), .MA17(n9842), .MA16(n9841), 
           .MA15(n9840), .MA14(n9839), .MA13(n9838), .MA12(n9837), .MA11(n9836), 
           .MA10(n9835), .MA9(n9834), .MA8(n9833), .MA7(n9832), .MA6(n9831), 
           .MA5(n9830), .MA4(n9829), .MA3(n9828), .MA2(n9827), .MA1(n9826), 
           .MA0(n9825), .MB35(n9933), .MB34(n9932), .MB33(n9931), .MB32(n9930), 
           .MB31(n9929), .MB30(n9928), .MB29(n9927), .MB28(n9926), .MB27(n9925), 
           .MB26(n9924), .MB25(n9923), .MB24(n9922), .MB23(n9921), .MB22(n9920), 
           .MB21(n9919), .MB20(n9918), .MB19(n9917), .MB18(n9916), .MB17(n9915), 
           .MB16(n9914), .MB15(n9913), .MB14(n9912), .MB13(n9911), .MB12(n9910), 
           .MB11(n9909), .MB10(n9908), .MB9(n9907), .MB8(n9906), .MB7(n9905), 
           .MB6(n9904), .MB5(n9903), .MB4(n9902), .MB3(n9901), .MB2(n9900), 
           .MB1(n9899), .MB0(n9898), .CIN53(n9969), .CIN52(n9968), .CIN51(n9967), 
           .CIN50(n9966), .CIN49(n9965), .CIN48(n9964), .CIN47(n9963), 
           .CIN46(n9962), .CIN45(n9961), .CIN44(n9960), .CIN43(n9959), 
           .CIN42(n9958), .CIN41(n9957), .CIN40(n9956), .CIN39(n9955), 
           .CIN38(n9954), .CIN37(n9953), .CIN36(n9952), .CIN35(n9951), 
           .CIN34(n9950), .CIN33(n9949), .CIN32(n9948), .CIN31(n9947), 
           .CIN30(n9946), .CIN29(n9945), .CIN28(n9944), .CIN27(n9943), 
           .CIN26(n9942), .CIN25(n9941), .CIN24(n9940), .CIN23(n9939), 
           .CIN22(n9938), .CIN21(n9937), .CIN20(n9936), .CIN19(n9935), 
           .CIN18(n9934), .CIN17(a_inv_c_1), .CIN16(a_inv_c_0), .CIN15(n9626), 
           .CIN14(n9627), .CIN13(n9628), .CIN12(n9629), .CIN11(n9630), 
           .CIN10(n9631), .CIN9(n9632), .CIN8(n9633), .CIN7(n9634), 
           .CIN6(n9635), .CIN5(n9636), .CIN4(n9637), .CIN3(n9638), .CIN2(n9639), 
           .CIN1(n9640), .CIN0(n9641), .OP10(GND_net), .OP9(VCC_net), 
           .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), .OP5(GND_net), 
           .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), .OP1(GND_net), 
           .OP0(VCC_net), .R13(prod_a[31]), .R12(prod_a[30]), .R11(prod_a[29]), 
           .R10(a_inv_c_12), .R9(a_inv_c_11), .R8(a_inv_c_10), .R7(a_inv_c_9), 
           .R6(a_inv_c_8), .R5(a_inv_c_7), .R4(a_inv_c_6), .R3(a_inv_c_5), 
           .R2(a_inv_c_4), .R1(a_inv_c_3), .R0(a_inv_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam lat_alu_4.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_4.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_4.REG_FLAG_CLK = "NONE";
    defparam lat_alu_4.REG_FLAG_CE = "CE0";
    defparam lat_alu_4.REG_FLAG_RST = "RST0";
    defparam lat_alu_4.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASK01 = "0x00000000000000";
    defparam lat_alu_4.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_4.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_4.CLK0_DIV = "ENABLED";
    defparam lat_alu_4.CLK1_DIV = "ENABLED";
    defparam lat_alu_4.CLK2_DIV = "ENABLED";
    defparam lat_alu_4.CLK3_DIV = "ENABLED";
    defparam lat_alu_4.MCPAT = "0x00000000000000";
    defparam lat_alu_4.MASKPAT = "0x00000000000000";
    defparam lat_alu_4.RNDPAT = "0x00000000000000";
    defparam lat_alu_4.GSR = "DISABLED";
    defparam lat_alu_4.RESETMODE = "SYNC";
    defparam lat_alu_4.MULT9_MODE = "DISABLED";
    defparam lat_alu_4.LEGACY = "DISABLED";
    ALU54B lat_alu_3 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n9678), .SIGNEDIB(n9751), .SIGNEDCIN(GND_net), .A35(n9677), 
           .A34(n9676), .A33(n9675), .A32(n9674), .A31(n9673), .A30(n9672), 
           .A29(n9671), .A28(n9670), .A27(n9669), .A26(n9668), .A25(n9667), 
           .A24(n9666), .A23(n9665), .A22(n9664), .A21(n9663), .A20(n9662), 
           .A19(n9661), .A18(n9660), .A17(n9659), .A16(n9658), .A15(n9657), 
           .A14(n9656), .A13(n9655), .A12(n9654), .A11(n9653), .A10(n9652), 
           .A9(n9651), .A8(n9650), .A7(n9649), .A6(n9648), .A5(n9647), 
           .A4(n9646), .A3(n9645), .A2(n9644), .A1(n9643), .A0(n9642), 
           .B35(n9750), .B34(n9749), .B33(n9748), .B32(n9747), .B31(n9746), 
           .B30(n9745), .B29(n9744), .B28(n9743), .B27(n9742), .B26(n9741), 
           .B25(n9740), .B24(n9739), .B23(n9738), .B22(n9737), .B21(n9736), 
           .B20(n9735), .B19(n9734), .B18(n9733), .B17(n9732), .B16(n9731), 
           .B15(n9730), .B14(n9729), .B13(n9728), .B12(n9727), .B11(n9726), 
           .B10(n9725), .B9(n9724), .B8(n9723), .B7(n9722), .B6(n9721), 
           .B5(n9720), .B4(n9719), .B3(n9718), .B2(n9717), .B1(n9716), 
           .B0(n9715), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n9714), .MA34(n9713), .MA33(n9712), .MA32(n9711), .MA31(n9710), 
           .MA30(n9709), .MA29(n9708), .MA28(n9707), .MA27(n9706), .MA26(n9705), 
           .MA25(n9704), .MA24(n9703), .MA23(n9702), .MA22(n9701), .MA21(n9700), 
           .MA20(n9699), .MA19(n9698), .MA18(n9697), .MA17(n9696), .MA16(n9695), 
           .MA15(n9694), .MA14(n9693), .MA13(n9692), .MA12(n9691), .MA11(n9690), 
           .MA10(n9689), .MA9(n9688), .MA8(n9687), .MA7(n9686), .MA6(n9685), 
           .MA5(n9684), .MA4(n9683), .MA3(n9682), .MA2(n9681), .MA1(n9680), 
           .MA0(n9679), .MB35(n9787), .MB34(n9786), .MB33(n9785), .MB32(n9784), 
           .MB31(n9783), .MB30(n9782), .MB29(n9781), .MB28(n9780), .MB27(n9779), 
           .MB26(n9778), .MB25(n9777), .MB24(n9776), .MB23(n9775), .MB22(n9774), 
           .MB21(n9773), .MB20(n9772), .MB19(n9771), .MB18(n9770), .MB17(n9769), 
           .MB16(n9768), .MB15(n9767), .MB14(n9766), .MB13(n9765), .MB12(n9764), 
           .MB11(n9763), .MB10(n9762), .MB9(n9761), .MB8(n9760), .MB7(n9759), 
           .MB6(n9758), .MB5(n9757), .MB4(n9756), .MB3(n9755), .MB2(n9754), 
           .MB1(n9753), .MB0(n9752), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n9969), 
           .R52(n9968), .R51(n9967), .R50(n9966), .R49(n9965), .R48(n9964), 
           .R47(n9963), .R46(n9962), .R45(n9961), .R44(n9960), .R43(n9959), 
           .R42(n9958), .R41(n9957), .R40(n9956), .R39(n9955), .R38(n9954), 
           .R37(n9953), .R36(n9952), .R35(n9951), .R34(n9950), .R33(n9949), 
           .R32(n9948), .R31(n9947), .R30(n9946), .R29(n9945), .R28(n9944), 
           .R27(n9943), .R26(n9942), .R25(n9941), .R24(n9940), .R23(n9939), 
           .R22(n9938), .R21(n9937), .R20(n9936), .R19(n9935), .R18(n9934), 
           .R17(a_inv_c_1), .R16(a_inv_c_0), .R15(n9626), .R14(n9627), 
           .R13(n9628), .R12(n9629), .R11(n9630), .R10(n9631), .R9(n9632), 
           .R8(n9633), .R7(n9634), .R6(n9635), .R5(n9636), .R4(n9637), 
           .R3(n9638), .R2(n9639), .R1(n9640), .R0(n9641), .SIGNEDR(n9970));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam lat_alu_3.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_3.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_3.REG_FLAG_CLK = "NONE";
    defparam lat_alu_3.REG_FLAG_CE = "CE0";
    defparam lat_alu_3.REG_FLAG_RST = "RST0";
    defparam lat_alu_3.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASK01 = "0x00000000000000";
    defparam lat_alu_3.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_3.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_3.CLK0_DIV = "ENABLED";
    defparam lat_alu_3.CLK1_DIV = "ENABLED";
    defparam lat_alu_3.CLK2_DIV = "ENABLED";
    defparam lat_alu_3.CLK3_DIV = "ENABLED";
    defparam lat_alu_3.MCPAT = "0x00000000000000";
    defparam lat_alu_3.MASKPAT = "0x00000000000000";
    defparam lat_alu_3.RNDPAT = "0x00000000000000";
    defparam lat_alu_3.GSR = "DISABLED";
    defparam lat_alu_3.RESETMODE = "SYNC";
    defparam lat_alu_3.MULT9_MODE = "DISABLED";
    defparam lat_alu_3.LEGACY = "DISABLED";
    MULT18X18D lat_mult_2 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68_adj_185), .B16(n68_adj_185), 
            .B15(n68_adj_185), .B14(n68_adj_185), .B13(n68_adj_185), .B12(n68_adj_185), 
            .B11(n68_adj_185), .B10(n68_adj_185), .B9(n68_adj_185), .B8(n68_adj_185), 
            .B7(n68_adj_185), .B6(n68_adj_185), .B5(n68_adj_185), .B4(n68_adj_185), 
            .B3(n68_adj_185), .B2(n68_adj_185), .B1(n68_adj_185), .B0(n68_adj_185), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n9878), .ROA16(n9877), 
            .ROA15(n9876), .ROA14(n9875), .ROA13(n9874), .ROA12(n9873), 
            .ROA11(n9872), .ROA10(n9871), .ROA9(n9870), .ROA8(n9869), 
            .ROA7(n9868), .ROA6(n9867), .ROA5(n9866), .ROA4(n9865), 
            .ROA3(n9864), .ROA2(n9863), .ROA1(n9862), .ROA0(n9861), 
            .ROB17(n9896), .ROB16(n9895), .ROB15(n9894), .ROB14(n9893), 
            .ROB13(n9892), .ROB12(n9891), .ROB11(n9890), .ROB10(n9889), 
            .ROB9(n9888), .ROB8(n9887), .ROB7(n9886), .ROB6(n9885), 
            .ROB5(n9884), .ROB4(n9883), .ROB3(n9882), .ROB2(n9881), 
            .ROB1(n9880), .ROB0(n9879), .P35(n9933), .P34(n9932), .P33(n9931), 
            .P32(n9930), .P31(n9929), .P30(n9928), .P29(n9927), .P28(n9926), 
            .P27(n9925), .P26(n9924), .P25(n9923), .P24(n9922), .P23(n9921), 
            .P22(n9920), .P21(n9919), .P20(n9918), .P19(n9917), .P18(n9916), 
            .P17(n9915), .P16(n9914), .P15(n9913), .P14(n9912), .P13(n9911), 
            .P12(n9910), .P11(n9909), .P10(n9908), .P9(n9907), .P8(n9906), 
            .P7(n9905), .P6(n9904), .P5(n9903), .P4(n9902), .P3(n9901), 
            .P2(n9900), .P1(n9899), .P0(n9898), .SIGNEDP(n9897));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam lat_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_2.REG_INPUTA_CE = "CE3";
    defparam lat_mult_2.REG_INPUTA_RST = "RST3";
    defparam lat_mult_2.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTB_CE = "CE0";
    defparam lat_mult_2.REG_INPUTB_RST = "RST0";
    defparam lat_mult_2.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTC_CE = "CE0";
    defparam lat_mult_2.REG_INPUTC_RST = "RST0";
    defparam lat_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_2.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_2.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_2.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_2.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_2.CLK0_DIV = "ENABLED";
    defparam lat_mult_2.CLK1_DIV = "ENABLED";
    defparam lat_mult_2.CLK2_DIV = "ENABLED";
    defparam lat_mult_2.CLK3_DIV = "ENABLED";
    defparam lat_mult_2.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_2.GSR = "DISABLED";
    defparam lat_mult_2.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_2.MULT_BYPASS = "DISABLED";
    defparam lat_mult_2.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_1 (.A17(n47), .A16(n48), .A15(n49), .A14(n50), 
            .A13(n51), .A12(n52), .A11(n53), .A10(n54), .A9(n55), 
            .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), .A3(n61), 
            .A2(n62), .A1(n63), .A0(n64), .B17(n68_adj_185), .B16(n68_adj_185), 
            .B15(n68_adj_185), .B14(n68_adj_185), .B13(n68_adj_185), .B12(n68_adj_185), 
            .B11(n68_adj_185), .B10(n68_adj_185), .B9(n68_adj_185), .B8(n68_adj_185), 
            .B7(n68_adj_185), .B6(n68_adj_185), .B5(n68_adj_185), .B4(n68_adj_185), 
            .B3(n68_adj_185), .B2(n68_adj_185), .B1(n68_adj_185), .B0(n68_adj_185), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n9805), .ROA16(n9804), 
            .ROA15(n9803), .ROA14(n9802), .ROA13(n9801), .ROA12(n9800), 
            .ROA11(n9799), .ROA10(n9798), .ROA9(n9797), .ROA8(n9796), 
            .ROA7(n9795), .ROA6(n9794), .ROA5(n9793), .ROA4(n9792), 
            .ROA3(n9791), .ROA2(n9790), .ROA1(n9789), .ROA0(n9788), 
            .ROB17(n9823), .ROB16(n9822), .ROB15(n9821), .ROB14(n9820), 
            .ROB13(n9819), .ROB12(n9818), .ROB11(n9817), .ROB10(n9816), 
            .ROB9(n9815), .ROB8(n9814), .ROB7(n9813), .ROB6(n9812), 
            .ROB5(n9811), .ROB4(n9810), .ROB3(n9809), .ROB2(n9808), 
            .ROB1(n9807), .ROB0(n9806), .P35(n9860), .P34(n9859), .P33(n9858), 
            .P32(n9857), .P31(n9856), .P30(n9855), .P29(n9854), .P28(n9853), 
            .P27(n9852), .P26(n9851), .P25(n9850), .P24(n9849), .P23(n9848), 
            .P22(n9847), .P21(n9846), .P20(n9845), .P19(n9844), .P18(n9843), 
            .P17(n9842), .P16(n9841), .P15(n9840), .P14(n9839), .P13(n9838), 
            .P12(n9837), .P11(n9836), .P10(n9835), .P9(n9834), .P8(n9833), 
            .P7(n9832), .P6(n9831), .P5(n9830), .P4(n9829), .P3(n9828), 
            .P2(n9827), .P1(n9826), .P0(n9825), .SIGNEDP(n9824));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam lat_mult_1.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_1.REG_INPUTA_CE = "CE3";
    defparam lat_mult_1.REG_INPUTA_RST = "RST3";
    defparam lat_mult_1.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTB_CE = "CE0";
    defparam lat_mult_1.REG_INPUTB_RST = "RST0";
    defparam lat_mult_1.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTC_CE = "CE0";
    defparam lat_mult_1.REG_INPUTC_RST = "RST0";
    defparam lat_mult_1.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_1.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_1.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_1.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_1.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_1.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_1.CLK0_DIV = "ENABLED";
    defparam lat_mult_1.CLK1_DIV = "ENABLED";
    defparam lat_mult_1.CLK2_DIV = "ENABLED";
    defparam lat_mult_1.CLK3_DIV = "ENABLED";
    defparam lat_mult_1.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_1.GSR = "DISABLED";
    defparam lat_mult_1.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_1.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_1.MULT_BYPASS = "DISABLED";
    defparam lat_mult_1.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_0 (.A17(n33), .A16(n33), .A15(n33), .A14(n33), 
            .A13(n33), .A12(n34), .A11(n35), .A10(n36), .A9(n37), 
            .A8(n38), .A7(n39), .A6(n40), .A5(n41), .A4(n42), .A3(n43), 
            .A2(n44), .A1(n45), .A0(n46), .B17(n68_adj_185), .B16(n68_adj_185), 
            .B15(n68_adj_185), .B14(n102_adj_170), .B13(n104_adj_184), 
            .B12(n106_adj_183), .B11(n108_adj_182), .B10(n110_adj_181), 
            .B9(n112_adj_180), .B8(n114_adj_179), .B7(n116_adj_178), .B6(n118_adj_177), 
            .B5(n120_adj_176), .B4(n122_adj_175), .B3(n124_adj_174), .B2(n126_adj_173), 
            .B1(n128_adj_172), .B0(n130_adj_171), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(clk_c), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(GND_net), 
            .RST3(reset_c), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .ROA17(n9732), .ROA16(n9731), .ROA15(n9730), .ROA14(n9729), 
            .ROA13(n9728), .ROA12(n9727), .ROA11(n9726), .ROA10(n9725), 
            .ROA9(n9724), .ROA8(n9723), .ROA7(n9722), .ROA6(n9721), 
            .ROA5(n9720), .ROA4(n9719), .ROA3(n9718), .ROA2(n9717), 
            .ROA1(n9716), .ROA0(n9715), .ROB17(n9750), .ROB16(n9749), 
            .ROB15(n9748), .ROB14(n9747), .ROB13(n9746), .ROB12(n9745), 
            .ROB11(n9744), .ROB10(n9743), .ROB9(n9742), .ROB8(n9741), 
            .ROB7(n9740), .ROB6(n9739), .ROB5(n9738), .ROB4(n9737), 
            .ROB3(n9736), .ROB2(n9735), .ROB1(n9734), .ROB0(n9733), 
            .P35(n9787), .P34(n9786), .P33(n9785), .P32(n9784), .P31(n9783), 
            .P30(n9782), .P29(n9781), .P28(n9780), .P27(n9779), .P26(n9778), 
            .P25(n9777), .P24(n9776), .P23(n9775), .P22(n9774), .P21(n9773), 
            .P20(n9772), .P19(n9771), .P18(n9770), .P17(n9769), .P16(n9768), 
            .P15(n9767), .P14(n9766), .P13(n9765), .P12(n9764), .P11(n9763), 
            .P10(n9762), .P9(n9761), .P8(n9760), .P7(n9759), .P6(n9758), 
            .P5(n9757), .P4(n9756), .P3(n9755), .P2(n9754), .P1(n9753), 
            .P0(n9752), .SIGNEDP(n9751));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam lat_mult_0.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_0.REG_INPUTA_CE = "CE3";
    defparam lat_mult_0.REG_INPUTA_RST = "RST3";
    defparam lat_mult_0.REG_INPUTB_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTB_CE = "CE0";
    defparam lat_mult_0.REG_INPUTB_RST = "RST0";
    defparam lat_mult_0.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTC_CE = "CE0";
    defparam lat_mult_0.REG_INPUTC_RST = "RST0";
    defparam lat_mult_0.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_0.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_0.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_0.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_0.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_0.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_0.CLK0_DIV = "ENABLED";
    defparam lat_mult_0.CLK1_DIV = "ENABLED";
    defparam lat_mult_0.CLK2_DIV = "ENABLED";
    defparam lat_mult_0.CLK3_DIV = "ENABLED";
    defparam lat_mult_0.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_0.GSR = "DISABLED";
    defparam lat_mult_0.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_0.MULT_BYPASS = "DISABLED";
    defparam lat_mult_0.RESETMODE = "ASYNC";
    LUT4 i393_2_lut (.A(prod_c[30]), .B(prod_c[29]), .Z(c_inv_c_14)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i393_2_lut.init = 16'h6666;
    MULT18X18D d_reg_15__I_0_mult_2 (.A17(n47), .A16(n48), .A15(n49), 
            .A14(n50), .A13(n51), .A12(n52), .A11(n53), .A10(n54), 
            .A9(n55), .A8(n56), .A7(n57), .A6(n58), .A5(n59), .A4(n60), 
            .A3(n61), .A2(n62), .A1(n63), .A0(n64), .B17(n68_adj_185), 
            .B16(n68_adj_185), .B15(n68_adj_185), .B14(n102_adj_170), 
            .B13(n104_adj_184), .B12(n106_adj_183), .B11(n108_adj_182), 
            .B10(n110_adj_181), .B9(n112_adj_180), .B8(n114_adj_179), 
            .B7(n116_adj_178), .B6(n118_adj_177), .B5(n120_adj_176), .B4(n122_adj_175), 
            .B3(n124_adj_174), .B2(n126_adj_173), .B1(n128_adj_172), .B0(n130_adj_171), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(clk_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(GND_net), .RST3(reset_c), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n9659), .ROA16(n9658), 
            .ROA15(n9657), .ROA14(n9656), .ROA13(n9655), .ROA12(n9654), 
            .ROA11(n9653), .ROA10(n9652), .ROA9(n9651), .ROA8(n9650), 
            .ROA7(n9649), .ROA6(n9648), .ROA5(n9647), .ROA4(n9646), 
            .ROA3(n9645), .ROA2(n9644), .ROA1(n9643), .ROA0(n9642), 
            .ROB17(n9677), .ROB16(n9676), .ROB15(n9675), .ROB14(n9674), 
            .ROB13(n9673), .ROB12(n9672), .ROB11(n9671), .ROB10(n9670), 
            .ROB9(n9669), .ROB8(n9668), .ROB7(n9667), .ROB6(n9666), 
            .ROB5(n9665), .ROB4(n9664), .ROB3(n9663), .ROB2(n9662), 
            .ROB1(n9661), .ROB0(n9660), .P35(n9714), .P34(n9713), .P33(n9712), 
            .P32(n9711), .P31(n9710), .P30(n9709), .P29(n9708), .P28(n9707), 
            .P27(n9706), .P26(n9705), .P25(n9704), .P24(n9703), .P23(n9702), 
            .P22(n9701), .P21(n9700), .P20(n9699), .P19(n9698), .P18(n9697), 
            .P17(n9696), .P16(n9695), .P15(n9694), .P14(n9693), .P13(n9692), 
            .P12(n9691), .P11(n9690), .P10(n9689), .P9(n9688), .P8(n9687), 
            .P7(n9686), .P6(n9685), .P5(n9684), .P4(n9683), .P3(n9682), 
            .P2(n9681), .P1(n9680), .P0(n9679), .SIGNEDP(n9678));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam d_reg_15__I_0_mult_2.REG_INPUTA_CE = "CE3";
    defparam d_reg_15__I_0_mult_2.REG_INPUTA_RST = "RST3";
    defparam d_reg_15__I_0_mult_2.REG_INPUTB_CLK = "NONE";
    defparam d_reg_15__I_0_mult_2.REG_INPUTB_CE = "CE0";
    defparam d_reg_15__I_0_mult_2.REG_INPUTB_RST = "RST0";
    defparam d_reg_15__I_0_mult_2.REG_INPUTC_CLK = "NONE";
    defparam d_reg_15__I_0_mult_2.REG_INPUTC_CE = "CE0";
    defparam d_reg_15__I_0_mult_2.REG_INPUTC_RST = "RST0";
    defparam d_reg_15__I_0_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam d_reg_15__I_0_mult_2.REG_PIPELINE_CE = "CE0";
    defparam d_reg_15__I_0_mult_2.REG_PIPELINE_RST = "RST0";
    defparam d_reg_15__I_0_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam d_reg_15__I_0_mult_2.REG_OUTPUT_CE = "CE0";
    defparam d_reg_15__I_0_mult_2.REG_OUTPUT_RST = "RST0";
    defparam d_reg_15__I_0_mult_2.CLK0_DIV = "ENABLED";
    defparam d_reg_15__I_0_mult_2.CLK1_DIV = "ENABLED";
    defparam d_reg_15__I_0_mult_2.CLK2_DIV = "ENABLED";
    defparam d_reg_15__I_0_mult_2.CLK3_DIV = "ENABLED";
    defparam d_reg_15__I_0_mult_2.HIGHSPEED_CLK = "NONE";
    defparam d_reg_15__I_0_mult_2.GSR = "DISABLED";
    defparam d_reg_15__I_0_mult_2.CAS_MATCH_REG = "FALSE";
    defparam d_reg_15__I_0_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam d_reg_15__I_0_mult_2.MULT_BYPASS = "DISABLED";
    defparam d_reg_15__I_0_mult_2.RESETMODE = "ASYNC";
    LUT4 i400_3_lut (.A(prod_c[31]), .B(prod_c[30]), .C(prod_c[29]), .Z(c_inv_c_15)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i400_3_lut.init = 16'h6a6a;
    LUT4 mux_294_i1_3_lut_rep_84 (.A(n68_adj_1394), .B(n68_adj_1426), .C(n1536), 
         .Z(n13020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_294_i1_3_lut_rep_84.init = 16'hcaca;
    LUT4 i1362_2_lut_4_lut (.A(n68_adj_1394), .B(n68_adj_1426), .C(n1536), 
         .D(det_zero), .Z(n42)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1362_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_295_i1_3_lut_rep_85 (.A(n68_adj_1330), .B(n68_adj_1362), .C(n1536), 
         .Z(n13021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_295_i1_3_lut_rep_85.init = 16'hcaca;
    LUT4 i1365_2_lut_4_lut (.A(n68_adj_1330), .B(n68_adj_1362), .C(n1536), 
         .D(det_zero), .Z(n41)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1365_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_296_i1_3_lut_rep_86 (.A(n68_adj_1268), .B(n68_adj_1299), .C(n1536), 
         .Z(n13022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_296_i1_3_lut_rep_86.init = 16'hcaca;
    LUT4 i1389_2_lut_4_lut (.A(n68_adj_1268), .B(n68_adj_1299), .C(n1536), 
         .D(det_zero), .Z(n40)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1389_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_304_i1_3_lut_rep_87 (.A(n68_adj_918), .B(n68_adj_886), .C(n1033), 
         .Z(n13023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_304_i1_3_lut_rep_87.init = 16'hcaca;
    LUT4 i1371_2_lut_4_lut (.A(n68_adj_918), .B(n68_adj_886), .C(n1033), 
         .D(det_zero), .Z(n38)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1371_2_lut_4_lut.init = 16'h0035;
    LUT4 i785_2_lut_4_lut (.A(n68_adj_918), .B(n68_adj_886), .C(n1033), 
         .D(n1067), .Z(n1503)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i785_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_303_i1_3_lut_rep_88 (.A(n68_adj_982), .B(n68_adj_950), .C(n1033), 
         .Z(n13024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_303_i1_3_lut_rep_88.init = 16'hcaca;
    LUT4 i369_1_lut (.A(prod_b[29]), .Z(b_inv_c_13)) /* synthesis lut_function=(!(A)) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i369_1_lut.init = 16'h5555;
    LUT4 i1374_2_lut_4_lut (.A(n68_adj_982), .B(n68_adj_950), .C(n1033), 
         .D(det_zero), .Z(n37)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1374_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_302_i1_3_lut_rep_89 (.A(n68_adj_1046), .B(n68_adj_1014), .C(n1033), 
         .Z(n13025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_302_i1_3_lut_rep_89.init = 16'hcaca;
    LUT4 i1377_2_lut_4_lut (.A(n68_adj_1046), .B(n68_adj_1014), .C(n1033), 
         .D(det_zero), .Z(n36)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1377_2_lut_4_lut.init = 16'h0035;
    FD1S3AX c_reg_i14 (.D(c_c_14), .CK(clk_c), .Q(c_reg[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i14.GSR = "ENABLED";
    LUT4 mux_301_i1_3_lut_rep_90 (.A(n68_adj_1110), .B(n68_adj_1078), .C(n1033), 
         .Z(n13026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_301_i1_3_lut_rep_90.init = 16'hcaca;
    CCU2C _add_1_609_add_4_23 (.A0(n101_adj_293), .B0(n3077), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_292), .B1(n3077), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11864), .COUT(n11865), .S0(n98_adj_196), 
          .S1(n95_adj_195));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_21 (.A0(n107_adj_295), .B0(n3077), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_294), .B1(n3077), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11863), .COUT(n11864), .S0(n104_adj_198), 
          .S1(n101_adj_197));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_21.INJECT1_1 = "NO";
    FD1S3AX c_reg_i13 (.D(c_c_13), .CK(clk_c), .Q(c_reg[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i13.GSR = "ENABLED";
    CCU2C _add_1_609_add_4_19 (.A0(n113_adj_297), .B0(n3077), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_296), .B1(n3077), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11862), .COUT(n11863), .S0(n110_adj_200), 
          .S1(n107_adj_199));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_17 (.A0(n119_adj_299), .B0(n3077), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_298), .B1(n3077), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11861), .COUT(n11862), .S0(n116_adj_202), 
          .S1(n113_adj_201));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_17.INJECT1_1 = "NO";
    FD1S3AX c_reg_i12 (.D(c_c_12), .CK(clk_c), .Q(c_reg[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i12.GSR = "ENABLED";
    CCU2C _add_1_609_add_4_15 (.A0(n125_adj_301), .B0(n3077), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_300), .B1(n3077), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11860), .COUT(n11861), .S0(n122_adj_204), 
          .S1(n119_adj_203));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_13 (.A0(n131_adj_303), .B0(n3077), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_302), .B1(n3077), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11859), .COUT(n11860), .S0(n128_adj_206), 
          .S1(n125_adj_205));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_11 (.A0(n137_adj_305), .B0(n3077), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_304), .B1(n3077), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11858), .COUT(n11859), .S0(n134_adj_208), 
          .S1(n131_adj_207));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_9 (.A0(n143_adj_307), .B0(n3077), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_306), .B1(n3077), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11857), .COUT(n11858), .S0(n140_adj_210), 
          .S1(n137_adj_209));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_9.INJECT1_1 = "NO";
    FD1S3AX c_reg_i11 (.D(c_c_11), .CK(clk_c), .Q(c_reg[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i11.GSR = "ENABLED";
    CCU2C _add_1_609_add_4_7 (.A0(n149_adj_309), .B0(n3077), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_308), .B1(n3077), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11856), .COUT(n11857), .S0(n146_adj_212), 
          .S1(n143_adj_211));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_5 (.A0(n155_adj_311), .B0(n3077), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_310), .B1(n3077), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11855), .COUT(n11856), .S0(n152_adj_214), 
          .S1(n149_adj_213));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_609_add_4_3 (.A0(n161_adj_313), .B0(n3077), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_312), .B1(n3077), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11854), .COUT(n11855), .S0(n158_adj_216), 
          .S1(n155_adj_215));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_609_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_3.INJECT1_1 = "NO";
    FD1S3AX c_reg_i10 (.D(c_c_10), .CK(clk_c), .Q(c_reg[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i10.GSR = "ENABLED";
    CCU2C _add_1_609_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n3077), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11854), .S1(n161_adj_217));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_609_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_609_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_609_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_609_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_33 (.A0(n1067), .B0(n13017), .C0(n71_adj_1907), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11853), .S0(n68_adj_218));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_435_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_435_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_31 (.A0(n77_adj_1909), .B0(n13017), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1908), .B1(n13017), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11852), .COUT(n11853), .S0(n74_adj_220), 
          .S1(n71_adj_219));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_29 (.A0(n83_adj_1911), .B0(n13017), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1910), .B1(n13017), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11851), .COUT(n11852), .S0(n80_adj_222), 
          .S1(n77_adj_221));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_29.INJECT1_1 = "NO";
    FD1S3AX c_reg_i9 (.D(c_c_9), .CK(clk_c), .Q(c_reg[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i9.GSR = "ENABLED";
    CCU2C _add_1_435_add_4_27 (.A0(n89_adj_1913), .B0(n13017), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1912), .B1(n13017), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11850), .COUT(n11851), .S0(n86_adj_224), 
          .S1(n83_adj_223));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_25 (.A0(n95_adj_1915), .B0(n13017), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1914), .B1(n13017), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11849), .COUT(n11850), .S0(n92_adj_226), 
          .S1(n89_adj_225));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_23 (.A0(n101_adj_1917), .B0(n13017), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1916), .B1(n13017), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11848), .COUT(n11849), .S0(n98_adj_228), 
          .S1(n95_adj_227));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_23.INJECT1_1 = "NO";
    FD1S3AX c_reg_i8 (.D(c_c_8), .CK(clk_c), .Q(c_reg[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i8.GSR = "ENABLED";
    CCU2C _add_1_435_add_4_21 (.A0(n107_adj_1919), .B0(n13017), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1918), .B1(n13017), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11847), .COUT(n11848), .S0(n104_adj_230), 
          .S1(n101_adj_229));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_19 (.A0(n113_adj_1921), .B0(n13017), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1920), .B1(n13017), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11846), .COUT(n11847), .S0(n110_adj_232), 
          .S1(n107_adj_231));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_17 (.A0(n119_adj_1923), .B0(n13017), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1922), .B1(n13017), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11845), .COUT(n11846), .S0(n116_adj_234), 
          .S1(n113_adj_233));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_15 (.A0(n125_adj_1925), .B0(n13017), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1924), .B1(n13017), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11844), .COUT(n11845), .S0(n122_adj_236), 
          .S1(n119_adj_235));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_15.INJECT1_1 = "NO";
    FD1S3AX c_reg_i7 (.D(c_c_7), .CK(clk_c), .Q(c_reg[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i7.GSR = "ENABLED";
    CCU2C _add_1_435_add_4_13 (.A0(n131_adj_1927), .B0(n13017), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1926), .B1(n13017), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11843), .COUT(n11844), .S0(n128_adj_238), 
          .S1(n125_adj_237));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_11 (.A0(n137_adj_1929), .B0(n13017), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1928), .B1(n13017), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11842), .COUT(n11843), .S0(n134_adj_240), 
          .S1(n131_adj_239));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_9 (.A0(n143_adj_1931), .B0(n13017), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1930), .B1(n13017), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11841), .COUT(n11842), .S0(n140_adj_242), 
          .S1(n137_adj_241));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_9.INJECT1_1 = "NO";
    FD1S3AX det_q4_28_res1_i28 (.D(det_q4_28_31__N_1[28]), .CK(clk_c), .Q(det_q4_28[28]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i28.GSR = "ENABLED";
    CCU2C _add_1_435_add_4_7 (.A0(n149_adj_1933), .B0(n13017), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1932), .B1(n13017), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11840), .COUT(n11841), .S0(n146_adj_244), 
          .S1(n143_adj_243));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_7.INJECT1_1 = "NO";
    FD1S3AX det_q4_28_res1_i29 (.D(det_q4_28_31__N_1[29]), .CK(clk_c), .Q(det_q4_28[29]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i29.GSR = "ENABLED";
    FD1S3AX c_reg_i6 (.D(c_c_6), .CK(clk_c), .Q(c_reg[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i6.GSR = "ENABLED";
    CCU2C _add_1_435_add_4_5 (.A0(n155_adj_1935), .B0(n13017), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1934), .B1(n13017), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11839), .COUT(n11840), .S0(n152_adj_246), 
          .S1(n149_adj_245));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_5.INJECT1_1 = "NO";
    FD1S3AX c_reg_i5 (.D(c_c_5), .CK(clk_c), .Q(c_reg[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i5.GSR = "ENABLED";
    CCU2C _add_1_435_add_4_3 (.A0(n161_adj_1937), .B0(n13017), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1936), .B1(n13017), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11838), .COUT(n11839), .S0(n158_adj_248), 
          .S1(n155_adj_247));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_435_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_435_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13017), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11838), .S1(n161_adj_249));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_435_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_435_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_435_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_435_add_4_1.INJECT1_1 = "NO";
    FD1S3AX det_q4_28_res1_i21 (.D(det_q4_28_31__N_1[21]), .CK(clk_c), .Q(det_q4_28[21]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i21.GSR = "ENABLED";
    CCU2C _add_1_606_add_4_33 (.A0(n74_adj_315), .B0(n2273), .C0(n71_adj_187), 
          .D0(n3112), .A1(n71_adj_314), .B1(n2273), .C1(n68_adj_186), 
          .D1(n3111), .CIN(n11836), .S0(n71_adj_251), .S1(n68_adj_250));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_33.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_33.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_33.INJECT1_1 = "NO";
    FD1S3AX det_q4_28_res1_i22 (.D(det_q4_28_31__N_1[22]), .CK(clk_c), .Q(det_q4_28[22]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i22.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i31 (.D(det_q4_28_31__N_1[31]), .CK(clk_c), .Q(det_q4_28[31]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i31.GSR = "ENABLED";
    FD1S3AX c_reg_i4 (.D(c_c_4), .CK(clk_c), .Q(c_reg[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i4.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i30 (.D(det_q4_28_31__N_1[30]), .CK(clk_c), .Q(det_q4_28[30]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i30.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i25 (.D(det_q4_28_31__N_1[25]), .CK(clk_c), .Q(det_q4_28[25]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i25.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i26 (.D(det_q4_28_31__N_1[26]), .CK(clk_c), .Q(det_q4_28[26]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i26.GSR = "ENABLED";
    FD1S3AX c_reg_i3 (.D(c_c_3), .CK(clk_c), .Q(c_reg[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i3.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i27 (.D(det_q4_28_31__N_1[27]), .CK(clk_c), .Q(det_q4_28[27]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i27.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i14 (.D(det_q4_28_31__N_1[14]), .CK(clk_c), .Q(det_q4_28[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i14.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i15 (.D(det_q4_28_31__N_1[15]), .CK(clk_c), .Q(det_q4_28[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i15.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i24 (.D(det_q4_28_31__N_1[24]), .CK(clk_c), .Q(det_q4_28[24]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i24.GSR = "ENABLED";
    FD1S3AX c_reg_i2 (.D(c_c_2), .CK(clk_c), .Q(c_reg[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i2.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i23 (.D(det_q4_28_31__N_1[23]), .CK(clk_c), .Q(det_q4_28[23]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i23.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i18 (.D(det_q4_28_31__N_1[18]), .CK(clk_c), .Q(det_q4_28[18]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i18.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i19 (.D(det_q4_28_31__N_1[19]), .CK(clk_c), .Q(det_q4_28[19]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i19.GSR = "ENABLED";
    FD1S3AX c_reg_i1 (.D(c_c_1), .CK(clk_c), .Q(c_reg[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i1.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i20 (.D(det_q4_28_31__N_1[20]), .CK(clk_c), .Q(det_q4_28[20]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i20.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i9 (.D(det_q4_28_31__N_1[9]), .CK(clk_c), .Q(det_q4_28[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i9.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i10 (.D(det_q4_28_31__N_1[10]), .CK(clk_c), .Q(det_q4_28[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i10.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i17 (.D(det_q4_28_31__N_1[17]), .CK(clk_c), .Q(det_q4_28[17]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i17.GSR = "ENABLED";
    FD1S3AX b_reg_i15 (.D(b_c_15), .CK(clk_c), .Q(b_reg[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i15.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i16 (.D(det_q4_28_31__N_1[16]), .CK(clk_c), .Q(det_q4_28[16]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i16.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i11 (.D(det_q4_28_31__N_1[11]), .CK(clk_c), .Q(det_q4_28[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i11.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i12 (.D(det_q4_28_31__N_1[12]), .CK(clk_c), .Q(det_q4_28[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i12.GSR = "ENABLED";
    FD1S3AX b_reg_i14 (.D(b_c_14), .CK(clk_c), .Q(b_reg[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i14.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i13 (.D(det_q4_28_31__N_1[13]), .CK(clk_c), .Q(det_q4_28[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i13.GSR = "ENABLED";
    FD1S3AX b_reg_i13 (.D(b_c_13), .CK(clk_c), .Q(b_reg[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i13.GSR = "ENABLED";
    IB a_pad_6 (.I(a[6]), .O(a_c_6));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_5 (.I(a[5]), .O(a_c_5));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB d_pad_14 (.I(d[14]), .O(d_c_14));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    FD1S3AX b_reg_i12 (.D(b_c_12), .CK(clk_c), .Q(b_reg[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i12.GSR = "ENABLED";
    IB d_pad_15 (.I(d[15]), .O(d_c_15));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB a_pad_4 (.I(a[4]), .O(a_c_4));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_3 (.I(a[3]), .O(a_c_3));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    FD1S3AX det_q4_28_res1_i3 (.D(det_q4_28_31__N_1[3]), .CK(clk_c), .Q(det_q4_28[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i3.GSR = "ENABLED";
    IB c_pad_4 (.I(c[4]), .O(c_c_4));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    LUT4 i371_2_lut (.A(prod_b[30]), .B(prod_b[29]), .Z(b_inv_c_14)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i371_2_lut.init = 16'h6666;
    LUT4 i378_3_lut (.A(prod_b[31]), .B(prod_b[30]), .C(prod_b[29]), .Z(b_inv_c_15)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i378_3_lut.init = 16'h6a6a;
    FD1S3AX b_reg_i11 (.D(b_c_11), .CK(clk_c), .Q(b_reg[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i11.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i2 (.D(det_q4_28_31__N_1[2]), .CK(clk_c), .Q(det_q4_28[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i2.GSR = "ENABLED";
    FD1S3AX b_reg_i10 (.D(b_c_10), .CK(clk_c), .Q(b_reg[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i10.GSR = "ENABLED";
    LUT4 i347_1_lut (.A(prod_a[29]), .Z(a_inv_c_13)) /* synthesis lut_function=(!(A)) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i347_1_lut.init = 16'h5555;
    LUT4 i349_2_lut (.A(prod_a[30]), .B(prod_a[29]), .Z(a_inv_c_14)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i349_2_lut.init = 16'h6666;
    FD1S3AX b_reg_i9 (.D(b_c_9), .CK(clk_c), .Q(b_reg[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i9.GSR = "ENABLED";
    LUT4 i807_2_lut_4_lut (.A(n68_adj_377), .B(n68_adj_345), .C(n2273), 
         .D(n1067), .Z(n3044)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i807_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_314_i1_3_lut_rep_69 (.A(n68_adj_472), .B(n68_adj_440), .C(n2273), 
         .Z(n13005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_314_i1_3_lut_rep_69.init = 16'hcaca;
    LUT4 i1443_2_lut_4_lut (.A(n68_adj_472), .B(n68_adj_440), .C(n2273), 
         .D(det_zero), .Z(n60)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1443_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_313_i1_3_lut_rep_70 (.A(n68_adj_536), .B(n68_adj_504), .C(n2273), 
         .Z(n13006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_313_i1_3_lut_rep_70.init = 16'hcaca;
    FD1S3AX b_reg_i8 (.D(b_c_8), .CK(clk_c), .Q(b_reg[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i8.GSR = "ENABLED";
    LUT4 i1434_2_lut_4_lut (.A(n68_adj_536), .B(n68_adj_504), .C(n2273), 
         .D(det_zero), .Z(n59)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1434_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_312_i1_3_lut_rep_71 (.A(n68_adj_600), .B(n68_adj_568), .C(n2273), 
         .Z(n13007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_312_i1_3_lut_rep_71.init = 16'hcaca;
    LUT4 i1437_2_lut_4_lut (.A(n68_adj_600), .B(n68_adj_568), .C(n2273), 
         .D(det_zero), .Z(n58)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1437_2_lut_4_lut.init = 16'h0035;
    FD1S3AX b_reg_i7 (.D(b_c_7), .CK(clk_c), .Q(b_reg[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i7.GSR = "ENABLED";
    LUT4 mux_311_i1_3_lut_rep_72 (.A(n68_adj_1681), .B(n68_adj_1649), .C(n2273), 
         .Z(n13008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_311_i1_3_lut_rep_72.init = 16'hcaca;
    LUT4 i1440_2_lut_4_lut (.A(n68_adj_1681), .B(n68_adj_1649), .C(n2273), 
         .D(det_zero), .Z(n57)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1440_2_lut_4_lut.init = 16'h0035;
    FD1S3AX b_reg_i6 (.D(b_c_6), .CK(clk_c), .Q(b_reg[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i6.GSR = "ENABLED";
    LUT4 mux_310_i1_3_lut_rep_73 (.A(n68_adj_1842), .B(n68_adj_1778), .C(n2273), 
         .Z(n13009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_310_i1_3_lut_rep_73.init = 16'hcaca;
    FD1S3AX b_reg_i5 (.D(b_c_5), .CK(clk_c), .Q(b_reg[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i5.GSR = "ENABLED";
    IB a_pad_1 (.I(a[1]), .O(a_c_1));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    LUT4 i1401_2_lut_4_lut (.A(n68_adj_1842), .B(n68_adj_1778), .C(n2273), 
         .D(det_zero), .Z(n56)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1401_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_309_i1_3_lut_rep_74 (.A(n68_adj_1970), .B(n68_adj_1938), .C(n2273), 
         .Z(n13010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_309_i1_3_lut_rep_74.init = 16'hcaca;
    LUT4 i1404_2_lut_4_lut (.A(n68_adj_1970), .B(n68_adj_1938), .C(n2273), 
         .D(det_zero), .Z(n55)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1404_2_lut_4_lut.init = 16'h0035;
    FD1S3AX b_reg_i4 (.D(b_c_4), .CK(clk_c), .Q(b_reg[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i4.GSR = "ENABLED";
    LUT4 mux_308_i1_3_lut_rep_75 (.A(n68_adj_2034), .B(n68_adj_2002), .C(n2273), 
         .Z(n13011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_308_i1_3_lut_rep_75.init = 16'hcaca;
    LUT4 i1431_2_lut_4_lut (.A(n68_adj_2034), .B(n68_adj_2002), .C(n2273), 
         .D(det_zero), .Z(n54)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1431_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_307_i1_3_lut_rep_76 (.A(n68_adj_664), .B(n68_adj_632), .C(n2273), 
         .Z(n13012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_307_i1_3_lut_rep_76.init = 16'hcaca;
    FD1S3AX b_reg_i3 (.D(b_c_3), .CK(clk_c), .Q(b_reg[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i3.GSR = "ENABLED";
    LUT4 i1428_2_lut_4_lut (.A(n68_adj_664), .B(n68_adj_632), .C(n2273), 
         .D(det_zero), .Z(n53)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1428_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_306_i1_3_lut_rep_77 (.A(n68_adj_728), .B(n68_adj_696), .C(n2273), 
         .Z(n13013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_306_i1_3_lut_rep_77.init = 16'hcaca;
    FD1S3AX b_reg_i2 (.D(b_c_2), .CK(clk_c), .Q(b_reg[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i2.GSR = "ENABLED";
    LUT4 i1413_2_lut_4_lut (.A(n68_adj_728), .B(n68_adj_696), .C(n2273), 
         .D(det_zero), .Z(n52)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1413_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_305_i1_3_lut_rep_78 (.A(n68_adj_792), .B(n68_adj_760), .C(n2273), 
         .Z(n13014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_305_i1_3_lut_rep_78.init = 16'hcaca;
    LUT4 i1416_2_lut_4_lut (.A(n68_adj_792), .B(n68_adj_760), .C(n2273), 
         .D(det_zero), .Z(n51)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1416_2_lut_4_lut.init = 16'h0035;
    FD1S3AX b_reg_i1 (.D(b_c_1), .CK(clk_c), .Q(b_reg[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i1.GSR = "ENABLED";
    LUT4 mux_297_i1_3_lut_rep_79 (.A(n68_adj_1143), .B(n68_adj_1175), .C(n2139), 
         .Z(n13015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_297_i1_3_lut_rep_79.init = 16'hcaca;
    LUT4 i1380_2_lut_4_lut (.A(n68_adj_1143), .B(n68_adj_1175), .C(n2139), 
         .D(det_zero), .Z(n49)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1380_2_lut_4_lut.init = 16'h0035;
    FD1S3AX b_reg_i0 (.D(b_c_0), .CK(clk_c), .Q(b_reg[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam b_reg_i0.GSR = "ENABLED";
    IB b_pad_15 (.I(b[15]), .O(b_c_15));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    LUT4 i732_2_lut_4_lut (.A(n68_adj_1143), .B(n68_adj_1175), .C(n2139), 
         .D(n1067), .Z(n2240)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i732_2_lut_4_lut.init = 16'h3500;
    OB d_inv_pad_2 (.I(d_inv_c_2), .O(d_inv[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_1 (.I(d_inv_c_1), .O(d_inv[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_0 (.I(d_inv_c_0), .O(d_inv[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB error_pad (.I(error_c), .O(error));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(19[26:31])
    OB d_inv_pad_12 (.I(d_inv_c_12), .O(d_inv[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    IB d_pad_6 (.I(d[6]), .O(d_c_6));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_5 (.I(d[5]), .O(d_c_5));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_2 (.I(d[2]), .O(d_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_1 (.I(d[1]), .O(d_c_1));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_0 (.I(d[0]), .O(d_c_0));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_11 (.I(d[11]), .O(d_c_11));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_10 (.I(d[10]), .O(d_c_10));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_3 (.I(d[3]), .O(d_c_3));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_4 (.I(d[4]), .O(d_c_4));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_9 (.I(d[9]), .O(d_c_9));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_8 (.I(d[8]), .O(d_c_8));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_7 (.I(d[7]), .O(d_c_7));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB clk_pad (.I(clk), .O(clk_c));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[20:23])
    IB reset_pad (.I(reset), .O(reset_c));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[25:30])
    IB a_pad_9 (.I(a[9]), .O(a_c_9));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_10 (.I(a[10]), .O(a_c_10));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_15 (.I(a[15]), .O(a_c_15));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_14 (.I(a[14]), .O(a_c_14));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_13 (.I(a[13]), .O(a_c_13));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB c_pad_11 (.I(c[11]), .O(c_c_11));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_10 (.I(c[10]), .O(c_c_10));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_1 (.I(c[1]), .O(c_c_1));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_2 (.I(c[2]), .O(c_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_7 (.I(c[7]), .O(c_c_7));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_6 (.I(c[6]), .O(c_c_6));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_5 (.I(c[5]), .O(c_c_5));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB b_pad_2 (.I(b[2]), .O(b_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB b_pad_1 (.I(b[1]), .O(b_c_1));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB c_pad_8 (.I(c[8]), .O(c_c_8));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_9 (.I(c[9]), .O(c_c_9));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_14 (.I(c[14]), .O(c_c_14));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_13 (.I(c[13]), .O(c_c_13));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_12 (.I(c[12]), .O(c_c_12));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB b_pad_9 (.I(b[9]), .O(b_c_9));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB b_pad_8 (.I(b[8]), .O(b_c_8));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB c_pad_15 (.I(c[15]), .O(c_c_15));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB b_pad_0 (.I(b[0]), .O(b_c_0));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB b_pad_5 (.I(b[5]), .O(b_c_5));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB b_pad_4 (.I(b[4]), .O(b_c_4));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    FD1S3AX det_q4_28_res1_i7 (.D(det_q4_28_31__N_1[7]), .CK(clk_c), .Q(det_q4_28[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i7.GSR = "ENABLED";
    IB b_pad_3 (.I(b[3]), .O(b_c_3));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB a_pad_2 (.I(a[2]), .O(a_c_2));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB a_pad_0 (.I(a[0]), .O(a_c_0));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    IB b_pad_6 (.I(b[6]), .O(b_c_6));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    OB a_inv_pad_15 (.I(a_inv_c_15), .O(a_inv[15]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[26:31])
    IB b_pad_7 (.I(b[7]), .O(b_c_7));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB b_pad_12 (.I(b[12]), .O(b_c_12));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    IB b_pad_11 (.I(b[11]), .O(b_c_11));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    GSR GSR_INST (.GSR(n11172));
    IB b_pad_10 (.I(b[10]), .O(b_c_10));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    OB d_inv_pad_13 (.I(d_inv_c_13), .O(d_inv[13]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    IB b_pad_14 (.I(b[14]), .O(b_c_14));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[29:30])
    FD1S3AX det_q4_28_res1_i6 (.D(det_q4_28_31__N_1[6]), .CK(clk_c), .Q(det_q4_28[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i6.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i5 (.D(det_q4_28_31__N_1[5]), .CK(clk_c), .Q(det_q4_28[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i5.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i4 (.D(det_q4_28_31__N_1[4]), .CK(clk_c), .Q(det_q4_28[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i4.GSR = "ENABLED";
    FD1S3AX det_q4_28_res1_i1 (.D(det_q4_28_31__N_1[1]), .CK(clk_c), .Q(det_q4_28[1]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam det_q4_28_res1_i1.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i2 (.D(d_c_1), .CK(clk_c), .Q(n128_adj_172));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i2.GSR = "ENABLED";
    LUT4 mux_290_i1_3_lut_rep_80 (.A(n68_adj_218), .B(n68_adj_1810), .C(n1536), 
         .Z(n13016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_290_i1_3_lut_rep_80.init = 16'hcaca;
    LUT4 i1407_2_lut_4_lut (.A(n68_adj_218), .B(n68_adj_1810), .C(n1536), 
         .D(det_zero), .Z(n46)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1407_2_lut_4_lut.init = 16'h0035;
    LUT4 i781_2_lut_4_lut (.A(n68_adj_218), .B(n68_adj_1810), .C(n1536), 
         .D(n1067), .Z(n2039)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i781_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_291_i1_3_lut_rep_81 (.A(n68_adj_1906), .B(n68_adj_1617), .C(n1536), 
         .Z(n13017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_291_i1_3_lut_rep_81.init = 16'hcaca;
    LUT4 i1392_2_lut_4_lut (.A(n68_adj_1906), .B(n68_adj_1617), .C(n1536), 
         .D(det_zero), .Z(n45)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1392_2_lut_4_lut.init = 16'h0035;
    IB d_pad_12 (.I(d[12]), .O(d_c_12));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB d_pad_13 (.I(d[13]), .O(d_c_13));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[35:36])
    IB c_pad_0 (.I(c[0]), .O(c_c_0));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    IB c_pad_3 (.I(c[3]), .O(c_c_3));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[32:33])
    OB d_inv_pad_3 (.I(d_inv_c_3), .O(d_inv[3]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_4 (.I(d_inv_c_4), .O(d_inv[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_5 (.I(d_inv_c_5), .O(d_inv[5]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_6 (.I(d_inv_c_6), .O(d_inv[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_7 (.I(d_inv_c_7), .O(d_inv[7]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_8 (.I(d_inv_c_8), .O(d_inv[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_9 (.I(d_inv_c_9), .O(d_inv[9]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_10 (.I(d_inv_c_10), .O(d_inv[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    OB d_inv_pad_11 (.I(d_inv_c_11), .O(d_inv[11]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(18[47:52])
    IB a_pad_12 (.I(a[12]), .O(a_c_12));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(17[26:27])
    LUT4 mux_292_i1_3_lut_rep_82 (.A(n68_adj_1522), .B(n68_adj_2098), .C(n1536), 
         .Z(n13018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_292_i1_3_lut_rep_82.init = 16'hcaca;
    LUT4 i1395_2_lut_4_lut (.A(n68_adj_1522), .B(n68_adj_2098), .C(n1536), 
         .D(det_zero), .Z(n44)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1395_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_293_i1_3_lut_rep_83 (.A(n68_adj_1458), .B(n68_adj_1490), .C(n1536), 
         .Z(n13019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_293_i1_3_lut_rep_83.init = 16'hcaca;
    LUT4 i1398_2_lut_4_lut (.A(n68_adj_1458), .B(n68_adj_1490), .C(n1536), 
         .D(det_zero), .Z(n43)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1398_2_lut_4_lut.init = 16'h0035;
    LUT4 det_zero_I_0_2_lut (.A(det_zero), .B(error_recip), .Z(error_c)) /* synthesis lut_function=(A+(B)) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(70[20:42])
    defparam det_zero_I_0_2_lut.init = 16'heeee;
    LUT4 i356_3_lut (.A(prod_a[31]), .B(prod_a[30]), .C(prod_a[29]), .Z(a_inv_c_15)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i356_3_lut.init = 16'h6a6a;
    LUT4 i724_1_lut (.A(reset_c), .Z(n11172)) /* synthesis lut_function=(!(A)) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[25:30])
    defparam i724_1_lut.init = 16'h5555;
    LUT4 i325_1_lut (.A(prod_d[29]), .Z(d_inv_c_13)) /* synthesis lut_function=(!(A)) */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(99[19:38])
    defparam i325_1_lut.init = 16'h5555;
    LUT4 i1244_2_lut (.A(det_q4_28[1]), .B(det_q4_28[0]), .Z(n161_adj_791)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1244_2_lut.init = 16'h6666;
    LUT4 i1248_2_lut (.A(n1098), .B(det_q4_28[0]), .Z(n161_adj_1174)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1248_2_lut.init = 16'h6666;
    CCU2C _add_1_606_add_4_31 (.A0(n80_adj_317), .B0(n2273), .C0(n77_adj_189), 
          .D0(n3114), .A1(n77_adj_316), .B1(n2273), .C1(n74_adj_188), 
          .D1(n3113), .CIN(n11835), .COUT(n11836), .S0(n77_adj_253), 
          .S1(n74_adj_252));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_29 (.A0(n86_adj_319), .B0(n2273), .C0(n83_adj_191), 
          .D0(n3116), .A1(n83_adj_318), .B1(n2273), .C1(n80_adj_190), 
          .D1(n3115), .CIN(n11834), .COUT(n11835), .S0(n83_adj_255), 
          .S1(n80_adj_254));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_27 (.A0(n92_adj_321), .B0(n2273), .C0(n89_adj_193), 
          .D0(n3118), .A1(n89_adj_320), .B1(n2273), .C1(n86_adj_192), 
          .D1(n3117), .CIN(n11833), .COUT(n11834), .S0(n89_adj_257), 
          .S1(n86_adj_256));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_25 (.A0(n98_adj_323), .B0(n2273), .C0(n95_adj_195), 
          .D0(n3120), .A1(n95_adj_322), .B1(n2273), .C1(n92_adj_194), 
          .D1(n3119), .CIN(n11832), .COUT(n11833), .S0(n95_adj_259), 
          .S1(n92_adj_258));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_23 (.A0(n104_adj_325), .B0(n2273), .C0(n101_adj_197), 
          .D0(n3122), .A1(n101_adj_324), .B1(n2273), .C1(n98_adj_196), 
          .D1(n3121), .CIN(n11831), .COUT(n11832), .S0(n101_adj_261), 
          .S1(n98_adj_260));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_21 (.A0(n110_adj_327), .B0(n2273), .C0(n107_adj_199), 
          .D0(n3124), .A1(n107_adj_326), .B1(n2273), .C1(n104_adj_198), 
          .D1(n3123), .CIN(n11830), .COUT(n11831), .S0(n107_adj_263), 
          .S1(n104_adj_262));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_19 (.A0(n116_adj_329), .B0(n2273), .C0(n113_adj_201), 
          .D0(n3126), .A1(n113_adj_328), .B1(n2273), .C1(n110_adj_200), 
          .D1(n3125), .CIN(n11829), .COUT(n11830), .S0(n113_adj_265), 
          .S1(n110_adj_264));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_17 (.A0(n122_adj_331), .B0(n2273), .C0(n119_adj_203), 
          .D0(n3128), .A1(n119_adj_330), .B1(n2273), .C1(n116_adj_202), 
          .D1(n3127), .CIN(n11828), .COUT(n11829), .S0(n119_adj_267), 
          .S1(n116_adj_266));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_15 (.A0(n128_adj_333), .B0(n2273), .C0(n125_adj_205), 
          .D0(n3130), .A1(n125_adj_332), .B1(n2273), .C1(n122_adj_204), 
          .D1(n3129), .CIN(n11827), .COUT(n11828), .S0(n125_adj_269), 
          .S1(n122_adj_268));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_13 (.A0(n134_adj_335), .B0(n2273), .C0(n131_adj_207), 
          .D0(n3132), .A1(n131_adj_334), .B1(n2273), .C1(n128_adj_206), 
          .D1(n3131), .CIN(n11826), .COUT(n11827), .S0(n131_adj_271), 
          .S1(n128_adj_270));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_11 (.A0(n140_adj_337), .B0(n2273), .C0(n137_adj_209), 
          .D0(n3134), .A1(n137_adj_336), .B1(n2273), .C1(n134_adj_208), 
          .D1(n3133), .CIN(n11825), .COUT(n11826), .S0(n137_adj_273), 
          .S1(n134_adj_272));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_9 (.A0(n146_adj_339), .B0(n2273), .C0(n143_adj_211), 
          .D0(n3136), .A1(n143_adj_338), .B1(n2273), .C1(n140_adj_210), 
          .D1(n3135), .CIN(n11824), .COUT(n11825), .S0(n143_adj_275), 
          .S1(n140_adj_274));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_7 (.A0(n152_adj_341), .B0(n2273), .C0(n149_adj_213), 
          .D0(n3138), .A1(n149_adj_340), .B1(n2273), .C1(n146_adj_212), 
          .D1(n3137), .CIN(n11823), .COUT(n11824), .S0(n149_adj_277), 
          .S1(n146_adj_276));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_5 (.A0(n158_adj_343), .B0(n2273), .C0(n155_adj_215), 
          .D0(n3140), .A1(n155_adj_342), .B1(n2273), .C1(n152_adj_214), 
          .D1(n3139), .CIN(n11822), .COUT(n11823), .S0(n155_adj_279), 
          .S1(n152_adj_278));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_606_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_3 (.A0(det_q4_28[0]), .B0(n2273), .C0(n161_adj_217), 
          .D0(n3142), .A1(n161_adj_344), .B1(n2273), .C1(n158_adj_216), 
          .D1(n3141), .CIN(n11821), .COUT(n11822), .S0(n161_adj_281), 
          .S1(n158_adj_280));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_606_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_606_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_606_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2273), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n11821));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_606_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_606_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_606_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_606_add_4_1.INJECT1_1 = "NO";
    CCU2C add_633_add_4_34 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11817), .S0(n1033));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_34.INIT0 = 16'hffff;
    defparam add_633_add_4_34.INIT1 = 16'h0000;
    defparam add_633_add_4_34.INJECT1_0 = "NO";
    defparam add_633_add_4_34.INJECT1_1 = "NO";
    CCU2C add_633_add_4_32 (.A0(det_q4_28[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11816), .COUT(n11817), .S0(n1035), .S1(n1034));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_32.INIT0 = 16'h5555;
    defparam add_633_add_4_32.INIT1 = 16'h5555;
    defparam add_633_add_4_32.INJECT1_0 = "NO";
    defparam add_633_add_4_32.INJECT1_1 = "NO";
    CCU2C add_633_add_4_30 (.A0(det_q4_28[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11815), .COUT(n11816), .S0(n1037), .S1(n1036));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_30.INIT0 = 16'h5555;
    defparam add_633_add_4_30.INIT1 = 16'h5555;
    defparam add_633_add_4_30.INJECT1_0 = "NO";
    defparam add_633_add_4_30.INJECT1_1 = "NO";
    CCU2C add_633_add_4_28 (.A0(det_q4_28[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11814), .COUT(n11815), .S0(n1039), .S1(n1038));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_28.INIT0 = 16'h5555;
    defparam add_633_add_4_28.INIT1 = 16'h5555;
    defparam add_633_add_4_28.INJECT1_0 = "NO";
    defparam add_633_add_4_28.INJECT1_1 = "NO";
    CCU2C add_633_add_4_26 (.A0(det_q4_28[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11813), .COUT(n11814), .S0(n1041), .S1(n1040));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_26.INIT0 = 16'h5555;
    defparam add_633_add_4_26.INIT1 = 16'h5555;
    defparam add_633_add_4_26.INJECT1_0 = "NO";
    defparam add_633_add_4_26.INJECT1_1 = "NO";
    CCU2C add_633_add_4_24 (.A0(det_q4_28[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11812), .COUT(n11813), .S0(n1043), .S1(n1042));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_24.INIT0 = 16'h5555;
    defparam add_633_add_4_24.INIT1 = 16'h5555;
    defparam add_633_add_4_24.INJECT1_0 = "NO";
    defparam add_633_add_4_24.INJECT1_1 = "NO";
    CCU2C add_633_add_4_22 (.A0(det_q4_28[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11811), .COUT(n11812), .S0(n1045), .S1(n1044));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_22.INIT0 = 16'h5555;
    defparam add_633_add_4_22.INIT1 = 16'h5555;
    defparam add_633_add_4_22.INJECT1_0 = "NO";
    defparam add_633_add_4_22.INJECT1_1 = "NO";
    CCU2C add_633_add_4_20 (.A0(det_q4_28[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11810), .COUT(n11811), .S0(n1047), .S1(n1046));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_20.INIT0 = 16'h5555;
    defparam add_633_add_4_20.INIT1 = 16'h5555;
    defparam add_633_add_4_20.INJECT1_0 = "NO";
    defparam add_633_add_4_20.INJECT1_1 = "NO";
    CCU2C add_633_add_4_18 (.A0(det_q4_28[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11809), .COUT(n11810), .S0(n1049), .S1(n1048));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_18.INIT0 = 16'h5555;
    defparam add_633_add_4_18.INIT1 = 16'h5555;
    defparam add_633_add_4_18.INJECT1_0 = "NO";
    defparam add_633_add_4_18.INJECT1_1 = "NO";
    CCU2C add_633_add_4_16 (.A0(det_q4_28[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11808), .COUT(n11809), .S0(n1051), .S1(n1050));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_16.INIT0 = 16'h5555;
    defparam add_633_add_4_16.INIT1 = 16'h5555;
    defparam add_633_add_4_16.INJECT1_0 = "NO";
    defparam add_633_add_4_16.INJECT1_1 = "NO";
    CCU2C add_633_add_4_14 (.A0(det_q4_28[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11807), .COUT(n11808), .S0(n1053), .S1(n1052));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_14.INIT0 = 16'h5555;
    defparam add_633_add_4_14.INIT1 = 16'h5555;
    defparam add_633_add_4_14.INJECT1_0 = "NO";
    defparam add_633_add_4_14.INJECT1_1 = "NO";
    CCU2C add_633_add_4_12 (.A0(det_q4_28[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11806), .COUT(n11807), .S0(n1055), .S1(n1054));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_12.INIT0 = 16'h5555;
    defparam add_633_add_4_12.INIT1 = 16'h5555;
    defparam add_633_add_4_12.INJECT1_0 = "NO";
    defparam add_633_add_4_12.INJECT1_1 = "NO";
    CCU2C add_633_add_4_10 (.A0(det_q4_28[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11805), .COUT(n11806), .S0(n1057), .S1(n1056));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_10.INIT0 = 16'h5555;
    defparam add_633_add_4_10.INIT1 = 16'h5555;
    defparam add_633_add_4_10.INJECT1_0 = "NO";
    defparam add_633_add_4_10.INJECT1_1 = "NO";
    CCU2C add_633_add_4_8 (.A0(det_q4_28[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11804), .COUT(n11805), .S0(n1059), .S1(n1058));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_8.INIT0 = 16'h5555;
    defparam add_633_add_4_8.INIT1 = 16'h5555;
    defparam add_633_add_4_8.INJECT1_0 = "NO";
    defparam add_633_add_4_8.INJECT1_1 = "NO";
    CCU2C add_633_add_4_6 (.A0(det_q4_28[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11803), .COUT(n11804), .S0(n1061), .S1(n1060));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_6.INIT0 = 16'h5555;
    defparam add_633_add_4_6.INIT1 = 16'h5555;
    defparam add_633_add_4_6.INJECT1_0 = "NO";
    defparam add_633_add_4_6.INJECT1_1 = "NO";
    CCU2C add_633_add_4_4 (.A0(det_q4_28[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n11802), .COUT(n11803), .S0(n1063), .S1(n1062));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_4.INIT0 = 16'h5555;
    defparam add_633_add_4_4.INIT1 = 16'h5555;
    defparam add_633_add_4_4.INJECT1_0 = "NO";
    defparam add_633_add_4_4.INJECT1_1 = "NO";
    CCU2C add_633_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(det_q4_28[1]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n11802), .S1(n1064));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam add_633_add_4_2.INIT0 = 16'h000f;
    defparam add_633_add_4_2.INIT1 = 16'h5555;
    defparam add_633_add_4_2.INJECT1_0 = "NO";
    defparam add_633_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_33 (.A0(n1067), .B0(n13005), .C0(n71_adj_441), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11801), .S0(n68_adj_345));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_597_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_597_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_31 (.A0(n77_adj_443), .B0(n13005), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_442), .B1(n13005), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11800), .COUT(n11801), .S0(n74_adj_347), 
          .S1(n71_adj_346));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_29 (.A0(n83_adj_445), .B0(n13005), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_444), .B1(n13005), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11799), .COUT(n11800), .S0(n80_adj_349), 
          .S1(n77_adj_348));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_27 (.A0(n89_adj_447), .B0(n13005), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_446), .B1(n13005), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11798), .COUT(n11799), .S0(n86_adj_351), 
          .S1(n83_adj_350));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_25 (.A0(n95_adj_449), .B0(n13005), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_448), .B1(n13005), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11797), .COUT(n11798), .S0(n92_adj_353), 
          .S1(n89_adj_352));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_23 (.A0(n101_adj_451), .B0(n13005), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_450), .B1(n13005), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11796), .COUT(n11797), .S0(n98_adj_355), 
          .S1(n95_adj_354));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_21 (.A0(n107_adj_453), .B0(n13005), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_452), .B1(n13005), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11795), .COUT(n11796), .S0(n104_adj_357), 
          .S1(n101_adj_356));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_19 (.A0(n113_adj_455), .B0(n13005), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_454), .B1(n13005), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11794), .COUT(n11795), .S0(n110_adj_359), 
          .S1(n107_adj_358));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_17 (.A0(n119_adj_457), .B0(n13005), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_456), .B1(n13005), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11793), .COUT(n11794), .S0(n116_adj_361), 
          .S1(n113_adj_360));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_15 (.A0(n125_adj_459), .B0(n13005), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_458), .B1(n13005), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11792), .COUT(n11793), .S0(n122_adj_363), 
          .S1(n119_adj_362));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_13 (.A0(n131_adj_461), .B0(n13005), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_460), .B1(n13005), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11791), .COUT(n11792), .S0(n128_adj_365), 
          .S1(n125_adj_364));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_11 (.A0(n137_adj_463), .B0(n13005), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_462), .B1(n13005), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11790), .COUT(n11791), .S0(n134_adj_367), 
          .S1(n131_adj_366));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_9 (.A0(n143_adj_465), .B0(n13005), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_464), .B1(n13005), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11789), .COUT(n11790), .S0(n140_adj_369), 
          .S1(n137_adj_368));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_7 (.A0(n149_adj_467), .B0(n13005), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_466), .B1(n13005), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11788), .COUT(n11789), .S0(n146_adj_371), 
          .S1(n143_adj_370));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_5 (.A0(n155_adj_469), .B0(n13005), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_468), .B1(n13005), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11787), .COUT(n11788), .S0(n152_adj_373), 
          .S1(n149_adj_372));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_3 (.A0(n161_adj_471), .B0(n13005), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_470), .B1(n13005), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11786), .COUT(n11787), .S0(n158_adj_375), 
          .S1(n155_adj_374));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_597_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_597_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13005), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11786), .S1(n161_adj_376));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_597_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_597_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_597_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_597_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_33 (.A0(n1067), .B0(n13005), .C0(n71_adj_473), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11785), .S0(n68_adj_377));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_594_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_594_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_31 (.A0(n77_adj_475), .B0(n13005), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_474), .B1(n13005), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11784), .COUT(n11785), .S0(n74_adj_379), 
          .S1(n71_adj_378));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_29 (.A0(n83_adj_477), .B0(n13005), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_476), .B1(n13005), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11783), .COUT(n11784), .S0(n80_adj_381), 
          .S1(n77_adj_380));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_27 (.A0(n89_adj_479), .B0(n13005), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_478), .B1(n13005), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11782), .COUT(n11783), .S0(n86_adj_383), 
          .S1(n83_adj_382));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_25 (.A0(n95_adj_481), .B0(n13005), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_480), .B1(n13005), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11781), .COUT(n11782), .S0(n92_adj_385), 
          .S1(n89_adj_384));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_23 (.A0(n101_adj_483), .B0(n13005), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_482), .B1(n13005), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11780), .COUT(n11781), .S0(n98_adj_387), 
          .S1(n95_adj_386));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_21 (.A0(n107_adj_485), .B0(n13005), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_484), .B1(n13005), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11779), .COUT(n11780), .S0(n104_adj_389), 
          .S1(n101_adj_388));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_19 (.A0(n113_adj_487), .B0(n13005), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_486), .B1(n13005), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11778), .COUT(n11779), .S0(n110_adj_391), 
          .S1(n107_adj_390));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_17 (.A0(n119_adj_489), .B0(n13005), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_488), .B1(n13005), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11777), .COUT(n11778), .S0(n116_adj_393), 
          .S1(n113_adj_392));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_15 (.A0(n125_adj_491), .B0(n13005), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_490), .B1(n13005), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11776), .COUT(n11777), .S0(n122_adj_395), 
          .S1(n119_adj_394));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_13 (.A0(n131_adj_493), .B0(n13005), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_492), .B1(n13005), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11775), .COUT(n11776), .S0(n128_adj_397), 
          .S1(n125_adj_396));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_11 (.A0(n137_adj_495), .B0(n13005), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_494), .B1(n13005), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11774), .COUT(n11775), .S0(n134_adj_399), 
          .S1(n131_adj_398));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_9 (.A0(n143_adj_497), .B0(n13005), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_496), .B1(n13005), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11773), .COUT(n11774), .S0(n140_adj_401), 
          .S1(n137_adj_400));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_7 (.A0(n149_adj_499), .B0(n13005), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_498), .B1(n13005), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11772), .COUT(n11773), .S0(n146_adj_403), 
          .S1(n143_adj_402));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_5 (.A0(n155_adj_501), .B0(n13005), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_500), .B1(n13005), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11771), .COUT(n11772), .S0(n152_adj_405), 
          .S1(n149_adj_404));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_3 (.A0(n161_adj_503), .B0(n13005), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_502), .B1(n13005), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11770), .COUT(n11771), .S0(n158_adj_407), 
          .S1(n155_adj_406));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_594_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_594_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13005), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11770), .S1(n161_adj_408));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_594_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_594_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_594_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_594_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_33 (.A0(n74_adj_1177), .B0(n2139), .C0(n71), .D0(n2241), 
          .A1(n71_adj_1176), .B1(n2139), .C1(n68_adj_169), .D1(n2240), 
          .CIN(n11768), .S0(n71_adj_409), .S1(n2273));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_33.INIT0 = 16'h74b8;
    defparam _add_1_add_4_33.INIT1 = 16'h74b8;
    defparam _add_1_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_31 (.A0(n80_adj_1179), .B0(n2139), .C0(n77), .D0(n2243), 
          .A1(n77_adj_1178), .B1(n2139), .C1(n74), .D1(n2242), .CIN(n11767), 
          .COUT(n11768), .S0(n77_adj_411), .S1(n74_adj_410));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_31.INIT0 = 16'h74b8;
    defparam _add_1_add_4_31.INIT1 = 16'h74b8;
    defparam _add_1_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_29 (.A0(n86_adj_1181), .B0(n2139), .C0(n83), .D0(n2245), 
          .A1(n83_adj_1180), .B1(n2139), .C1(n80), .D1(n2244), .CIN(n11766), 
          .COUT(n11767), .S0(n83_adj_413), .S1(n80_adj_412));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_29.INIT0 = 16'h74b8;
    defparam _add_1_add_4_29.INIT1 = 16'h74b8;
    defparam _add_1_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_27 (.A0(n92_adj_1183), .B0(n2139), .C0(n89), .D0(n2247), 
          .A1(n89_adj_1182), .B1(n2139), .C1(n86), .D1(n2246), .CIN(n11765), 
          .COUT(n11766), .S0(n89_adj_415), .S1(n86_adj_414));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_27.INIT0 = 16'h74b8;
    defparam _add_1_add_4_27.INIT1 = 16'h74b8;
    defparam _add_1_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_25 (.A0(n98_adj_1185), .B0(n2139), .C0(n95), .D0(n2249), 
          .A1(n95_adj_1184), .B1(n2139), .C1(n92), .D1(n2248), .CIN(n11764), 
          .COUT(n11765), .S0(n95_adj_417), .S1(n92_adj_416));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_25.INIT0 = 16'h74b8;
    defparam _add_1_add_4_25.INIT1 = 16'h74b8;
    defparam _add_1_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_23 (.A0(n104_adj_1187), .B0(n2139), .C0(n101), 
          .D0(n2251), .A1(n101_adj_1186), .B1(n2139), .C1(n98), .D1(n2250), 
          .CIN(n11763), .COUT(n11764), .S0(n101_adj_419), .S1(n98_adj_418));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_23.INIT0 = 16'h74b8;
    defparam _add_1_add_4_23.INIT1 = 16'h74b8;
    defparam _add_1_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_21 (.A0(n110_adj_1189), .B0(n2139), .C0(n107), 
          .D0(n2253), .A1(n107_adj_1188), .B1(n2139), .C1(n104_adj_168), 
          .D1(n2252), .CIN(n11762), .COUT(n11763), .S0(n107_adj_421), 
          .S1(n104_adj_420));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_21.INIT0 = 16'h74b8;
    defparam _add_1_add_4_21.INIT1 = 16'h74b8;
    defparam _add_1_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_19 (.A0(n116_adj_1191), .B0(n2139), .C0(n113), 
          .D0(n2255), .A1(n113_adj_1190), .B1(n2139), .C1(n110_adj_167), 
          .D1(n2254), .CIN(n11761), .COUT(n11762), .S0(n113_adj_423), 
          .S1(n110_adj_422));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_19.INIT0 = 16'h74b8;
    defparam _add_1_add_4_19.INIT1 = 16'h74b8;
    defparam _add_1_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_17 (.A0(n122_adj_1193), .B0(n2139), .C0(n119), 
          .D0(n2257), .A1(n119_adj_1192), .B1(n2139), .C1(n116_adj_166), 
          .D1(n2256), .CIN(n11760), .COUT(n11761), .S0(n119_adj_425), 
          .S1(n116_adj_424));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_17.INIT0 = 16'h74b8;
    defparam _add_1_add_4_17.INIT1 = 16'h74b8;
    defparam _add_1_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_15 (.A0(n128_adj_1195), .B0(n2139), .C0(n125), 
          .D0(n2259), .A1(n125_adj_1194), .B1(n2139), .C1(n122_adj_165), 
          .D1(n2258), .CIN(n11759), .COUT(n11760), .S0(n125_adj_427), 
          .S1(n122_adj_426));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_15.INIT0 = 16'h74b8;
    defparam _add_1_add_4_15.INIT1 = 16'h74b8;
    defparam _add_1_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_13 (.A0(n134_adj_1197), .B0(n2139), .C0(n131), 
          .D0(n2261), .A1(n131_adj_1196), .B1(n2139), .C1(n128_adj_164), 
          .D1(n2260), .CIN(n11758), .COUT(n11759), .S0(n131_adj_429), 
          .S1(n128_adj_428));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_13.INIT0 = 16'h74b8;
    defparam _add_1_add_4_13.INIT1 = 16'h74b8;
    defparam _add_1_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_11 (.A0(n140_adj_1199), .B0(n2139), .C0(n137), 
          .D0(n2263), .A1(n137_adj_1198), .B1(n2139), .C1(n134), .D1(n2262), 
          .CIN(n11757), .COUT(n11758), .S0(n137_adj_431), .S1(n134_adj_430));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_11.INIT0 = 16'h74b8;
    defparam _add_1_add_4_11.INIT1 = 16'h74b8;
    defparam _add_1_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_9 (.A0(n146_adj_1201), .B0(n2139), .C0(n143), .D0(n2265), 
          .A1(n143_adj_1200), .B1(n2139), .C1(n140), .D1(n2264), .CIN(n11756), 
          .COUT(n11757), .S0(n143_adj_433), .S1(n140_adj_432));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_9.INIT0 = 16'h74b8;
    defparam _add_1_add_4_9.INIT1 = 16'h74b8;
    defparam _add_1_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_7 (.A0(n152_adj_1203), .B0(n2139), .C0(n149), .D0(n2267), 
          .A1(n149_adj_1202), .B1(n2139), .C1(n146), .D1(n2266), .CIN(n11755), 
          .COUT(n11756), .S0(n149_adj_435), .S1(n146_adj_434));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_7.INIT0 = 16'h74b8;
    defparam _add_1_add_4_7.INIT1 = 16'h74b8;
    defparam _add_1_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_5 (.A0(n158_adj_1205), .B0(n2139), .C0(n155), .D0(n2269), 
          .A1(n155_adj_1204), .B1(n2139), .C1(n152), .D1(n2268), .CIN(n11754), 
          .COUT(n11755), .S0(n155_adj_437), .S1(n152_adj_436));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_5.INIT0 = 16'h74b8;
    defparam _add_1_add_4_5.INIT1 = 16'h74b8;
    defparam _add_1_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_3 (.A0(det_q4_28[0]), .B0(n2139), .C0(n161), .D0(n2271), 
          .A1(n161_adj_791), .B1(n2139), .C1(n158), .D1(n2270), .CIN(n11753), 
          .COUT(n11754), .S0(n161_adj_439), .S1(n158_adj_438));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_3.INIT0 = 16'h74b8;
    defparam _add_1_add_4_3.INIT1 = 16'h74b8;
    defparam _add_1_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n2139), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .COUT(n11753));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_33 (.A0(n1067), .B0(n13006), .C0(n71_adj_505), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11749), .S0(n68_adj_440));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_591_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_591_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_31 (.A0(n77_adj_507), .B0(n13006), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_506), .B1(n13006), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11748), .COUT(n11749), .S0(n74_adj_442), 
          .S1(n71_adj_441));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_29 (.A0(n83_adj_509), .B0(n13006), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_508), .B1(n13006), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11747), .COUT(n11748), .S0(n80_adj_444), 
          .S1(n77_adj_443));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_27 (.A0(n89_adj_511), .B0(n13006), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_510), .B1(n13006), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11746), .COUT(n11747), .S0(n86_adj_446), 
          .S1(n83_adj_445));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_25 (.A0(n95_adj_513), .B0(n13006), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_512), .B1(n13006), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11745), .COUT(n11746), .S0(n92_adj_448), 
          .S1(n89_adj_447));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_23 (.A0(n101_adj_515), .B0(n13006), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_514), .B1(n13006), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11744), .COUT(n11745), .S0(n98_adj_450), 
          .S1(n95_adj_449));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_21 (.A0(n107_adj_517), .B0(n13006), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_516), .B1(n13006), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11743), .COUT(n11744), .S0(n104_adj_452), 
          .S1(n101_adj_451));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_19 (.A0(n113_adj_519), .B0(n13006), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_518), .B1(n13006), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11742), .COUT(n11743), .S0(n110_adj_454), 
          .S1(n107_adj_453));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_17 (.A0(n119_adj_521), .B0(n13006), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_520), .B1(n13006), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11741), .COUT(n11742), .S0(n116_adj_456), 
          .S1(n113_adj_455));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_15 (.A0(n125_adj_523), .B0(n13006), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_522), .B1(n13006), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11740), .COUT(n11741), .S0(n122_adj_458), 
          .S1(n119_adj_457));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_13 (.A0(n131_adj_525), .B0(n13006), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_524), .B1(n13006), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11739), .COUT(n11740), .S0(n128_adj_460), 
          .S1(n125_adj_459));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_11 (.A0(n137_adj_527), .B0(n13006), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_526), .B1(n13006), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11738), .COUT(n11739), .S0(n134_adj_462), 
          .S1(n131_adj_461));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_9 (.A0(n143_adj_529), .B0(n13006), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_528), .B1(n13006), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11737), .COUT(n11738), .S0(n140_adj_464), 
          .S1(n137_adj_463));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_7 (.A0(n149_adj_531), .B0(n13006), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_530), .B1(n13006), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11736), .COUT(n11737), .S0(n146_adj_466), 
          .S1(n143_adj_465));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_5 (.A0(n155_adj_533), .B0(n13006), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_532), .B1(n13006), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11735), .COUT(n11736), .S0(n152_adj_468), 
          .S1(n149_adj_467));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_3 (.A0(n161_adj_535), .B0(n13006), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_534), .B1(n13006), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11734), .COUT(n11735), .S0(n158_adj_470), 
          .S1(n155_adj_469));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_591_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_591_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13006), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11734), .S1(n161_adj_471));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_591_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_591_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_591_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_591_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_33 (.A0(n1067), .B0(n13006), .C0(n71_adj_537), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11733), .S0(n68_adj_472));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_588_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_588_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_31 (.A0(n77_adj_539), .B0(n13006), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_538), .B1(n13006), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11732), .COUT(n11733), .S0(n74_adj_474), 
          .S1(n71_adj_473));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_29 (.A0(n83_adj_541), .B0(n13006), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_540), .B1(n13006), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11731), .COUT(n11732), .S0(n80_adj_476), 
          .S1(n77_adj_475));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_27 (.A0(n89_adj_543), .B0(n13006), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_542), .B1(n13006), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11730), .COUT(n11731), .S0(n86_adj_478), 
          .S1(n83_adj_477));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_25 (.A0(n95_adj_545), .B0(n13006), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_544), .B1(n13006), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11729), .COUT(n11730), .S0(n92_adj_480), 
          .S1(n89_adj_479));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_23 (.A0(n101_adj_547), .B0(n13006), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_546), .B1(n13006), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11728), .COUT(n11729), .S0(n98_adj_482), 
          .S1(n95_adj_481));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_21 (.A0(n107_adj_549), .B0(n13006), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_548), .B1(n13006), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11727), .COUT(n11728), .S0(n104_adj_484), 
          .S1(n101_adj_483));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_19 (.A0(n113_adj_551), .B0(n13006), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_550), .B1(n13006), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11726), .COUT(n11727), .S0(n110_adj_486), 
          .S1(n107_adj_485));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_17 (.A0(n119_adj_553), .B0(n13006), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_552), .B1(n13006), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11725), .COUT(n11726), .S0(n116_adj_488), 
          .S1(n113_adj_487));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_15 (.A0(n125_adj_555), .B0(n13006), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_554), .B1(n13006), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11724), .COUT(n11725), .S0(n122_adj_490), 
          .S1(n119_adj_489));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_13 (.A0(n131_adj_557), .B0(n13006), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_556), .B1(n13006), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11723), .COUT(n11724), .S0(n128_adj_492), 
          .S1(n125_adj_491));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_11 (.A0(n137_adj_559), .B0(n13006), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_558), .B1(n13006), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11722), .COUT(n11723), .S0(n134_adj_494), 
          .S1(n131_adj_493));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_9 (.A0(n143_adj_561), .B0(n13006), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_560), .B1(n13006), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11721), .COUT(n11722), .S0(n140_adj_496), 
          .S1(n137_adj_495));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_7 (.A0(n149_adj_563), .B0(n13006), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_562), .B1(n13006), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11720), .COUT(n11721), .S0(n146_adj_498), 
          .S1(n143_adj_497));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_5 (.A0(n155_adj_565), .B0(n13006), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_564), .B1(n13006), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11719), .COUT(n11720), .S0(n152_adj_500), 
          .S1(n149_adj_499));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_3 (.A0(n161_adj_567), .B0(n13006), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_566), .B1(n13006), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11718), .COUT(n11719), .S0(n158_adj_502), 
          .S1(n155_adj_501));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_588_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_588_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13006), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11718), .S1(n161_adj_503));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_588_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_588_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_588_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_588_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_33 (.A0(n1067), .B0(n13004), .C0(n71_adj_346), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11717), .S0(n68_adj_282));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_603_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_603_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_31 (.A0(n77_adj_348), .B0(n13004), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_347), .B1(n13004), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11716), .COUT(n11717), .S0(n74_adj_284), 
          .S1(n71_adj_283));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_29 (.A0(n83_adj_350), .B0(n13004), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_349), .B1(n13004), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11715), .COUT(n11716), .S0(n80_adj_286), 
          .S1(n77_adj_285));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_29.INJECT1_1 = "NO";
    FD1S3AX d_reg_15__I_0_e2__i3 (.D(d_c_2), .CK(clk_c), .Q(n126_adj_173));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i3.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i4 (.D(d_c_3), .CK(clk_c), .Q(n124_adj_174));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i4.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i5 (.D(d_c_4), .CK(clk_c), .Q(n122_adj_175));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i5.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i6 (.D(d_c_5), .CK(clk_c), .Q(n120_adj_176));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i6.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i7 (.D(d_c_6), .CK(clk_c), .Q(n118_adj_177));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i7.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i8 (.D(d_c_7), .CK(clk_c), .Q(n116_adj_178));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i8.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i9 (.D(d_c_8), .CK(clk_c), .Q(n114_adj_179));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i9.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i10 (.D(d_c_9), .CK(clk_c), .Q(n112_adj_180));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i10.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i11 (.D(d_c_10), .CK(clk_c), .Q(n110_adj_181));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i11.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i12 (.D(d_c_11), .CK(clk_c), .Q(n108_adj_182));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i12.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i13 (.D(d_c_12), .CK(clk_c), .Q(n106_adj_183));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i13.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i14 (.D(d_c_13), .CK(clk_c), .Q(n104_adj_184));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i14.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i15 (.D(d_c_14), .CK(clk_c), .Q(n102_adj_170));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i15.GSR = "ENABLED";
    FD1S3AX d_reg_15__I_0_e2__i16 (.D(d_c_15), .CK(clk_c), .Q(n68_adj_185));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(84[44:57])
    defparam d_reg_15__I_0_e2__i16.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i2 (.D(a_c_1), .CK(clk_c), .Q(n128));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i2.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i3 (.D(a_c_2), .CK(clk_c), .Q(n126));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i3.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i4 (.D(a_c_3), .CK(clk_c), .Q(n124));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i4.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i5 (.D(a_c_4), .CK(clk_c), .Q(n122));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i5.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i6 (.D(a_c_5), .CK(clk_c), .Q(n120));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i6.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i7 (.D(a_c_6), .CK(clk_c), .Q(n118));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i7.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i8 (.D(a_c_7), .CK(clk_c), .Q(n116));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i8.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i9 (.D(a_c_8), .CK(clk_c), .Q(n114));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i9.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i10 (.D(a_c_9), .CK(clk_c), .Q(n112));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i10.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i11 (.D(a_c_10), .CK(clk_c), .Q(n110));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i11.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i12 (.D(a_c_11), .CK(clk_c), .Q(n108));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i12.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i13 (.D(a_c_12), .CK(clk_c), .Q(n106));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i13.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i14 (.D(a_c_13), .CK(clk_c), .Q(n104));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i14.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i15 (.D(a_c_14), .CK(clk_c), .Q(n102));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i15.GSR = "ENABLED";
    FD1S3AX a_reg_15__I_0_e2__i16 (.D(a_c_15), .CK(clk_c), .Q(n68));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(87[44:57])
    defparam a_reg_15__I_0_e2__i16.GSR = "ENABLED";
    LUT4 i1356_2_lut_4_lut (.A(n68_adj_1110), .B(n68_adj_1078), .C(n1033), 
         .D(det_zero), .Z(n35)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1356_2_lut_4_lut.init = 16'h0035;
    FD1S3AX c_reg_i0 (.D(c_c_0), .CK(clk_c), .Q(c_reg[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(41[18] 49[12])
    defparam c_reg_i0.GSR = "ENABLED";
    CCU2C _add_1_603_add_4_27 (.A0(n89_adj_352), .B0(n13004), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_351), .B1(n13004), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11714), .COUT(n11715), .S0(n86_adj_288), 
          .S1(n83_adj_287));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_25 (.A0(n95_adj_354), .B0(n13004), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_353), .B1(n13004), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11713), .COUT(n11714), .S0(n92_adj_290), 
          .S1(n89_adj_289));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_23 (.A0(n101_adj_356), .B0(n13004), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_355), .B1(n13004), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11712), .COUT(n11713), .S0(n98_adj_292), 
          .S1(n95_adj_291));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_21 (.A0(n107_adj_358), .B0(n13004), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_357), .B1(n13004), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11711), .COUT(n11712), .S0(n104_adj_294), 
          .S1(n101_adj_293));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_19 (.A0(n113_adj_360), .B0(n13004), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_359), .B1(n13004), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11710), .COUT(n11711), .S0(n110_adj_296), 
          .S1(n107_adj_295));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_17 (.A0(n119_adj_362), .B0(n13004), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_361), .B1(n13004), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11709), .COUT(n11710), .S0(n116_adj_298), 
          .S1(n113_adj_297));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_15 (.A0(n125_adj_364), .B0(n13004), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_363), .B1(n13004), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11708), .COUT(n11709), .S0(n122_adj_300), 
          .S1(n119_adj_299));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_13 (.A0(n131_adj_366), .B0(n13004), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_365), .B1(n13004), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11707), .COUT(n11708), .S0(n128_adj_302), 
          .S1(n125_adj_301));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_11 (.A0(n137_adj_368), .B0(n13004), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_367), .B1(n13004), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11706), .COUT(n11707), .S0(n134_adj_304), 
          .S1(n131_adj_303));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_9 (.A0(n143_adj_370), .B0(n13004), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_369), .B1(n13004), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11705), .COUT(n11706), .S0(n140_adj_306), 
          .S1(n137_adj_305));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_7 (.A0(n149_adj_372), .B0(n13004), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_371), .B1(n13004), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11704), .COUT(n11705), .S0(n146_adj_308), 
          .S1(n143_adj_307));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_5 (.A0(n155_adj_374), .B0(n13004), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_373), .B1(n13004), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11703), .COUT(n11704), .S0(n152_adj_310), 
          .S1(n149_adj_309));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_3 (.A0(n161_adj_376), .B0(n13004), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_375), .B1(n13004), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11702), .COUT(n11703), .S0(n158_adj_312), 
          .S1(n155_adj_311));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_603_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_603_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13004), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11702), .S1(n161_adj_313));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_603_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_603_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_603_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_603_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_33 (.A0(n1067), .B0(n13007), .C0(n71_adj_569), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11701), .S0(n68_adj_504));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_585_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_585_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_31 (.A0(n77_adj_571), .B0(n13007), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_570), .B1(n13007), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11700), .COUT(n11701), .S0(n74_adj_506), 
          .S1(n71_adj_505));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_29 (.A0(n83_adj_573), .B0(n13007), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_572), .B1(n13007), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11699), .COUT(n11700), .S0(n80_adj_508), 
          .S1(n77_adj_507));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_27 (.A0(n89_adj_575), .B0(n13007), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_574), .B1(n13007), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11698), .COUT(n11699), .S0(n86_adj_510), 
          .S1(n83_adj_509));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_25 (.A0(n95_adj_577), .B0(n13007), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_576), .B1(n13007), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11697), .COUT(n11698), .S0(n92_adj_512), 
          .S1(n89_adj_511));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_23 (.A0(n101_adj_579), .B0(n13007), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_578), .B1(n13007), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11696), .COUT(n11697), .S0(n98_adj_514), 
          .S1(n95_adj_513));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_21 (.A0(n107_adj_581), .B0(n13007), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_580), .B1(n13007), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11695), .COUT(n11696), .S0(n104_adj_516), 
          .S1(n101_adj_515));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_19 (.A0(n113_adj_583), .B0(n13007), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_582), .B1(n13007), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11694), .COUT(n11695), .S0(n110_adj_518), 
          .S1(n107_adj_517));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_17 (.A0(n119_adj_585), .B0(n13007), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_584), .B1(n13007), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11693), .COUT(n11694), .S0(n116_adj_520), 
          .S1(n113_adj_519));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_15 (.A0(n125_adj_587), .B0(n13007), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_586), .B1(n13007), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11692), .COUT(n11693), .S0(n122_adj_522), 
          .S1(n119_adj_521));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_13 (.A0(n131_adj_589), .B0(n13007), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_588), .B1(n13007), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11691), .COUT(n11692), .S0(n128_adj_524), 
          .S1(n125_adj_523));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_11 (.A0(n137_adj_591), .B0(n13007), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_590), .B1(n13007), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11690), .COUT(n11691), .S0(n134_adj_526), 
          .S1(n131_adj_525));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_9 (.A0(n143_adj_593), .B0(n13007), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_592), .B1(n13007), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11689), .COUT(n11690), .S0(n140_adj_528), 
          .S1(n137_adj_527));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_7 (.A0(n149_adj_595), .B0(n13007), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_594), .B1(n13007), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11688), .COUT(n11689), .S0(n146_adj_530), 
          .S1(n143_adj_529));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_5 (.A0(n155_adj_597), .B0(n13007), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_596), .B1(n13007), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11687), .COUT(n11688), .S0(n152_adj_532), 
          .S1(n149_adj_531));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_3 (.A0(n161_adj_599), .B0(n13007), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_598), .B1(n13007), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11686), .COUT(n11687), .S0(n158_adj_534), 
          .S1(n155_adj_533));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_585_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_585_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13007), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11686), .S1(n161_adj_535));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_585_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_585_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_585_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_585_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_300_i1_3_lut_rep_91 (.A(n68_adj_1713), .B(n68_adj_1554), .C(n1033), 
         .Z(n13027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_300_i1_3_lut_rep_91.init = 16'hcaca;
    LUT4 i1359_2_lut_4_lut (.A(n68_adj_1713), .B(n68_adj_1554), .C(n1033), 
         .D(det_zero), .Z(n34)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1359_2_lut_4_lut.init = 16'h0035;
    LUT4 mux_299_i1_3_lut_rep_92 (.A(n68_adj_2066), .B(n68_adj_1874), .C(n1033), 
         .Z(n13028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_299_i1_3_lut_rep_92.init = 16'hcaca;
    LUT4 i1368_2_lut_4_lut (.A(n68_adj_2066), .B(n68_adj_1874), .C(n1033), 
         .D(det_zero), .Z(n33)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i1368_2_lut_4_lut.init = 16'h0035;
    VLO i1 (.Z(GND_net));
    reciprocal_q16_16 u_recip (.error_recip(error_recip), .clk_c(clk_c), 
            .det_zero(det_zero), .n1081(n1081), .det_q4_28({det_q4_28}), 
            .n13023(n13023), .n1517(n1517), .n1080(n1080), .n1516(n1516), 
            .n1079(n1079), .n1515(n1515), .n1078(n1078), .n1514(n1514), 
            .n1077(n1077), .n1513(n1513), .n1076(n1076), .n1512(n1512), 
            .n1075(n1075), .n1511(n1511), .n1092(n1092), .n13016(n13016), 
            .n2064(n2064), .n1091(n1091), .n2063(n2063), .n1074(n1074), 
            .n1510(n1510), .n1073(n1073), .n1509(n1509), .n1072(n1072), 
            .n1508(n1508), .n1071(n1071), .n1507(n1507), .n1070(n1070), 
            .n1506(n1506), .n1090(n1090), .n2062(n2062), .n1069(n1069), 
            .n1505(n1505), .n1068(n1068), .n1504(n1504), .n1098(n1098), 
            .n2070(n2070), .n1097(n1097), .n2069(n2069), .n1089(n1089), 
            .n2061(n2061), .n1096(n1096), .n2068(n2068), .n1095(n1095), 
            .n2067(n2067), .n1094(n1094), .n2066(n2066), .n1088(n1088), 
            .n2060(n2060), .n1087(n1087), .n2059(n2059), .n1086(n1086), 
            .n2058(n2058), .n1085(n1085), .n2057(n2057), .n1084(n1084), 
            .n2056(n2056), .n1083(n1083), .n2055(n2055), .n1082(n1082), 
            .n2054(n2054), .n2053(n2053), .n2052(n2052), .n2051(n2051), 
            .n2050(n2050), .n2049(n2049), .n2048(n2048), .n2047(n2047), 
            .n2046(n2046), .n2045(n2045), .n2044(n2044), .n2043(n2043), 
            .n2042(n2042), .n2041(n2041), .n2040(n2040), .n1093(n1093), 
            .n2065(n2065), .n3077(n3077), .n3110({n3111, n3112, n3113, 
            n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
            n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
            n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, 
            n3138, n3139, n3140, n3141, n3142}), .n1067(n1067), 
            .n13015(n13015), .n2241(n2241), .n2243(n2243), .n2242(n2242), 
            .n2245(n2245), .n2244(n2244), .n2247(n2247), .n2246(n2246), 
            .n2249(n2249), .n2248(n2248), .n2251(n2251), .n2250(n2250), 
            .n2253(n2253), .n2252(n2252), .n2255(n2255), .n2254(n2254), 
            .n2257(n2257), .n2256(n2256), .n2259(n2259), .n2258(n2258), 
            .n2261(n2261), .n2260(n2260), .n2263(n2263), .n2262(n2262), 
            .n2265(n2265), .n2264(n2264), .n2267(n2267), .n2266(n2266), 
            .n2269(n2269), .n2268(n2268), .n2271(n2271), .n2270(n2270), 
            .n13004(n13004), .n3075(n3075), .n3074(n3074), .n3073(n3073), 
            .n3072(n3072), .n3071(n3071), .n3070(n3070), .n3069(n3069), 
            .n3068(n3068), .n3067(n3067), .n3066(n3066), .n3065(n3065), 
            .n3064(n3064), .n3063(n3063), .n3062(n3062), .n3061(n3061), 
            .n3060(n3060), .n3059(n3059), .n3058(n3058), .n3057(n3057), 
            .n3056(n3056), .n3055(n3055), .n3054(n3054), .n3053(n3053), 
            .n3052(n3052), .n3051(n3051), .n3050(n3050), .n3049(n3049), 
            .n3048(n3048), .n1536(n1536), .n39(n39), .n68(n68_adj_1777), 
            .n68_adj_1(n68_adj_1142), .n68_adj_2(n68_adj_250), .n64(n64), 
            .n63(n63), .n62(n62), .n3047(n3047), .n3046(n3046), .n3045(n3045), 
            .n1534(n1534), .n1533(n1533), .n1532(n1532), .n1531(n1531), 
            .n1530(n1530), .n1529(n1529), .n1528(n1528), .n1527(n1527), 
            .n1526(n1526), .n1525(n1525), .n1524(n1524), .n1523(n1523), 
            .n1522(n1522), .n1521(n1521), .n2273(n2273), .n50(n50), 
            .n2139(n2139), .n48(n48), .n2072(n2072), .n47(n47), .GND_net(GND_net), 
            .n1520(n1520), .n1519(n1519), .n1518(n1518), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(61[23] 67[6])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2C _add_1_612_add_4_3 (.A0(n161_adj_1174), .B0(n13015), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1173), .B1(n13015), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11870), .COUT(n11871), .S0(n158), .S1(n155));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_5 (.A0(n155_adj_1172), .B0(n13015), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1171), .B1(n13015), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11871), .COUT(n11872), .S0(n152), .S1(n149));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_7 (.A0(n149_adj_1170), .B0(n13015), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1169), .B1(n13015), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11872), .COUT(n11873), .S0(n146), .S1(n143));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_9 (.A0(n143_adj_1168), .B0(n13015), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1167), .B1(n13015), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11873), .COUT(n11874), .S0(n140), .S1(n137));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_11 (.A0(n137_adj_1166), .B0(n13015), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1165), .B1(n13015), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11874), .COUT(n11875), .S0(n134), .S1(n131));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_13 (.A0(n131_adj_1164), .B0(n13015), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1163), .B1(n13015), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11875), .COUT(n11876), .S0(n128_adj_164), 
          .S1(n125));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_15 (.A0(n125_adj_1162), .B0(n13015), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1161), .B1(n13015), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11876), .COUT(n11877), .S0(n122_adj_165), 
          .S1(n119));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_17 (.A0(n119_adj_1160), .B0(n13015), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1159), .B1(n13015), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11877), .COUT(n11878), .S0(n116_adj_166), 
          .S1(n113));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_19 (.A0(n113_adj_1158), .B0(n13015), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1157), .B1(n13015), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11878), .COUT(n11879), .S0(n110_adj_167), 
          .S1(n107));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_21 (.A0(n107_adj_1156), .B0(n13015), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1155), .B1(n13015), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11879), .COUT(n11880), .S0(n104_adj_168), 
          .S1(n101));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_23 (.A0(n101_adj_1154), .B0(n13015), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1153), .B1(n13015), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11880), .COUT(n11881), .S0(n98), .S1(n95));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_25 (.A0(n95_adj_1152), .B0(n13015), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1151), .B1(n13015), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11881), .COUT(n11882), .S0(n92), .S1(n89));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_27 (.A0(n89_adj_1150), .B0(n13015), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1149), .B1(n13015), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11882), .COUT(n11883), .S0(n86), .S1(n83));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_29 (.A0(n83_adj_1148), .B0(n13015), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1147), .B1(n13015), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11883), .COUT(n11884), .S0(n80), .S1(n77));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_31 (.A0(n77_adj_1146), .B0(n13015), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1145), .B1(n13015), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11884), .COUT(n11885), .S0(n74), .S1(n71));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_612_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_612_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_612_add_4_33 (.A0(n1067), .B0(n13015), .C0(n71_adj_1144), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11885), .S0(n68_adj_169));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_612_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_612_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_612_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_612_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2273), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n11889));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_600_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_600_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_3 (.A0(n3075), .B0(n2273), .C0(det_q4_28[0]), 
          .D0(VCC_net), .A1(n3074), .B1(n2273), .C1(n161_adj_408), .D1(VCC_net), 
          .CIN(n11889), .COUT(n11890), .S0(n161_adj_344), .S1(n158_adj_343));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_3.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_3.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_5 (.A0(n3073), .B0(n2273), .C0(n158_adj_407), 
          .D0(VCC_net), .A1(n3072), .B1(n2273), .C1(n155_adj_406), .D1(VCC_net), 
          .CIN(n11890), .COUT(n11891), .S0(n155_adj_342), .S1(n152_adj_341));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_5.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_5.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_7 (.A0(n3071), .B0(n2273), .C0(n152_adj_405), 
          .D0(VCC_net), .A1(n3070), .B1(n2273), .C1(n149_adj_404), .D1(VCC_net), 
          .CIN(n11891), .COUT(n11892), .S0(n149_adj_340), .S1(n146_adj_339));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_7.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_7.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_9 (.A0(n3069), .B0(n2273), .C0(n146_adj_403), 
          .D0(VCC_net), .A1(n3068), .B1(n2273), .C1(n143_adj_402), .D1(VCC_net), 
          .CIN(n11892), .COUT(n11893), .S0(n143_adj_338), .S1(n140_adj_337));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_9.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_9.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_11 (.A0(n3067), .B0(n2273), .C0(n140_adj_401), 
          .D0(VCC_net), .A1(n3066), .B1(n2273), .C1(n137_adj_400), .D1(VCC_net), 
          .CIN(n11893), .COUT(n11894), .S0(n137_adj_336), .S1(n134_adj_335));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_11.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_11.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_13 (.A0(n3065), .B0(n2273), .C0(n134_adj_399), 
          .D0(VCC_net), .A1(n3064), .B1(n2273), .C1(n131_adj_398), .D1(VCC_net), 
          .CIN(n11894), .COUT(n11895), .S0(n131_adj_334), .S1(n128_adj_333));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_13.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_13.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_15 (.A0(n3063), .B0(n2273), .C0(n128_adj_397), 
          .D0(VCC_net), .A1(n3062), .B1(n2273), .C1(n125_adj_396), .D1(VCC_net), 
          .CIN(n11895), .COUT(n11896), .S0(n125_adj_332), .S1(n122_adj_331));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_15.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_15.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_17 (.A0(n3061), .B0(n2273), .C0(n122_adj_395), 
          .D0(VCC_net), .A1(n3060), .B1(n2273), .C1(n119_adj_394), .D1(VCC_net), 
          .CIN(n11896), .COUT(n11897), .S0(n119_adj_330), .S1(n116_adj_329));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_17.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_17.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_19 (.A0(n3059), .B0(n2273), .C0(n116_adj_393), 
          .D0(VCC_net), .A1(n3058), .B1(n2273), .C1(n113_adj_392), .D1(VCC_net), 
          .CIN(n11897), .COUT(n11898), .S0(n113_adj_328), .S1(n110_adj_327));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_19.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_19.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_21 (.A0(n3057), .B0(n2273), .C0(n110_adj_391), 
          .D0(VCC_net), .A1(n3056), .B1(n2273), .C1(n107_adj_390), .D1(VCC_net), 
          .CIN(n11898), .COUT(n11899), .S0(n107_adj_326), .S1(n104_adj_325));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_21.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_21.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_23 (.A0(n3055), .B0(n2273), .C0(n104_adj_389), 
          .D0(VCC_net), .A1(n3054), .B1(n2273), .C1(n101_adj_388), .D1(VCC_net), 
          .CIN(n11899), .COUT(n11900), .S0(n101_adj_324), .S1(n98_adj_323));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_23.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_23.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_25 (.A0(n3053), .B0(n2273), .C0(n98_adj_387), 
          .D0(VCC_net), .A1(n3052), .B1(n2273), .C1(n95_adj_386), .D1(VCC_net), 
          .CIN(n11900), .COUT(n11901), .S0(n95_adj_322), .S1(n92_adj_321));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_25.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_25.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_27 (.A0(n3051), .B0(n2273), .C0(n92_adj_385), 
          .D0(VCC_net), .A1(n3050), .B1(n2273), .C1(n89_adj_384), .D1(VCC_net), 
          .CIN(n11901), .COUT(n11902), .S0(n89_adj_320), .S1(n86_adj_319));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_27.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_27.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_29 (.A0(n3049), .B0(n2273), .C0(n86_adj_383), 
          .D0(VCC_net), .A1(n3048), .B1(n2273), .C1(n83_adj_382), .D1(VCC_net), 
          .CIN(n11902), .COUT(n11903), .S0(n83_adj_318), .S1(n80_adj_317));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_29.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_29.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_31 (.A0(n3047), .B0(n2273), .C0(n80_adj_381), 
          .D0(VCC_net), .A1(n3046), .B1(n2273), .C1(n77_adj_380), .D1(VCC_net), 
          .CIN(n11903), .COUT(n11904), .S0(n77_adj_316), .S1(n74_adj_315));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_31.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_31.INIT1 = 16'h1212;
    defparam _add_1_600_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_600_add_4_33 (.A0(n3045), .B0(n2273), .C0(n74_adj_379), 
          .D0(VCC_net), .A1(n71_adj_378), .B1(n2273), .C1(n68_adj_282), 
          .D1(n3044), .CIN(n11904), .S0(n71_adj_314), .S1(n3077));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_600_add_4_33.INIT0 = 16'h1212;
    defparam _add_1_600_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_600_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_600_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13007), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11906), .S1(n161_adj_567));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_582_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_3 (.A0(n161_adj_631), .B0(n13007), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_630), .B1(n13007), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11906), .COUT(n11907), .S0(n158_adj_566), 
          .S1(n155_adj_565));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_5 (.A0(n155_adj_629), .B0(n13007), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_628), .B1(n13007), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11907), .COUT(n11908), .S0(n152_adj_564), 
          .S1(n149_adj_563));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_7 (.A0(n149_adj_627), .B0(n13007), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_626), .B1(n13007), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11908), .COUT(n11909), .S0(n146_adj_562), 
          .S1(n143_adj_561));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_9 (.A0(n143_adj_625), .B0(n13007), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_624), .B1(n13007), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11909), .COUT(n11910), .S0(n140_adj_560), 
          .S1(n137_adj_559));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_11 (.A0(n137_adj_623), .B0(n13007), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_622), .B1(n13007), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11910), .COUT(n11911), .S0(n134_adj_558), 
          .S1(n131_adj_557));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_13 (.A0(n131_adj_621), .B0(n13007), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_620), .B1(n13007), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11911), .COUT(n11912), .S0(n128_adj_556), 
          .S1(n125_adj_555));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_15 (.A0(n125_adj_619), .B0(n13007), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_618), .B1(n13007), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11912), .COUT(n11913), .S0(n122_adj_554), 
          .S1(n119_adj_553));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_17 (.A0(n119_adj_617), .B0(n13007), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_616), .B1(n13007), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11913), .COUT(n11914), .S0(n116_adj_552), 
          .S1(n113_adj_551));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_19 (.A0(n113_adj_615), .B0(n13007), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_614), .B1(n13007), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11914), .COUT(n11915), .S0(n110_adj_550), 
          .S1(n107_adj_549));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_21 (.A0(n107_adj_613), .B0(n13007), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_612), .B1(n13007), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11915), .COUT(n11916), .S0(n104_adj_548), 
          .S1(n101_adj_547));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_23 (.A0(n101_adj_611), .B0(n13007), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_610), .B1(n13007), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11916), .COUT(n11917), .S0(n98_adj_546), 
          .S1(n95_adj_545));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_25 (.A0(n95_adj_609), .B0(n13007), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_608), .B1(n13007), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11917), .COUT(n11918), .S0(n92_adj_544), 
          .S1(n89_adj_543));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_27 (.A0(n89_adj_607), .B0(n13007), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_606), .B1(n13007), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11918), .COUT(n11919), .S0(n86_adj_542), 
          .S1(n83_adj_541));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_29 (.A0(n83_adj_605), .B0(n13007), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_604), .B1(n13007), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11919), .COUT(n11920), .S0(n80_adj_540), 
          .S1(n77_adj_539));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_31 (.A0(n77_adj_603), .B0(n13007), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_602), .B1(n13007), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11920), .COUT(n11921), .S0(n74_adj_538), 
          .S1(n71_adj_537));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_582_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_582_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_582_add_4_33 (.A0(n1067), .B0(n13007), .C0(n71_adj_601), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11921), .S0(n68_adj_536));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_582_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_582_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_582_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_582_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13008), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11922), .S1(n161_adj_599));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_579_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_3 (.A0(n161_adj_1680), .B0(n13008), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1679), .B1(n13008), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11922), .COUT(n11923), .S0(n158_adj_598), 
          .S1(n155_adj_597));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_5 (.A0(n155_adj_1678), .B0(n13008), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1677), .B1(n13008), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11923), .COUT(n11924), .S0(n152_adj_596), 
          .S1(n149_adj_595));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_7 (.A0(n149_adj_1676), .B0(n13008), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1675), .B1(n13008), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11924), .COUT(n11925), .S0(n146_adj_594), 
          .S1(n143_adj_593));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_9 (.A0(n143_adj_1674), .B0(n13008), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1673), .B1(n13008), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11925), .COUT(n11926), .S0(n140_adj_592), 
          .S1(n137_adj_591));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_11 (.A0(n137_adj_1672), .B0(n13008), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1671), .B1(n13008), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11926), .COUT(n11927), .S0(n134_adj_590), 
          .S1(n131_adj_589));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_13 (.A0(n131_adj_1670), .B0(n13008), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1669), .B1(n13008), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11927), .COUT(n11928), .S0(n128_adj_588), 
          .S1(n125_adj_587));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_15 (.A0(n125_adj_1668), .B0(n13008), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1667), .B1(n13008), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11928), .COUT(n11929), .S0(n122_adj_586), 
          .S1(n119_adj_585));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_17 (.A0(n119_adj_1666), .B0(n13008), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1665), .B1(n13008), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11929), .COUT(n11930), .S0(n116_adj_584), 
          .S1(n113_adj_583));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_19 (.A0(n113_adj_1664), .B0(n13008), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1663), .B1(n13008), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11930), .COUT(n11931), .S0(n110_adj_582), 
          .S1(n107_adj_581));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_21 (.A0(n107_adj_1662), .B0(n13008), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1661), .B1(n13008), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11931), .COUT(n11932), .S0(n104_adj_580), 
          .S1(n101_adj_579));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_23 (.A0(n101_adj_1660), .B0(n13008), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1659), .B1(n13008), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11932), .COUT(n11933), .S0(n98_adj_578), 
          .S1(n95_adj_577));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_25 (.A0(n95_adj_1658), .B0(n13008), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1657), .B1(n13008), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11933), .COUT(n11934), .S0(n92_adj_576), 
          .S1(n89_adj_575));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_27 (.A0(n89_adj_1656), .B0(n13008), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1655), .B1(n13008), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11934), .COUT(n11935), .S0(n86_adj_574), 
          .S1(n83_adj_573));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_29 (.A0(n83_adj_1654), .B0(n13008), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1653), .B1(n13008), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11935), .COUT(n11936), .S0(n80_adj_572), 
          .S1(n77_adj_571));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_31 (.A0(n77_adj_1652), .B0(n13008), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1651), .B1(n13008), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11936), .COUT(n11937), .S0(n74_adj_570), 
          .S1(n71_adj_569));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_579_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_579_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_579_add_4_33 (.A0(n1067), .B0(n13008), .C0(n71_adj_1650), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11937), .S0(n68_adj_568));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_579_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_579_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_579_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_579_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13008), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11938), .S1(n161_adj_631));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_576_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_3 (.A0(n161_adj_1712), .B0(n13008), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1711), .B1(n13008), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11938), .COUT(n11939), .S0(n158_adj_630), 
          .S1(n155_adj_629));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_5 (.A0(n155_adj_1710), .B0(n13008), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1709), .B1(n13008), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11939), .COUT(n11940), .S0(n152_adj_628), 
          .S1(n149_adj_627));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_7 (.A0(n149_adj_1708), .B0(n13008), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1707), .B1(n13008), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11940), .COUT(n11941), .S0(n146_adj_626), 
          .S1(n143_adj_625));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_9 (.A0(n143_adj_1706), .B0(n13008), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1705), .B1(n13008), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11941), .COUT(n11942), .S0(n140_adj_624), 
          .S1(n137_adj_623));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_11 (.A0(n137_adj_1704), .B0(n13008), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1703), .B1(n13008), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11942), .COUT(n11943), .S0(n134_adj_622), 
          .S1(n131_adj_621));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_13 (.A0(n131_adj_1702), .B0(n13008), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1701), .B1(n13008), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11943), .COUT(n11944), .S0(n128_adj_620), 
          .S1(n125_adj_619));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_15 (.A0(n125_adj_1700), .B0(n13008), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1699), .B1(n13008), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11944), .COUT(n11945), .S0(n122_adj_618), 
          .S1(n119_adj_617));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_17 (.A0(n119_adj_1698), .B0(n13008), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1697), .B1(n13008), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11945), .COUT(n11946), .S0(n116_adj_616), 
          .S1(n113_adj_615));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_19 (.A0(n113_adj_1696), .B0(n13008), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1695), .B1(n13008), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11946), .COUT(n11947), .S0(n110_adj_614), 
          .S1(n107_adj_613));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_21 (.A0(n107_adj_1694), .B0(n13008), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1693), .B1(n13008), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11947), .COUT(n11948), .S0(n104_adj_612), 
          .S1(n101_adj_611));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_23 (.A0(n101_adj_1692), .B0(n13008), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1691), .B1(n13008), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11948), .COUT(n11949), .S0(n98_adj_610), 
          .S1(n95_adj_609));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_25 (.A0(n95_adj_1690), .B0(n13008), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1689), .B1(n13008), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11949), .COUT(n11950), .S0(n92_adj_608), 
          .S1(n89_adj_607));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_27 (.A0(n89_adj_1688), .B0(n13008), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1687), .B1(n13008), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11950), .COUT(n11951), .S0(n86_adj_606), 
          .S1(n83_adj_605));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_29 (.A0(n83_adj_1686), .B0(n13008), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1685), .B1(n13008), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11951), .COUT(n11952), .S0(n80_adj_604), 
          .S1(n77_adj_603));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_31 (.A0(n77_adj_1684), .B0(n13008), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1683), .B1(n13008), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11952), .COUT(n11953), .S0(n74_adj_602), 
          .S1(n71_adj_601));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_576_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_576_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_576_add_4_33 (.A0(n1067), .B0(n13008), .C0(n71_adj_1682), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11953), .S0(n68_adj_600));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_576_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_576_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_576_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_576_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13013), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11954), .S1(n161_adj_663));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_549_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_3 (.A0(n161_adj_727), .B0(n13013), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_726), .B1(n13013), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11954), .COUT(n11955), .S0(n158_adj_662), 
          .S1(n155_adj_661));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_5 (.A0(n155_adj_725), .B0(n13013), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_724), .B1(n13013), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11955), .COUT(n11956), .S0(n152_adj_660), 
          .S1(n149_adj_659));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_7 (.A0(n149_adj_723), .B0(n13013), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_722), .B1(n13013), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11956), .COUT(n11957), .S0(n146_adj_658), 
          .S1(n143_adj_657));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_9 (.A0(n143_adj_721), .B0(n13013), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_720), .B1(n13013), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11957), .COUT(n11958), .S0(n140_adj_656), 
          .S1(n137_adj_655));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_11 (.A0(n137_adj_719), .B0(n13013), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_718), .B1(n13013), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11958), .COUT(n11959), .S0(n134_adj_654), 
          .S1(n131_adj_653));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_13 (.A0(n131_adj_717), .B0(n13013), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_716), .B1(n13013), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11959), .COUT(n11960), .S0(n128_adj_652), 
          .S1(n125_adj_651));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_15 (.A0(n125_adj_715), .B0(n13013), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_714), .B1(n13013), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11960), .COUT(n11961), .S0(n122_adj_650), 
          .S1(n119_adj_649));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_17 (.A0(n119_adj_713), .B0(n13013), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_712), .B1(n13013), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11961), .COUT(n11962), .S0(n116_adj_648), 
          .S1(n113_adj_647));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_19 (.A0(n113_adj_711), .B0(n13013), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_710), .B1(n13013), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11962), .COUT(n11963), .S0(n110_adj_646), 
          .S1(n107_adj_645));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_21 (.A0(n107_adj_709), .B0(n13013), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_708), .B1(n13013), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11963), .COUT(n11964), .S0(n104_adj_644), 
          .S1(n101_adj_643));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_23 (.A0(n101_adj_707), .B0(n13013), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_706), .B1(n13013), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11964), .COUT(n11965), .S0(n98_adj_642), 
          .S1(n95_adj_641));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_25 (.A0(n95_adj_705), .B0(n13013), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_704), .B1(n13013), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11965), .COUT(n11966), .S0(n92_adj_640), 
          .S1(n89_adj_639));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_27 (.A0(n89_adj_703), .B0(n13013), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_702), .B1(n13013), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11966), .COUT(n11967), .S0(n86_adj_638), 
          .S1(n83_adj_637));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_29 (.A0(n83_adj_701), .B0(n13013), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_700), .B1(n13013), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11967), .COUT(n11968), .S0(n80_adj_636), 
          .S1(n77_adj_635));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_31 (.A0(n77_adj_699), .B0(n13013), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_698), .B1(n13013), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11968), .COUT(n11969), .S0(n74_adj_634), 
          .S1(n71_adj_633));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_549_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_549_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_549_add_4_33 (.A0(n1067), .B0(n13013), .C0(n71_adj_697), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11969), .S0(n68_adj_632));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_549_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_549_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_549_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_549_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13013), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11970), .S1(n161_adj_695));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_546_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_3 (.A0(n161_adj_759), .B0(n13013), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_758), .B1(n13013), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11970), .COUT(n11971), .S0(n158_adj_694), 
          .S1(n155_adj_693));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_5 (.A0(n155_adj_757), .B0(n13013), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_756), .B1(n13013), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11971), .COUT(n11972), .S0(n152_adj_692), 
          .S1(n149_adj_691));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_7 (.A0(n149_adj_755), .B0(n13013), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_754), .B1(n13013), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11972), .COUT(n11973), .S0(n146_adj_690), 
          .S1(n143_adj_689));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_9 (.A0(n143_adj_753), .B0(n13013), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_752), .B1(n13013), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11973), .COUT(n11974), .S0(n140_adj_688), 
          .S1(n137_adj_687));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_11 (.A0(n137_adj_751), .B0(n13013), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_750), .B1(n13013), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11974), .COUT(n11975), .S0(n134_adj_686), 
          .S1(n131_adj_685));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_13 (.A0(n131_adj_749), .B0(n13013), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_748), .B1(n13013), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11975), .COUT(n11976), .S0(n128_adj_684), 
          .S1(n125_adj_683));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_15 (.A0(n125_adj_747), .B0(n13013), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_746), .B1(n13013), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11976), .COUT(n11977), .S0(n122_adj_682), 
          .S1(n119_adj_681));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_17 (.A0(n119_adj_745), .B0(n13013), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_744), .B1(n13013), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11977), .COUT(n11978), .S0(n116_adj_680), 
          .S1(n113_adj_679));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_19 (.A0(n113_adj_743), .B0(n13013), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_742), .B1(n13013), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11978), .COUT(n11979), .S0(n110_adj_678), 
          .S1(n107_adj_677));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_21 (.A0(n107_adj_741), .B0(n13013), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_740), .B1(n13013), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11979), .COUT(n11980), .S0(n104_adj_676), 
          .S1(n101_adj_675));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_23 (.A0(n101_adj_739), .B0(n13013), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_738), .B1(n13013), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11980), .COUT(n11981), .S0(n98_adj_674), 
          .S1(n95_adj_673));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_25 (.A0(n95_adj_737), .B0(n13013), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_736), .B1(n13013), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11981), .COUT(n11982), .S0(n92_adj_672), 
          .S1(n89_adj_671));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_27 (.A0(n89_adj_735), .B0(n13013), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_734), .B1(n13013), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11982), .COUT(n11983), .S0(n86_adj_670), 
          .S1(n83_adj_669));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_29 (.A0(n83_adj_733), .B0(n13013), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_732), .B1(n13013), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11983), .COUT(n11984), .S0(n80_adj_668), 
          .S1(n77_adj_667));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_31 (.A0(n77_adj_731), .B0(n13013), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_730), .B1(n13013), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n11984), .COUT(n11985), .S0(n74_adj_666), 
          .S1(n71_adj_665));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_546_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_546_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_546_add_4_33 (.A0(n1067), .B0(n13013), .C0(n71_adj_729), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11985), .S0(n68_adj_664));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_546_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_546_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_546_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_546_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13014), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n11986), .S1(n161_adj_727));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_543_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_3 (.A0(n161_adj_791), .B0(n13014), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_790), .B1(n13014), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n11986), .COUT(n11987), .S0(n158_adj_726), 
          .S1(n155_adj_725));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_5 (.A0(n155_adj_789), .B0(n13014), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_788), .B1(n13014), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n11987), .COUT(n11988), .S0(n152_adj_724), 
          .S1(n149_adj_723));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_7 (.A0(n149_adj_787), .B0(n13014), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_786), .B1(n13014), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n11988), .COUT(n11989), .S0(n146_adj_722), 
          .S1(n143_adj_721));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_9 (.A0(n143_adj_785), .B0(n13014), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_784), .B1(n13014), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n11989), .COUT(n11990), .S0(n140_adj_720), 
          .S1(n137_adj_719));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_11 (.A0(n137_adj_783), .B0(n13014), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_782), .B1(n13014), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n11990), .COUT(n11991), .S0(n134_adj_718), 
          .S1(n131_adj_717));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_13 (.A0(n131_adj_781), .B0(n13014), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_780), .B1(n13014), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n11991), .COUT(n11992), .S0(n128_adj_716), 
          .S1(n125_adj_715));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_15 (.A0(n125_adj_779), .B0(n13014), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_778), .B1(n13014), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n11992), .COUT(n11993), .S0(n122_adj_714), 
          .S1(n119_adj_713));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_17 (.A0(n119_adj_777), .B0(n13014), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_776), .B1(n13014), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n11993), .COUT(n11994), .S0(n116_adj_712), 
          .S1(n113_adj_711));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_19 (.A0(n113_adj_775), .B0(n13014), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_774), .B1(n13014), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n11994), .COUT(n11995), .S0(n110_adj_710), 
          .S1(n107_adj_709));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_21 (.A0(n107_adj_773), .B0(n13014), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_772), .B1(n13014), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n11995), .COUT(n11996), .S0(n104_adj_708), 
          .S1(n101_adj_707));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_23 (.A0(n101_adj_771), .B0(n13014), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_770), .B1(n13014), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n11996), .COUT(n11997), .S0(n98_adj_706), 
          .S1(n95_adj_705));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_25 (.A0(n95_adj_769), .B0(n13014), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_768), .B1(n13014), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n11997), .COUT(n11998), .S0(n92_adj_704), 
          .S1(n89_adj_703));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_27 (.A0(n89_adj_767), .B0(n13014), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_766), .B1(n13014), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n11998), .COUT(n11999), .S0(n86_adj_702), 
          .S1(n83_adj_701));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_29 (.A0(n83_adj_765), .B0(n13014), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_764), .B1(n13014), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n11999), .COUT(n12000), .S0(n80_adj_700), 
          .S1(n77_adj_699));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_31 (.A0(n77_adj_763), .B0(n13014), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_762), .B1(n13014), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12000), .COUT(n12001), .S0(n74_adj_698), 
          .S1(n71_adj_697));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_543_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_543_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_543_add_4_33 (.A0(n1067), .B0(n13014), .C0(n71_adj_761), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12001), .S0(n68_adj_696));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_543_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_543_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_543_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_543_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13014), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12002), .S1(n161_adj_759));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_540_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_3 (.A0(n161_adj_1174), .B0(n13014), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_822), .B1(n13014), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12002), .COUT(n12003), .S0(n158_adj_758), 
          .S1(n155_adj_757));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_5 (.A0(n155_adj_821), .B0(n13014), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_820), .B1(n13014), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12003), .COUT(n12004), .S0(n152_adj_756), 
          .S1(n149_adj_755));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_7 (.A0(n149_adj_819), .B0(n13014), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_818), .B1(n13014), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12004), .COUT(n12005), .S0(n146_adj_754), 
          .S1(n143_adj_753));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_9 (.A0(n143_adj_817), .B0(n13014), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_816), .B1(n13014), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12005), .COUT(n12006), .S0(n140_adj_752), 
          .S1(n137_adj_751));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_11 (.A0(n137_adj_815), .B0(n13014), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_814), .B1(n13014), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12006), .COUT(n12007), .S0(n134_adj_750), 
          .S1(n131_adj_749));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_13 (.A0(n131_adj_813), .B0(n13014), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_812), .B1(n13014), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12007), .COUT(n12008), .S0(n128_adj_748), 
          .S1(n125_adj_747));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_15 (.A0(n125_adj_811), .B0(n13014), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_810), .B1(n13014), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12008), .COUT(n12009), .S0(n122_adj_746), 
          .S1(n119_adj_745));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_17 (.A0(n119_adj_809), .B0(n13014), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_808), .B1(n13014), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12009), .COUT(n12010), .S0(n116_adj_744), 
          .S1(n113_adj_743));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_19 (.A0(n113_adj_807), .B0(n13014), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_806), .B1(n13014), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12010), .COUT(n12011), .S0(n110_adj_742), 
          .S1(n107_adj_741));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_21 (.A0(n107_adj_805), .B0(n13014), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_804), .B1(n13014), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12011), .COUT(n12012), .S0(n104_adj_740), 
          .S1(n101_adj_739));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_23 (.A0(n101_adj_803), .B0(n13014), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_802), .B1(n13014), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12012), .COUT(n12013), .S0(n98_adj_738), 
          .S1(n95_adj_737));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_25 (.A0(n95_adj_801), .B0(n13014), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_800), .B1(n13014), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12013), .COUT(n12014), .S0(n92_adj_736), 
          .S1(n89_adj_735));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_27 (.A0(n89_adj_799), .B0(n13014), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_798), .B1(n13014), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12014), .COUT(n12015), .S0(n86_adj_734), 
          .S1(n83_adj_733));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_29 (.A0(n83_adj_797), .B0(n13014), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_796), .B1(n13014), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12015), .COUT(n12016), .S0(n80_adj_732), 
          .S1(n77_adj_731));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_31 (.A0(n77_adj_795), .B0(n13014), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_794), .B1(n13014), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12016), .COUT(n12017), .S0(n74_adj_730), 
          .S1(n71_adj_729));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_540_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_540_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_540_add_4_33 (.A0(n1067), .B0(n13014), .C0(n71_adj_793), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12017), .S0(n68_adj_728));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_540_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_540_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_540_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_540_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_439), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12019), .S1(n158_adj_790));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_537_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_438), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_437), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12019), .COUT(n12020), .S0(n155_adj_789), 
          .S1(n152_adj_788));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_436), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_435), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12020), .COUT(n12021), .S0(n149_adj_787), 
          .S1(n146_adj_786));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_434), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_433), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12021), .COUT(n12022), .S0(n143_adj_785), 
          .S1(n140_adj_784));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_432), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_431), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12022), .COUT(n12023), .S0(n137_adj_783), 
          .S1(n134_adj_782));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_430), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_429), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12023), .COUT(n12024), .S0(n131_adj_781), 
          .S1(n128_adj_780));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_428), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_427), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12024), .COUT(n12025), .S0(n125_adj_779), 
          .S1(n122_adj_778));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_426), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_425), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12025), .COUT(n12026), .S0(n119_adj_777), 
          .S1(n116_adj_776));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_424), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_423), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12026), .COUT(n12027), .S0(n113_adj_775), 
          .S1(n110_adj_774));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_422), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_421), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12027), .COUT(n12028), .S0(n107_adj_773), 
          .S1(n104_adj_772));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_420), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_419), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12028), .COUT(n12029), .S0(n101_adj_771), 
          .S1(n98_adj_770));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_418), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_417), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12029), .COUT(n12030), .S0(n95_adj_769), 
          .S1(n92_adj_768));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_416), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_415), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12030), .COUT(n12031), .S0(n89_adj_767), 
          .S1(n86_adj_766));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_414), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_413), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12031), .COUT(n12032), .S0(n83_adj_765), 
          .S1(n80_adj_764));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_412), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_411), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12032), .COUT(n12033), .S0(n77_adj_763), 
          .S1(n74_adj_762));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_537_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_537_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_410), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_409), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12033), .S0(n71_adj_761), .S1(n68_adj_760));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_537_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_537_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_537_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_537_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_2 (.A0(n1098), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1097), .B1(n161_adj_439), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12036), .S1(n158_adj_822));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_534_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_4 (.A0(n1096), .B0(n158_adj_438), .C0(GND_net), 
          .D0(VCC_net), .A1(n1095), .B1(n155_adj_437), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12036), .COUT(n12037), .S0(n155_adj_821), 
          .S1(n152_adj_820));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_6 (.A0(n1094), .B0(n152_adj_436), .C0(GND_net), 
          .D0(VCC_net), .A1(n1093), .B1(n149_adj_435), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12037), .COUT(n12038), .S0(n149_adj_819), 
          .S1(n146_adj_818));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_8 (.A0(n1092), .B0(n146_adj_434), .C0(GND_net), 
          .D0(VCC_net), .A1(n1091), .B1(n143_adj_433), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12038), .COUT(n12039), .S0(n143_adj_817), 
          .S1(n140_adj_816));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_10 (.A0(n1090), .B0(n140_adj_432), .C0(GND_net), 
          .D0(VCC_net), .A1(n1089), .B1(n137_adj_431), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12039), .COUT(n12040), .S0(n137_adj_815), 
          .S1(n134_adj_814));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_12 (.A0(n1088), .B0(n134_adj_430), .C0(GND_net), 
          .D0(VCC_net), .A1(n1087), .B1(n131_adj_429), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12040), .COUT(n12041), .S0(n131_adj_813), 
          .S1(n128_adj_812));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_14 (.A0(n1086), .B0(n128_adj_428), .C0(GND_net), 
          .D0(VCC_net), .A1(n1085), .B1(n125_adj_427), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12041), .COUT(n12042), .S0(n125_adj_811), 
          .S1(n122_adj_810));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_16 (.A0(n1084), .B0(n122_adj_426), .C0(GND_net), 
          .D0(VCC_net), .A1(n1083), .B1(n119_adj_425), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12042), .COUT(n12043), .S0(n119_adj_809), 
          .S1(n116_adj_808));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_18 (.A0(n1082), .B0(n116_adj_424), .C0(GND_net), 
          .D0(VCC_net), .A1(n1081), .B1(n113_adj_423), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12043), .COUT(n12044), .S0(n113_adj_807), 
          .S1(n110_adj_806));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_20 (.A0(n1080), .B0(n110_adj_422), .C0(GND_net), 
          .D0(VCC_net), .A1(n1079), .B1(n107_adj_421), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12044), .COUT(n12045), .S0(n107_adj_805), 
          .S1(n104_adj_804));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_22 (.A0(n1078), .B0(n104_adj_420), .C0(GND_net), 
          .D0(VCC_net), .A1(n1077), .B1(n101_adj_419), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12045), .COUT(n12046), .S0(n101_adj_803), 
          .S1(n98_adj_802));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_24 (.A0(n1076), .B0(n98_adj_418), .C0(GND_net), 
          .D0(VCC_net), .A1(n1075), .B1(n95_adj_417), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12046), .COUT(n12047), .S0(n95_adj_801), 
          .S1(n92_adj_800));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_26 (.A0(n1074), .B0(n92_adj_416), .C0(GND_net), 
          .D0(VCC_net), .A1(n1073), .B1(n89_adj_415), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12047), .COUT(n12048), .S0(n89_adj_799), 
          .S1(n86_adj_798));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_28 (.A0(n1072), .B0(n86_adj_414), .C0(GND_net), 
          .D0(VCC_net), .A1(n1071), .B1(n83_adj_413), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12048), .COUT(n12049), .S0(n83_adj_797), 
          .S1(n80_adj_796));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_30 (.A0(n1070), .B0(n80_adj_412), .C0(GND_net), 
          .D0(VCC_net), .A1(n1069), .B1(n77_adj_411), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12049), .COUT(n12050), .S0(n77_adj_795), 
          .S1(n74_adj_794));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_534_add_4_32 (.A0(n1068), .B0(n74_adj_410), .C0(GND_net), 
          .D0(VCC_net), .A1(n1067), .B1(n71_adj_409), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12050), .S0(n71_adj_793), .S1(n68_adj_792));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_534_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_534_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_534_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_534_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n1033), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12055));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_531_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_531_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_3 (.A0(det_q4_28[0]), .B0(n1033), .C0(n161_adj_885), 
          .D0(n1534), .A1(n161_adj_917), .B1(n1033), .C1(n158_adj_884), 
          .D1(n1533), .CIN(n12055), .COUT(n12056), .S0(n161_adj_853), 
          .S1(n158_adj_852));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_3.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_3.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_5 (.A0(n158_adj_916), .B0(n1033), .C0(n155_adj_883), 
          .D0(n1532), .A1(n155_adj_915), .B1(n1033), .C1(n152_adj_882), 
          .D1(n1531), .CIN(n12056), .COUT(n12057), .S0(n155_adj_851), 
          .S1(n152_adj_850));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_5.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_5.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_7 (.A0(n152_adj_914), .B0(n1033), .C0(n149_adj_881), 
          .D0(n1530), .A1(n149_adj_913), .B1(n1033), .C1(n146_adj_880), 
          .D1(n1529), .CIN(n12057), .COUT(n12058), .S0(n149_adj_849), 
          .S1(n146_adj_848));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_7.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_7.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_9 (.A0(n146_adj_912), .B0(n1033), .C0(n143_adj_879), 
          .D0(n1528), .A1(n143_adj_911), .B1(n1033), .C1(n140_adj_878), 
          .D1(n1527), .CIN(n12058), .COUT(n12059), .S0(n143_adj_847), 
          .S1(n140_adj_846));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_9.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_9.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_11 (.A0(n140_adj_910), .B0(n1033), .C0(n137_adj_877), 
          .D0(n1526), .A1(n137_adj_909), .B1(n1033), .C1(n134_adj_876), 
          .D1(n1525), .CIN(n12059), .COUT(n12060), .S0(n137_adj_845), 
          .S1(n134_adj_844));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_11.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_11.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_13 (.A0(n134_adj_908), .B0(n1033), .C0(n131_adj_875), 
          .D0(n1524), .A1(n131_adj_907), .B1(n1033), .C1(n128_adj_874), 
          .D1(n1523), .CIN(n12060), .COUT(n12061), .S0(n131_adj_843), 
          .S1(n128_adj_842));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_13.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_13.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_15 (.A0(n128_adj_906), .B0(n1033), .C0(n125_adj_873), 
          .D0(n1522), .A1(n125_adj_905), .B1(n1033), .C1(n122_adj_872), 
          .D1(n1521), .CIN(n12061), .COUT(n12062), .S0(n125_adj_841), 
          .S1(n122_adj_840));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_15.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_15.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_17 (.A0(n122_adj_904), .B0(n1033), .C0(n119_adj_871), 
          .D0(n1520), .A1(n119_adj_903), .B1(n1033), .C1(n116_adj_870), 
          .D1(n1519), .CIN(n12062), .COUT(n12063), .S0(n119_adj_839), 
          .S1(n116_adj_838));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_17.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_17.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_19 (.A0(n116_adj_902), .B0(n1033), .C0(n113_adj_869), 
          .D0(n1518), .A1(n113_adj_901), .B1(n1033), .C1(n110_adj_868), 
          .D1(n1517), .CIN(n12063), .COUT(n12064), .S0(n113_adj_837), 
          .S1(n110_adj_836));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_19.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_19.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_21 (.A0(n110_adj_900), .B0(n1033), .C0(n107_adj_867), 
          .D0(n1516), .A1(n107_adj_899), .B1(n1033), .C1(n104_adj_866), 
          .D1(n1515), .CIN(n12064), .COUT(n12065), .S0(n107_adj_835), 
          .S1(n104_adj_834));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_21.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_21.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_23 (.A0(n104_adj_898), .B0(n1033), .C0(n101_adj_865), 
          .D0(n1514), .A1(n101_adj_897), .B1(n1033), .C1(n98_adj_864), 
          .D1(n1513), .CIN(n12065), .COUT(n12066), .S0(n101_adj_833), 
          .S1(n98_adj_832));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_23.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_23.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_25 (.A0(n98_adj_896), .B0(n1033), .C0(n95_adj_863), 
          .D0(n1512), .A1(n95_adj_895), .B1(n1033), .C1(n92_adj_862), 
          .D1(n1511), .CIN(n12066), .COUT(n12067), .S0(n95_adj_831), 
          .S1(n92_adj_830));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_25.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_25.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_27 (.A0(n92_adj_894), .B0(n1033), .C0(n89_adj_861), 
          .D0(n1510), .A1(n89_adj_893), .B1(n1033), .C1(n86_adj_860), 
          .D1(n1509), .CIN(n12067), .COUT(n12068), .S0(n89_adj_829), 
          .S1(n86_adj_828));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_27.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_27.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_29 (.A0(n86_adj_892), .B0(n1033), .C0(n83_adj_859), 
          .D0(n1508), .A1(n83_adj_891), .B1(n1033), .C1(n80_adj_858), 
          .D1(n1507), .CIN(n12068), .COUT(n12069), .S0(n83_adj_827), 
          .S1(n80_adj_826));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_29.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_29.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_31 (.A0(n80_adj_890), .B0(n1033), .C0(n77_adj_857), 
          .D0(n1506), .A1(n77_adj_889), .B1(n1033), .C1(n74_adj_856), 
          .D1(n1505), .CIN(n12069), .COUT(n12070), .S0(n77_adj_825), 
          .S1(n74_adj_824));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_31.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_31.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_531_add_4_33 (.A0(n74_adj_888), .B0(n1033), .C0(n71_adj_855), 
          .D0(n1504), .A1(n71_adj_887), .B1(n1033), .C1(n68_adj_854), 
          .D1(n1503), .CIN(n12070), .S0(n71_adj_823), .S1(n1536));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_531_add_4_33.INIT0 = 16'h74b8;
    defparam _add_1_531_add_4_33.INIT1 = 16'h74b8;
    defparam _add_1_531_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_531_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13023), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12072), .S1(n161_adj_885));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_528_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_3 (.A0(n161_adj_949), .B0(n13023), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_948), .B1(n13023), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12072), .COUT(n12073), .S0(n158_adj_884), 
          .S1(n155_adj_883));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_5 (.A0(n155_adj_947), .B0(n13023), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_946), .B1(n13023), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12073), .COUT(n12074), .S0(n152_adj_882), 
          .S1(n149_adj_881));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_7 (.A0(n149_adj_945), .B0(n13023), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_944), .B1(n13023), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12074), .COUT(n12075), .S0(n146_adj_880), 
          .S1(n143_adj_879));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_9 (.A0(n143_adj_943), .B0(n13023), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_942), .B1(n13023), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12075), .COUT(n12076), .S0(n140_adj_878), 
          .S1(n137_adj_877));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_11 (.A0(n137_adj_941), .B0(n13023), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_940), .B1(n13023), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12076), .COUT(n12077), .S0(n134_adj_876), 
          .S1(n131_adj_875));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_13 (.A0(n131_adj_939), .B0(n13023), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_938), .B1(n13023), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12077), .COUT(n12078), .S0(n128_adj_874), 
          .S1(n125_adj_873));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_15 (.A0(n125_adj_937), .B0(n13023), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_936), .B1(n13023), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12078), .COUT(n12079), .S0(n122_adj_872), 
          .S1(n119_adj_871));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_17 (.A0(n119_adj_935), .B0(n13023), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_934), .B1(n13023), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12079), .COUT(n12080), .S0(n116_adj_870), 
          .S1(n113_adj_869));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_19 (.A0(n113_adj_933), .B0(n13023), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_932), .B1(n13023), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12080), .COUT(n12081), .S0(n110_adj_868), 
          .S1(n107_adj_867));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_21 (.A0(n107_adj_931), .B0(n13023), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_930), .B1(n13023), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12081), .COUT(n12082), .S0(n104_adj_866), 
          .S1(n101_adj_865));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_23 (.A0(n101_adj_929), .B0(n13023), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_928), .B1(n13023), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12082), .COUT(n12083), .S0(n98_adj_864), 
          .S1(n95_adj_863));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_25 (.A0(n95_adj_927), .B0(n13023), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_926), .B1(n13023), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12083), .COUT(n12084), .S0(n92_adj_862), 
          .S1(n89_adj_861));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_27 (.A0(n89_adj_925), .B0(n13023), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_924), .B1(n13023), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12084), .COUT(n12085), .S0(n86_adj_860), 
          .S1(n83_adj_859));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_29 (.A0(n83_adj_923), .B0(n13023), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_922), .B1(n13023), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12085), .COUT(n12086), .S0(n80_adj_858), 
          .S1(n77_adj_857));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_31 (.A0(n77_adj_921), .B0(n13023), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_920), .B1(n13023), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12086), .COUT(n12087), .S0(n74_adj_856), 
          .S1(n71_adj_855));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_528_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_528_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_528_add_4_33 (.A0(n1067), .B0(n13023), .C0(n71_adj_919), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12087), .S0(n68_adj_854));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_528_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_528_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_528_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_528_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13024), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12088), .S1(n161_adj_917));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_525_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_3 (.A0(n161_adj_981), .B0(n13024), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_980), .B1(n13024), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12088), .COUT(n12089), .S0(n158_adj_916), 
          .S1(n155_adj_915));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_5 (.A0(n155_adj_979), .B0(n13024), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_978), .B1(n13024), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12089), .COUT(n12090), .S0(n152_adj_914), 
          .S1(n149_adj_913));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_7 (.A0(n149_adj_977), .B0(n13024), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_976), .B1(n13024), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12090), .COUT(n12091), .S0(n146_adj_912), 
          .S1(n143_adj_911));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_9 (.A0(n143_adj_975), .B0(n13024), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_974), .B1(n13024), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12091), .COUT(n12092), .S0(n140_adj_910), 
          .S1(n137_adj_909));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_11 (.A0(n137_adj_973), .B0(n13024), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_972), .B1(n13024), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12092), .COUT(n12093), .S0(n134_adj_908), 
          .S1(n131_adj_907));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_13 (.A0(n131_adj_971), .B0(n13024), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_970), .B1(n13024), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12093), .COUT(n12094), .S0(n128_adj_906), 
          .S1(n125_adj_905));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_15 (.A0(n125_adj_969), .B0(n13024), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_968), .B1(n13024), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12094), .COUT(n12095), .S0(n122_adj_904), 
          .S1(n119_adj_903));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_17 (.A0(n119_adj_967), .B0(n13024), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_966), .B1(n13024), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12095), .COUT(n12096), .S0(n116_adj_902), 
          .S1(n113_adj_901));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_19 (.A0(n113_adj_965), .B0(n13024), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_964), .B1(n13024), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12096), .COUT(n12097), .S0(n110_adj_900), 
          .S1(n107_adj_899));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_21 (.A0(n107_adj_963), .B0(n13024), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_962), .B1(n13024), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12097), .COUT(n12098), .S0(n104_adj_898), 
          .S1(n101_adj_897));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_23 (.A0(n101_adj_961), .B0(n13024), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_960), .B1(n13024), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12098), .COUT(n12099), .S0(n98_adj_896), 
          .S1(n95_adj_895));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_25 (.A0(n95_adj_959), .B0(n13024), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_958), .B1(n13024), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12099), .COUT(n12100), .S0(n92_adj_894), 
          .S1(n89_adj_893));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_27 (.A0(n89_adj_957), .B0(n13024), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_956), .B1(n13024), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12100), .COUT(n12101), .S0(n86_adj_892), 
          .S1(n83_adj_891));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_29 (.A0(n83_adj_955), .B0(n13024), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_954), .B1(n13024), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12101), .COUT(n12102), .S0(n80_adj_890), 
          .S1(n77_adj_889));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_31 (.A0(n77_adj_953), .B0(n13024), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_952), .B1(n13024), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12102), .COUT(n12103), .S0(n74_adj_888), 
          .S1(n71_adj_887));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_525_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_525_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_525_add_4_33 (.A0(n1067), .B0(n13024), .C0(n71_adj_951), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12103), .S0(n68_adj_886));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_525_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_525_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_525_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_525_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13024), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12104), .S1(n161_adj_949));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_522_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_3 (.A0(n161_adj_1013), .B0(n13024), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1012), .B1(n13024), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12104), .COUT(n12105), .S0(n158_adj_948), 
          .S1(n155_adj_947));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_5 (.A0(n155_adj_1011), .B0(n13024), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1010), .B1(n13024), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12105), .COUT(n12106), .S0(n152_adj_946), 
          .S1(n149_adj_945));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_7 (.A0(n149_adj_1009), .B0(n13024), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1008), .B1(n13024), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12106), .COUT(n12107), .S0(n146_adj_944), 
          .S1(n143_adj_943));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_9 (.A0(n143_adj_1007), .B0(n13024), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1006), .B1(n13024), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12107), .COUT(n12108), .S0(n140_adj_942), 
          .S1(n137_adj_941));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_11 (.A0(n137_adj_1005), .B0(n13024), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1004), .B1(n13024), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12108), .COUT(n12109), .S0(n134_adj_940), 
          .S1(n131_adj_939));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_13 (.A0(n131_adj_1003), .B0(n13024), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1002), .B1(n13024), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12109), .COUT(n12110), .S0(n128_adj_938), 
          .S1(n125_adj_937));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_15 (.A0(n125_adj_1001), .B0(n13024), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1000), .B1(n13024), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12110), .COUT(n12111), .S0(n122_adj_936), 
          .S1(n119_adj_935));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_17 (.A0(n119_adj_999), .B0(n13024), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_998), .B1(n13024), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12111), .COUT(n12112), .S0(n116_adj_934), 
          .S1(n113_adj_933));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_19 (.A0(n113_adj_997), .B0(n13024), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_996), .B1(n13024), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12112), .COUT(n12113), .S0(n110_adj_932), 
          .S1(n107_adj_931));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_21 (.A0(n107_adj_995), .B0(n13024), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_994), .B1(n13024), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12113), .COUT(n12114), .S0(n104_adj_930), 
          .S1(n101_adj_929));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_23 (.A0(n101_adj_993), .B0(n13024), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_992), .B1(n13024), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12114), .COUT(n12115), .S0(n98_adj_928), 
          .S1(n95_adj_927));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_25 (.A0(n95_adj_991), .B0(n13024), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_990), .B1(n13024), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12115), .COUT(n12116), .S0(n92_adj_926), 
          .S1(n89_adj_925));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_27 (.A0(n89_adj_989), .B0(n13024), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_988), .B1(n13024), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12116), .COUT(n12117), .S0(n86_adj_924), 
          .S1(n83_adj_923));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_29 (.A0(n83_adj_987), .B0(n13024), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_986), .B1(n13024), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12117), .COUT(n12118), .S0(n80_adj_922), 
          .S1(n77_adj_921));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_31 (.A0(n77_adj_985), .B0(n13024), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_984), .B1(n13024), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12118), .COUT(n12119), .S0(n74_adj_920), 
          .S1(n71_adj_919));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_522_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_522_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_522_add_4_33 (.A0(n1067), .B0(n13024), .C0(n71_adj_983), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12119), .S0(n68_adj_918));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_522_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_522_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_522_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_522_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13025), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12120), .S1(n161_adj_981));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_519_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_3 (.A0(n161_adj_1045), .B0(n13025), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1044), .B1(n13025), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12120), .COUT(n12121), .S0(n158_adj_980), 
          .S1(n155_adj_979));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_5 (.A0(n155_adj_1043), .B0(n13025), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1042), .B1(n13025), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12121), .COUT(n12122), .S0(n152_adj_978), 
          .S1(n149_adj_977));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_7 (.A0(n149_adj_1041), .B0(n13025), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1040), .B1(n13025), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12122), .COUT(n12123), .S0(n146_adj_976), 
          .S1(n143_adj_975));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_9 (.A0(n143_adj_1039), .B0(n13025), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1038), .B1(n13025), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12123), .COUT(n12124), .S0(n140_adj_974), 
          .S1(n137_adj_973));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_11 (.A0(n137_adj_1037), .B0(n13025), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1036), .B1(n13025), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12124), .COUT(n12125), .S0(n134_adj_972), 
          .S1(n131_adj_971));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_13 (.A0(n131_adj_1035), .B0(n13025), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1034), .B1(n13025), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12125), .COUT(n12126), .S0(n128_adj_970), 
          .S1(n125_adj_969));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_15 (.A0(n125_adj_1033), .B0(n13025), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1032), .B1(n13025), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12126), .COUT(n12127), .S0(n122_adj_968), 
          .S1(n119_adj_967));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_17 (.A0(n119_adj_1031), .B0(n13025), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1030), .B1(n13025), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12127), .COUT(n12128), .S0(n116_adj_966), 
          .S1(n113_adj_965));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_19 (.A0(n113_adj_1029), .B0(n13025), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1028), .B1(n13025), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12128), .COUT(n12129), .S0(n110_adj_964), 
          .S1(n107_adj_963));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_21 (.A0(n107_adj_1027), .B0(n13025), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1026), .B1(n13025), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12129), .COUT(n12130), .S0(n104_adj_962), 
          .S1(n101_adj_961));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_23 (.A0(n101_adj_1025), .B0(n13025), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1024), .B1(n13025), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12130), .COUT(n12131), .S0(n98_adj_960), 
          .S1(n95_adj_959));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_25 (.A0(n95_adj_1023), .B0(n13025), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1022), .B1(n13025), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12131), .COUT(n12132), .S0(n92_adj_958), 
          .S1(n89_adj_957));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_27 (.A0(n89_adj_1021), .B0(n13025), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1020), .B1(n13025), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12132), .COUT(n12133), .S0(n86_adj_956), 
          .S1(n83_adj_955));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_29 (.A0(n83_adj_1019), .B0(n13025), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1018), .B1(n13025), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12133), .COUT(n12134), .S0(n80_adj_954), 
          .S1(n77_adj_953));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_31 (.A0(n77_adj_1017), .B0(n13025), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1016), .B1(n13025), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12134), .COUT(n12135), .S0(n74_adj_952), 
          .S1(n71_adj_951));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_519_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_519_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_519_add_4_33 (.A0(n1067), .B0(n13025), .C0(n71_adj_1015), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12135), .S0(n68_adj_950));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_519_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_519_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_519_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_519_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13025), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12136), .S1(n161_adj_1013));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_516_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_3 (.A0(n161_adj_1077), .B0(n13025), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1076), .B1(n13025), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12136), .COUT(n12137), .S0(n158_adj_1012), 
          .S1(n155_adj_1011));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_5 (.A0(n155_adj_1075), .B0(n13025), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1074), .B1(n13025), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12137), .COUT(n12138), .S0(n152_adj_1010), 
          .S1(n149_adj_1009));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_7 (.A0(n149_adj_1073), .B0(n13025), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1072), .B1(n13025), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12138), .COUT(n12139), .S0(n146_adj_1008), 
          .S1(n143_adj_1007));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_9 (.A0(n143_adj_1071), .B0(n13025), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1070), .B1(n13025), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12139), .COUT(n12140), .S0(n140_adj_1006), 
          .S1(n137_adj_1005));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_11 (.A0(n137_adj_1069), .B0(n13025), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1068), .B1(n13025), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12140), .COUT(n12141), .S0(n134_adj_1004), 
          .S1(n131_adj_1003));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_13 (.A0(n131_adj_1067), .B0(n13025), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1066), .B1(n13025), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12141), .COUT(n12142), .S0(n128_adj_1002), 
          .S1(n125_adj_1001));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_15 (.A0(n125_adj_1065), .B0(n13025), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1064), .B1(n13025), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12142), .COUT(n12143), .S0(n122_adj_1000), 
          .S1(n119_adj_999));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_17 (.A0(n119_adj_1063), .B0(n13025), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1062), .B1(n13025), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12143), .COUT(n12144), .S0(n116_adj_998), 
          .S1(n113_adj_997));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_19 (.A0(n113_adj_1061), .B0(n13025), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1060), .B1(n13025), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12144), .COUT(n12145), .S0(n110_adj_996), 
          .S1(n107_adj_995));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_21 (.A0(n107_adj_1059), .B0(n13025), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1058), .B1(n13025), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12145), .COUT(n12146), .S0(n104_adj_994), 
          .S1(n101_adj_993));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_23 (.A0(n101_adj_1057), .B0(n13025), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1056), .B1(n13025), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12146), .COUT(n12147), .S0(n98_adj_992), 
          .S1(n95_adj_991));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_25 (.A0(n95_adj_1055), .B0(n13025), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1054), .B1(n13025), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12147), .COUT(n12148), .S0(n92_adj_990), 
          .S1(n89_adj_989));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_27 (.A0(n89_adj_1053), .B0(n13025), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1052), .B1(n13025), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12148), .COUT(n12149), .S0(n86_adj_988), 
          .S1(n83_adj_987));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_29 (.A0(n83_adj_1051), .B0(n13025), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1050), .B1(n13025), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12149), .COUT(n12150), .S0(n80_adj_986), 
          .S1(n77_adj_985));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_31 (.A0(n77_adj_1049), .B0(n13025), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1048), .B1(n13025), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12150), .COUT(n12151), .S0(n74_adj_984), 
          .S1(n71_adj_983));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_516_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_516_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_516_add_4_33 (.A0(n1067), .B0(n13025), .C0(n71_adj_1047), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12151), .S0(n68_adj_982));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_516_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_516_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_516_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_516_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13026), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12152), .S1(n161_adj_1045));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_513_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_3 (.A0(n161_adj_1109), .B0(n13026), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1108), .B1(n13026), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12152), .COUT(n12153), .S0(n158_adj_1044), 
          .S1(n155_adj_1043));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_5 (.A0(n155_adj_1107), .B0(n13026), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1106), .B1(n13026), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12153), .COUT(n12154), .S0(n152_adj_1042), 
          .S1(n149_adj_1041));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_7 (.A0(n149_adj_1105), .B0(n13026), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1104), .B1(n13026), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12154), .COUT(n12155), .S0(n146_adj_1040), 
          .S1(n143_adj_1039));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_9 (.A0(n143_adj_1103), .B0(n13026), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1102), .B1(n13026), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12155), .COUT(n12156), .S0(n140_adj_1038), 
          .S1(n137_adj_1037));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_11 (.A0(n137_adj_1101), .B0(n13026), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1100), .B1(n13026), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12156), .COUT(n12157), .S0(n134_adj_1036), 
          .S1(n131_adj_1035));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_13 (.A0(n131_adj_1099), .B0(n13026), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1098), .B1(n13026), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12157), .COUT(n12158), .S0(n128_adj_1034), 
          .S1(n125_adj_1033));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_15 (.A0(n125_adj_1097), .B0(n13026), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1096), .B1(n13026), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12158), .COUT(n12159), .S0(n122_adj_1032), 
          .S1(n119_adj_1031));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_17 (.A0(n119_adj_1095), .B0(n13026), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1094), .B1(n13026), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12159), .COUT(n12160), .S0(n116_adj_1030), 
          .S1(n113_adj_1029));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_19 (.A0(n113_adj_1093), .B0(n13026), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1092), .B1(n13026), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12160), .COUT(n12161), .S0(n110_adj_1028), 
          .S1(n107_adj_1027));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_21 (.A0(n107_adj_1091), .B0(n13026), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1090), .B1(n13026), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12161), .COUT(n12162), .S0(n104_adj_1026), 
          .S1(n101_adj_1025));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_23 (.A0(n101_adj_1089), .B0(n13026), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1088), .B1(n13026), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12162), .COUT(n12163), .S0(n98_adj_1024), 
          .S1(n95_adj_1023));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_25 (.A0(n95_adj_1087), .B0(n13026), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1086), .B1(n13026), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12163), .COUT(n12164), .S0(n92_adj_1022), 
          .S1(n89_adj_1021));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_27 (.A0(n89_adj_1085), .B0(n13026), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1084), .B1(n13026), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12164), .COUT(n12165), .S0(n86_adj_1020), 
          .S1(n83_adj_1019));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_29 (.A0(n83_adj_1083), .B0(n13026), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1082), .B1(n13026), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12165), .COUT(n12166), .S0(n80_adj_1018), 
          .S1(n77_adj_1017));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_31 (.A0(n77_adj_1081), .B0(n13026), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1080), .B1(n13026), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12166), .COUT(n12167), .S0(n74_adj_1016), 
          .S1(n71_adj_1015));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_513_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_513_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_513_add_4_33 (.A0(n1067), .B0(n13026), .C0(n71_adj_1079), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12167), .S0(n68_adj_1014));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_513_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_513_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_513_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_513_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13026), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12168), .S1(n161_adj_1077));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_510_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_3 (.A0(n161_adj_1141), .B0(n13026), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1140), .B1(n13026), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12168), .COUT(n12169), .S0(n158_adj_1076), 
          .S1(n155_adj_1075));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_5 (.A0(n155_adj_1139), .B0(n13026), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1138), .B1(n13026), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12169), .COUT(n12170), .S0(n152_adj_1074), 
          .S1(n149_adj_1073));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_7 (.A0(n149_adj_1137), .B0(n13026), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1136), .B1(n13026), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12170), .COUT(n12171), .S0(n146_adj_1072), 
          .S1(n143_adj_1071));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_9 (.A0(n143_adj_1135), .B0(n13026), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1134), .B1(n13026), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12171), .COUT(n12172), .S0(n140_adj_1070), 
          .S1(n137_adj_1069));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_11 (.A0(n137_adj_1133), .B0(n13026), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1132), .B1(n13026), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12172), .COUT(n12173), .S0(n134_adj_1068), 
          .S1(n131_adj_1067));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_13 (.A0(n131_adj_1131), .B0(n13026), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1130), .B1(n13026), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12173), .COUT(n12174), .S0(n128_adj_1066), 
          .S1(n125_adj_1065));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_15 (.A0(n125_adj_1129), .B0(n13026), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1128), .B1(n13026), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12174), .COUT(n12175), .S0(n122_adj_1064), 
          .S1(n119_adj_1063));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_17 (.A0(n119_adj_1127), .B0(n13026), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1126), .B1(n13026), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12175), .COUT(n12176), .S0(n116_adj_1062), 
          .S1(n113_adj_1061));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_19 (.A0(n113_adj_1125), .B0(n13026), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1124), .B1(n13026), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12176), .COUT(n12177), .S0(n110_adj_1060), 
          .S1(n107_adj_1059));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_21 (.A0(n107_adj_1123), .B0(n13026), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1122), .B1(n13026), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12177), .COUT(n12178), .S0(n104_adj_1058), 
          .S1(n101_adj_1057));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_23 (.A0(n101_adj_1121), .B0(n13026), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1120), .B1(n13026), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12178), .COUT(n12179), .S0(n98_adj_1056), 
          .S1(n95_adj_1055));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_25 (.A0(n95_adj_1119), .B0(n13026), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1118), .B1(n13026), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12179), .COUT(n12180), .S0(n92_adj_1054), 
          .S1(n89_adj_1053));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_27 (.A0(n89_adj_1117), .B0(n13026), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1116), .B1(n13026), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12180), .COUT(n12181), .S0(n86_adj_1052), 
          .S1(n83_adj_1051));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_29 (.A0(n83_adj_1115), .B0(n13026), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1114), .B1(n13026), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12181), .COUT(n12182), .S0(n80_adj_1050), 
          .S1(n77_adj_1049));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_31 (.A0(n77_adj_1113), .B0(n13026), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1112), .B1(n13026), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12182), .COUT(n12183), .S0(n74_adj_1048), 
          .S1(n71_adj_1047));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_510_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_510_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_510_add_4_33 (.A0(n1067), .B0(n13026), .C0(n71_adj_1111), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12183), .S0(n68_adj_1046));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_510_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_510_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_510_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_510_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12184), .S1(c_s[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_420_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_420_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_3 (.A0(c_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12184), .COUT(n12185), .S0(c_s[1]), .S1(c_s[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_5 (.A0(c_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12185), .COUT(n12186), .S0(c_s[3]), .S1(c_s[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_7 (.A0(c_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12186), .COUT(n12187), .S0(c_s[5]), .S1(c_s[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_9 (.A0(c_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12187), .COUT(n12188), .S0(c_s[7]), .S1(c_s[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_11 (.A0(c_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12188), .COUT(n12189), .S0(c_s[9]), .S1(c_s[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_13 (.A0(c_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12189), .COUT(n12190), .S0(c_s[11]), .S1(c_s[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_13.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_15 (.A0(c_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12190), .COUT(n12191), .S0(c_s[13]), .S1(c_s[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_15.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_15.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_420_add_4_17 (.A0(c_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(c_reg[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12191), .S0(c_s[15]), .S1(c_s[16]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(80[30:58])
    defparam _add_1_420_add_4_17.INIT0 = 16'h5555;
    defparam _add_1_420_add_4_17.INIT1 = 16'h5555;
    defparam _add_1_420_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_420_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13027), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12193), .S1(n161_adj_1109));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_507_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_3 (.A0(n161_adj_1585), .B0(n13027), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1584), .B1(n13027), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12193), .COUT(n12194), .S0(n158_adj_1108), 
          .S1(n155_adj_1107));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_5 (.A0(n155_adj_1583), .B0(n13027), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1582), .B1(n13027), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12194), .COUT(n12195), .S0(n152_adj_1106), 
          .S1(n149_adj_1105));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_7 (.A0(n149_adj_1581), .B0(n13027), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1580), .B1(n13027), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12195), .COUT(n12196), .S0(n146_adj_1104), 
          .S1(n143_adj_1103));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_9 (.A0(n143_adj_1579), .B0(n13027), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1578), .B1(n13027), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12196), .COUT(n12197), .S0(n140_adj_1102), 
          .S1(n137_adj_1101));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_11 (.A0(n137_adj_1577), .B0(n13027), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1576), .B1(n13027), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12197), .COUT(n12198), .S0(n134_adj_1100), 
          .S1(n131_adj_1099));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_13 (.A0(n131_adj_1575), .B0(n13027), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1574), .B1(n13027), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12198), .COUT(n12199), .S0(n128_adj_1098), 
          .S1(n125_adj_1097));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_15 (.A0(n125_adj_1573), .B0(n13027), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1572), .B1(n13027), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12199), .COUT(n12200), .S0(n122_adj_1096), 
          .S1(n119_adj_1095));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_17 (.A0(n119_adj_1571), .B0(n13027), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1570), .B1(n13027), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12200), .COUT(n12201), .S0(n116_adj_1094), 
          .S1(n113_adj_1093));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_19 (.A0(n113_adj_1569), .B0(n13027), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1568), .B1(n13027), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12201), .COUT(n12202), .S0(n110_adj_1092), 
          .S1(n107_adj_1091));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_21 (.A0(n107_adj_1567), .B0(n13027), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1566), .B1(n13027), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12202), .COUT(n12203), .S0(n104_adj_1090), 
          .S1(n101_adj_1089));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_23 (.A0(n101_adj_1565), .B0(n13027), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1564), .B1(n13027), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12203), .COUT(n12204), .S0(n98_adj_1088), 
          .S1(n95_adj_1087));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_25 (.A0(n95_adj_1563), .B0(n13027), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1562), .B1(n13027), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12204), .COUT(n12205), .S0(n92_adj_1086), 
          .S1(n89_adj_1085));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_27 (.A0(n89_adj_1561), .B0(n13027), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1560), .B1(n13027), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12205), .COUT(n12206), .S0(n86_adj_1084), 
          .S1(n83_adj_1083));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_29 (.A0(n83_adj_1559), .B0(n13027), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1558), .B1(n13027), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12206), .COUT(n12207), .S0(n80_adj_1082), 
          .S1(n77_adj_1081));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_31 (.A0(n77_adj_1557), .B0(n13027), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1556), .B1(n13027), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12207), .COUT(n12208), .S0(n74_adj_1080), 
          .S1(n71_adj_1079));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_507_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_507_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_507_add_4_33 (.A0(n1067), .B0(n13027), .C0(n71_adj_1555), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12208), .S0(n68_adj_1078));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_507_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_507_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_507_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_507_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13027), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12209), .S1(n161_adj_1141));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_504_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_3 (.A0(n161_adj_1744), .B0(n13027), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1743), .B1(n13027), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12209), .COUT(n12210), .S0(n158_adj_1140), 
          .S1(n155_adj_1139));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_5 (.A0(n155_adj_1742), .B0(n13027), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1741), .B1(n13027), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12210), .COUT(n12211), .S0(n152_adj_1138), 
          .S1(n149_adj_1137));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_7 (.A0(n149_adj_1740), .B0(n13027), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1739), .B1(n13027), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12211), .COUT(n12212), .S0(n146_adj_1136), 
          .S1(n143_adj_1135));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_9 (.A0(n143_adj_1738), .B0(n13027), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1737), .B1(n13027), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12212), .COUT(n12213), .S0(n140_adj_1134), 
          .S1(n137_adj_1133));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_11 (.A0(n137_adj_1736), .B0(n13027), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1735), .B1(n13027), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12213), .COUT(n12214), .S0(n134_adj_1132), 
          .S1(n131_adj_1131));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_13 (.A0(n131_adj_1734), .B0(n13027), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1733), .B1(n13027), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12214), .COUT(n12215), .S0(n128_adj_1130), 
          .S1(n125_adj_1129));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_15 (.A0(n125_adj_1732), .B0(n13027), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1731), .B1(n13027), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12215), .COUT(n12216), .S0(n122_adj_1128), 
          .S1(n119_adj_1127));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_17 (.A0(n119_adj_1730), .B0(n13027), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1729), .B1(n13027), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12216), .COUT(n12217), .S0(n116_adj_1126), 
          .S1(n113_adj_1125));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_19 (.A0(n113_adj_1728), .B0(n13027), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1727), .B1(n13027), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12217), .COUT(n12218), .S0(n110_adj_1124), 
          .S1(n107_adj_1123));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_21 (.A0(n107_adj_1726), .B0(n13027), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1725), .B1(n13027), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12218), .COUT(n12219), .S0(n104_adj_1122), 
          .S1(n101_adj_1121));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_23 (.A0(n101_adj_1724), .B0(n13027), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1723), .B1(n13027), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12219), .COUT(n12220), .S0(n98_adj_1120), 
          .S1(n95_adj_1119));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_25 (.A0(n95_adj_1722), .B0(n13027), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1721), .B1(n13027), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12220), .COUT(n12221), .S0(n92_adj_1118), 
          .S1(n89_adj_1117));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_27 (.A0(n89_adj_1720), .B0(n13027), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1719), .B1(n13027), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12221), .COUT(n12222), .S0(n86_adj_1116), 
          .S1(n83_adj_1115));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_29 (.A0(n83_adj_1718), .B0(n13027), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1717), .B1(n13027), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12222), .COUT(n12223), .S0(n80_adj_1114), 
          .S1(n77_adj_1113));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_31 (.A0(n77_adj_1716), .B0(n13027), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1715), .B1(n13027), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12223), .COUT(n12224), .S0(n74_adj_1112), 
          .S1(n71_adj_1111));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_504_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_504_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_504_add_4_33 (.A0(n1067), .B0(n13027), .C0(n71_adj_1714), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12224), .S0(n68_adj_1110));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_504_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_504_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_504_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_504_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_281), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12225));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_486_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_280), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_279), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12225), .COUT(n12226));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_278), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_277), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12226), .COUT(n12227));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_276), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_275), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12227), .COUT(n12228));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_274), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_273), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12228), .COUT(n12229));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_272), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_271), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12229), .COUT(n12230));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_270), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_269), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12230), .COUT(n12231));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_268), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_267), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12231), .COUT(n12232));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_266), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_265), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12232), .COUT(n12233));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_264), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_263), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12233), .COUT(n12234));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_262), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_261), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12234), .COUT(n12235));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_260), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_259), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12235), .COUT(n12236));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_258), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_257), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12236), .COUT(n12237));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_256), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_255), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12237), .COUT(n12238));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_254), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_253), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12238), .COUT(n12239));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_486_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_486_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_252), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_251), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12239), .S1(n68_adj_1142));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_486_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_486_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_486_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_486_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_2 (.A0(n1098), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1097), .B1(n161_adj_1236), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12242), .S1(n158_adj_1173));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_483_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_4 (.A0(n1096), .B0(n158_adj_1235), .C0(GND_net), 
          .D0(VCC_net), .A1(n1095), .B1(n155_adj_1234), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12242), .COUT(n12243), .S0(n155_adj_1172), 
          .S1(n152_adj_1171));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_6 (.A0(n1094), .B0(n152_adj_1233), .C0(GND_net), 
          .D0(VCC_net), .A1(n1093), .B1(n149_adj_1232), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12243), .COUT(n12244), .S0(n149_adj_1170), 
          .S1(n146_adj_1169));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_8 (.A0(n1092), .B0(n146_adj_1231), .C0(GND_net), 
          .D0(VCC_net), .A1(n1091), .B1(n143_adj_1230), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12244), .COUT(n12245), .S0(n143_adj_1168), 
          .S1(n140_adj_1167));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_10 (.A0(n1090), .B0(n140_adj_1229), .C0(GND_net), 
          .D0(VCC_net), .A1(n1089), .B1(n137_adj_1228), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12245), .COUT(n12246), .S0(n137_adj_1166), 
          .S1(n134_adj_1165));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_12 (.A0(n1088), .B0(n134_adj_1227), .C0(GND_net), 
          .D0(VCC_net), .A1(n1087), .B1(n131_adj_1226), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12246), .COUT(n12247), .S0(n131_adj_1164), 
          .S1(n128_adj_1163));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_14 (.A0(n1086), .B0(n128_adj_1225), .C0(GND_net), 
          .D0(VCC_net), .A1(n1085), .B1(n125_adj_1224), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12247), .COUT(n12248), .S0(n125_adj_1162), 
          .S1(n122_adj_1161));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_16 (.A0(n1084), .B0(n122_adj_1223), .C0(GND_net), 
          .D0(VCC_net), .A1(n1083), .B1(n119_adj_1222), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12248), .COUT(n12249), .S0(n119_adj_1160), 
          .S1(n116_adj_1159));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_18 (.A0(n1082), .B0(n116_adj_1221), .C0(GND_net), 
          .D0(VCC_net), .A1(n1081), .B1(n113_adj_1220), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12249), .COUT(n12250), .S0(n113_adj_1158), 
          .S1(n110_adj_1157));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_20 (.A0(n1080), .B0(n110_adj_1219), .C0(GND_net), 
          .D0(VCC_net), .A1(n1079), .B1(n107_adj_1218), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12250), .COUT(n12251), .S0(n107_adj_1156), 
          .S1(n104_adj_1155));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_22 (.A0(n1078), .B0(n104_adj_1217), .C0(GND_net), 
          .D0(VCC_net), .A1(n1077), .B1(n101_adj_1216), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12251), .COUT(n12252), .S0(n101_adj_1154), 
          .S1(n98_adj_1153));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_24 (.A0(n1076), .B0(n98_adj_1215), .C0(GND_net), 
          .D0(VCC_net), .A1(n1075), .B1(n95_adj_1214), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12252), .COUT(n12253), .S0(n95_adj_1152), 
          .S1(n92_adj_1151));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_26 (.A0(n1074), .B0(n92_adj_1213), .C0(GND_net), 
          .D0(VCC_net), .A1(n1073), .B1(n89_adj_1212), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12253), .COUT(n12254), .S0(n89_adj_1150), 
          .S1(n86_adj_1149));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_28 (.A0(n1072), .B0(n86_adj_1211), .C0(GND_net), 
          .D0(VCC_net), .A1(n1071), .B1(n83_adj_1210), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12254), .COUT(n12255), .S0(n83_adj_1148), 
          .S1(n80_adj_1147));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_30 (.A0(n1070), .B0(n80_adj_1209), .C0(GND_net), 
          .D0(VCC_net), .A1(n1069), .B1(n77_adj_1208), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12255), .COUT(n12256), .S0(n77_adj_1146), 
          .S1(n74_adj_1145));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_483_add_4_32 (.A0(n1068), .B0(n74_adj_1207), .C0(GND_net), 
          .D0(VCC_net), .A1(n1067), .B1(n71_adj_1206), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12256), .S0(n71_adj_1144), .S1(n68_adj_1143));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_483_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_483_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_483_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_483_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_1236), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12259), .S1(n158_adj_1205));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_480_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_1235), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_1234), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12259), .COUT(n12260), .S0(n155_adj_1204), 
          .S1(n152_adj_1203));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_1233), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_1232), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12260), .COUT(n12261), .S0(n149_adj_1202), 
          .S1(n146_adj_1201));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_1231), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_1230), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12261), .COUT(n12262), .S0(n143_adj_1200), 
          .S1(n140_adj_1199));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_1229), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_1228), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12262), .COUT(n12263), .S0(n137_adj_1198), 
          .S1(n134_adj_1197));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_1227), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_1226), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12263), .COUT(n12264), .S0(n131_adj_1196), 
          .S1(n128_adj_1195));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_1225), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_1224), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12264), .COUT(n12265), .S0(n125_adj_1194), 
          .S1(n122_adj_1193));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_1223), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_1222), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12265), .COUT(n12266), .S0(n119_adj_1192), 
          .S1(n116_adj_1191));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_1221), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_1220), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12266), .COUT(n12267), .S0(n113_adj_1190), 
          .S1(n110_adj_1189));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_1219), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_1218), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12267), .COUT(n12268), .S0(n107_adj_1188), 
          .S1(n104_adj_1187));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_1217), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_1216), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12268), .COUT(n12269), .S0(n101_adj_1186), 
          .S1(n98_adj_1185));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_1215), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_1214), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12269), .COUT(n12270), .S0(n95_adj_1184), 
          .S1(n92_adj_1183));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_1213), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_1212), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12270), .COUT(n12271), .S0(n89_adj_1182), 
          .S1(n86_adj_1181));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_1211), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_1210), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12271), .COUT(n12272), .S0(n83_adj_1180), 
          .S1(n80_adj_1179));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_1209), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_1208), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12272), .COUT(n12273), .S0(n77_adj_1178), 
          .S1(n74_adj_1177));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_480_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_480_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_1207), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_1206), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12273), .S0(n71_adj_1176), .S1(n68_adj_1175));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_480_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_480_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_480_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_480_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n2072), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12278));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_477_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_477_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_3 (.A0(det_q4_28[0]), .B0(n2072), .C0(n161_adj_791), 
          .D0(n1098), .A1(n161_adj_1616), .B1(n2072), .C1(n158_adj_1267), 
          .D1(n1097), .CIN(n12278), .COUT(n12279), .S0(n161_adj_1236), 
          .S1(n158_adj_1235));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_5 (.A0(n158_adj_1615), .B0(n2072), .C0(n155_adj_1266), 
          .D0(n1096), .A1(n155_adj_1614), .B1(n2072), .C1(n152_adj_1265), 
          .D1(n1095), .CIN(n12279), .COUT(n12280), .S0(n155_adj_1234), 
          .S1(n152_adj_1233));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_7 (.A0(n152_adj_1613), .B0(n2072), .C0(n149_adj_1264), 
          .D0(n1094), .A1(n149_adj_1612), .B1(n2072), .C1(n146_adj_1263), 
          .D1(n1093), .CIN(n12280), .COUT(n12281), .S0(n149_adj_1232), 
          .S1(n146_adj_1231));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_9 (.A0(n146_adj_1611), .B0(n2072), .C0(n143_adj_1262), 
          .D0(n1092), .A1(n143_adj_1610), .B1(n2072), .C1(n140_adj_1261), 
          .D1(n1091), .CIN(n12281), .COUT(n12282), .S0(n143_adj_1230), 
          .S1(n140_adj_1229));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_11 (.A0(n140_adj_1609), .B0(n2072), .C0(n137_adj_1260), 
          .D0(n1090), .A1(n137_adj_1608), .B1(n2072), .C1(n134_adj_1259), 
          .D1(n1089), .CIN(n12282), .COUT(n12283), .S0(n137_adj_1228), 
          .S1(n134_adj_1227));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_13 (.A0(n134_adj_1607), .B0(n2072), .C0(n131_adj_1258), 
          .D0(n1088), .A1(n131_adj_1606), .B1(n2072), .C1(n128_adj_1257), 
          .D1(n1087), .CIN(n12283), .COUT(n12284), .S0(n131_adj_1226), 
          .S1(n128_adj_1225));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_15 (.A0(n128_adj_1605), .B0(n2072), .C0(n125_adj_1256), 
          .D0(n1086), .A1(n125_adj_1604), .B1(n2072), .C1(n122_adj_1255), 
          .D1(n1085), .CIN(n12284), .COUT(n12285), .S0(n125_adj_1224), 
          .S1(n122_adj_1223));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_17 (.A0(n122_adj_1603), .B0(n2072), .C0(n119_adj_1254), 
          .D0(n1084), .A1(n119_adj_1602), .B1(n2072), .C1(n116_adj_1253), 
          .D1(n1083), .CIN(n12285), .COUT(n12286), .S0(n119_adj_1222), 
          .S1(n116_adj_1221));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_19 (.A0(n116_adj_1601), .B0(n2072), .C0(n113_adj_1252), 
          .D0(n1082), .A1(n113_adj_1600), .B1(n2072), .C1(n110_adj_1251), 
          .D1(n1081), .CIN(n12286), .COUT(n12287), .S0(n113_adj_1220), 
          .S1(n110_adj_1219));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_21 (.A0(n110_adj_1599), .B0(n2072), .C0(n107_adj_1250), 
          .D0(n1080), .A1(n107_adj_1598), .B1(n2072), .C1(n104_adj_1249), 
          .D1(n1079), .CIN(n12287), .COUT(n12288), .S0(n107_adj_1218), 
          .S1(n104_adj_1217));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_23 (.A0(n104_adj_1597), .B0(n2072), .C0(n101_adj_1248), 
          .D0(n1078), .A1(n101_adj_1596), .B1(n2072), .C1(n98_adj_1247), 
          .D1(n1077), .CIN(n12288), .COUT(n12289), .S0(n101_adj_1216), 
          .S1(n98_adj_1215));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_25 (.A0(n98_adj_1595), .B0(n2072), .C0(n95_adj_1246), 
          .D0(n1076), .A1(n95_adj_1594), .B1(n2072), .C1(n92_adj_1245), 
          .D1(n1075), .CIN(n12289), .COUT(n12290), .S0(n95_adj_1214), 
          .S1(n92_adj_1213));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_27 (.A0(n92_adj_1593), .B0(n2072), .C0(n89_adj_1244), 
          .D0(n1074), .A1(n89_adj_1592), .B1(n2072), .C1(n86_adj_1243), 
          .D1(n1073), .CIN(n12290), .COUT(n12291), .S0(n89_adj_1212), 
          .S1(n86_adj_1211));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_29 (.A0(n86_adj_1591), .B0(n2072), .C0(n83_adj_1242), 
          .D0(n1072), .A1(n83_adj_1590), .B1(n2072), .C1(n80_adj_1241), 
          .D1(n1071), .CIN(n12291), .COUT(n12292), .S0(n83_adj_1210), 
          .S1(n80_adj_1209));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_31 (.A0(n80_adj_1589), .B0(n2072), .C0(n77_adj_1240), 
          .D0(n1070), .A1(n77_adj_1588), .B1(n2072), .C1(n74_adj_1239), 
          .D1(n1069), .CIN(n12292), .COUT(n12293), .S0(n77_adj_1208), 
          .S1(n74_adj_1207));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_477_add_4_33 (.A0(n74_adj_1587), .B0(n2072), .C0(n71_adj_1238), 
          .D0(n1068), .A1(n71_adj_1586), .B1(n2072), .C1(n68_adj_1237), 
          .D1(n1067), .CIN(n12293), .S0(n71_adj_1206), .S1(n2139));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_477_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_477_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_477_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_477_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_1616), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12296), .S1(n158_adj_1267));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_474_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_1615), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_1614), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12296), .COUT(n12297), .S0(n155_adj_1266), 
          .S1(n152_adj_1265));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_1613), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_1612), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12297), .COUT(n12298), .S0(n149_adj_1264), 
          .S1(n146_adj_1263));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_1611), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_1610), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12298), .COUT(n12299), .S0(n143_adj_1262), 
          .S1(n140_adj_1261));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_1609), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_1608), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12299), .COUT(n12300), .S0(n137_adj_1260), 
          .S1(n134_adj_1259));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_1607), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_1606), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12300), .COUT(n12301), .S0(n131_adj_1258), 
          .S1(n128_adj_1257));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_1605), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_1604), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12301), .COUT(n12302), .S0(n125_adj_1256), 
          .S1(n122_adj_1255));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_1603), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_1602), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12302), .COUT(n12303), .S0(n119_adj_1254), 
          .S1(n116_adj_1253));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_1601), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_1600), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12303), .COUT(n12304), .S0(n113_adj_1252), 
          .S1(n110_adj_1251));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_1599), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_1598), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12304), .COUT(n12305), .S0(n107_adj_1250), 
          .S1(n104_adj_1249));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_1597), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_1596), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12305), .COUT(n12306), .S0(n101_adj_1248), 
          .S1(n98_adj_1247));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_1595), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_1594), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12306), .COUT(n12307), .S0(n95_adj_1246), 
          .S1(n92_adj_1245));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_1593), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_1592), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12307), .COUT(n12308), .S0(n89_adj_1244), 
          .S1(n86_adj_1243));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_1591), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_1590), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12308), .COUT(n12309), .S0(n83_adj_1242), 
          .S1(n80_adj_1241));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_1589), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_1588), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12309), .COUT(n12310), .S0(n77_adj_1240), 
          .S1(n74_adj_1239));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_474_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_474_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_1587), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_1586), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12310), .S0(n71_adj_1238), .S1(n68_adj_1237));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_474_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_474_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_474_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_474_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_2 (.A0(n1098), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1097), .B1(n161_adj_853), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12313), .S1(n158_adj_1298));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_471_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_4 (.A0(n1096), .B0(n158_adj_852), .C0(GND_net), 
          .D0(VCC_net), .A1(n1095), .B1(n155_adj_851), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12313), .COUT(n12314), .S0(n155_adj_1297), 
          .S1(n152_adj_1296));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_6 (.A0(n1094), .B0(n152_adj_850), .C0(GND_net), 
          .D0(VCC_net), .A1(n1093), .B1(n149_adj_849), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12314), .COUT(n12315), .S0(n149_adj_1295), 
          .S1(n146_adj_1294));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_8 (.A0(n1092), .B0(n146_adj_848), .C0(GND_net), 
          .D0(VCC_net), .A1(n1091), .B1(n143_adj_847), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12315), .COUT(n12316), .S0(n143_adj_1293), 
          .S1(n140_adj_1292));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_10 (.A0(n1090), .B0(n140_adj_846), .C0(GND_net), 
          .D0(VCC_net), .A1(n1089), .B1(n137_adj_845), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12316), .COUT(n12317), .S0(n137_adj_1291), 
          .S1(n134_adj_1290));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_12 (.A0(n1088), .B0(n134_adj_844), .C0(GND_net), 
          .D0(VCC_net), .A1(n1087), .B1(n131_adj_843), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12317), .COUT(n12318), .S0(n131_adj_1289), 
          .S1(n128_adj_1288));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_14 (.A0(n1086), .B0(n128_adj_842), .C0(GND_net), 
          .D0(VCC_net), .A1(n1085), .B1(n125_adj_841), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12318), .COUT(n12319), .S0(n125_adj_1287), 
          .S1(n122_adj_1286));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_16 (.A0(n1084), .B0(n122_adj_840), .C0(GND_net), 
          .D0(VCC_net), .A1(n1083), .B1(n119_adj_839), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12319), .COUT(n12320), .S0(n119_adj_1285), 
          .S1(n116_adj_1284));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_18 (.A0(n1082), .B0(n116_adj_838), .C0(GND_net), 
          .D0(VCC_net), .A1(n1081), .B1(n113_adj_837), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12320), .COUT(n12321), .S0(n113_adj_1283), 
          .S1(n110_adj_1282));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_20 (.A0(n1080), .B0(n110_adj_836), .C0(GND_net), 
          .D0(VCC_net), .A1(n1079), .B1(n107_adj_835), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12321), .COUT(n12322), .S0(n107_adj_1281), 
          .S1(n104_adj_1280));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_22 (.A0(n1078), .B0(n104_adj_834), .C0(GND_net), 
          .D0(VCC_net), .A1(n1077), .B1(n101_adj_833), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12322), .COUT(n12323), .S0(n101_adj_1279), 
          .S1(n98_adj_1278));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_24 (.A0(n1076), .B0(n98_adj_832), .C0(GND_net), 
          .D0(VCC_net), .A1(n1075), .B1(n95_adj_831), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12323), .COUT(n12324), .S0(n95_adj_1277), 
          .S1(n92_adj_1276));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_26 (.A0(n1074), .B0(n92_adj_830), .C0(GND_net), 
          .D0(VCC_net), .A1(n1073), .B1(n89_adj_829), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12324), .COUT(n12325), .S0(n89_adj_1275), 
          .S1(n86_adj_1274));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_28 (.A0(n1072), .B0(n86_adj_828), .C0(GND_net), 
          .D0(VCC_net), .A1(n1071), .B1(n83_adj_827), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12325), .COUT(n12326), .S0(n83_adj_1273), 
          .S1(n80_adj_1272));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_30 (.A0(n1070), .B0(n80_adj_826), .C0(GND_net), 
          .D0(VCC_net), .A1(n1069), .B1(n77_adj_825), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12326), .COUT(n12327), .S0(n77_adj_1271), 
          .S1(n74_adj_1270));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_471_add_4_32 (.A0(n1068), .B0(n74_adj_824), .C0(GND_net), 
          .D0(VCC_net), .A1(n1067), .B1(n71_adj_823), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12327), .S0(n71_adj_1269), .S1(n68_adj_1268));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_471_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_471_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_471_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_471_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_2 (.A0(det_q4_28[1]), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[2]), .B1(n161_adj_853), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12330), .S1(n158_adj_1329));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_468_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_4 (.A0(det_q4_28[3]), .B0(n158_adj_852), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[4]), .B1(n155_adj_851), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12330), .COUT(n12331), .S0(n155_adj_1328), 
          .S1(n152_adj_1327));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_6 (.A0(det_q4_28[5]), .B0(n152_adj_850), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[6]), .B1(n149_adj_849), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12331), .COUT(n12332), .S0(n149_adj_1326), 
          .S1(n146_adj_1325));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_8 (.A0(det_q4_28[7]), .B0(n146_adj_848), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[8]), .B1(n143_adj_847), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12332), .COUT(n12333), .S0(n143_adj_1324), 
          .S1(n140_adj_1323));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_10 (.A0(det_q4_28[9]), .B0(n140_adj_846), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[10]), .B1(n137_adj_845), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12333), .COUT(n12334), .S0(n137_adj_1322), 
          .S1(n134_adj_1321));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_12 (.A0(det_q4_28[11]), .B0(n134_adj_844), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[12]), .B1(n131_adj_843), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12334), .COUT(n12335), .S0(n131_adj_1320), 
          .S1(n128_adj_1319));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_14 (.A0(det_q4_28[13]), .B0(n128_adj_842), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[14]), .B1(n125_adj_841), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12335), .COUT(n12336), .S0(n125_adj_1318), 
          .S1(n122_adj_1317));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_16 (.A0(det_q4_28[15]), .B0(n122_adj_840), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[16]), .B1(n119_adj_839), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12336), .COUT(n12337), .S0(n119_adj_1316), 
          .S1(n116_adj_1315));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_18 (.A0(det_q4_28[17]), .B0(n116_adj_838), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[18]), .B1(n113_adj_837), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12337), .COUT(n12338), .S0(n113_adj_1314), 
          .S1(n110_adj_1313));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_20 (.A0(det_q4_28[19]), .B0(n110_adj_836), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[20]), .B1(n107_adj_835), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12338), .COUT(n12339), .S0(n107_adj_1312), 
          .S1(n104_adj_1311));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_22 (.A0(det_q4_28[21]), .B0(n104_adj_834), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[22]), .B1(n101_adj_833), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12339), .COUT(n12340), .S0(n101_adj_1310), 
          .S1(n98_adj_1309));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_24 (.A0(det_q4_28[23]), .B0(n98_adj_832), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[24]), .B1(n95_adj_831), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12340), .COUT(n12341), .S0(n95_adj_1308), 
          .S1(n92_adj_1307));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_26 (.A0(det_q4_28[25]), .B0(n92_adj_830), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[26]), .B1(n89_adj_829), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12341), .COUT(n12342), .S0(n89_adj_1306), 
          .S1(n86_adj_1305));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_28 (.A0(det_q4_28[27]), .B0(n86_adj_828), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[28]), .B1(n83_adj_827), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12342), .COUT(n12343), .S0(n83_adj_1304), 
          .S1(n80_adj_1303));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_30 (.A0(det_q4_28[29]), .B0(n80_adj_826), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[30]), .B1(n77_adj_825), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12343), .COUT(n12344), .S0(n77_adj_1302), 
          .S1(n74_adj_1301));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_468_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_468_add_4_32 (.A0(det_q4_28[31]), .B0(n74_adj_824), .C0(GND_net), 
          .D0(VCC_net), .A1(n71_adj_823), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12344), .S0(n71_adj_1300), .S1(n68_adj_1299));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_468_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_468_add_4_32.INIT1 = 16'haaa0;
    defparam _add_1_468_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_468_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13022), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12346), .S1(n161_adj_1361));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_465_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_3 (.A0(n161_adj_1174), .B0(n13022), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1298), .B1(n13022), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12346), .COUT(n12347), .S0(n158_adj_1360), 
          .S1(n155_adj_1359));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_5 (.A0(n155_adj_1297), .B0(n13022), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1296), .B1(n13022), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12347), .COUT(n12348), .S0(n152_adj_1358), 
          .S1(n149_adj_1357));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_7 (.A0(n149_adj_1295), .B0(n13022), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1294), .B1(n13022), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12348), .COUT(n12349), .S0(n146_adj_1356), 
          .S1(n143_adj_1355));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_9 (.A0(n143_adj_1293), .B0(n13022), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1292), .B1(n13022), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12349), .COUT(n12350), .S0(n140_adj_1354), 
          .S1(n137_adj_1353));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_11 (.A0(n137_adj_1291), .B0(n13022), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1290), .B1(n13022), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12350), .COUT(n12351), .S0(n134_adj_1352), 
          .S1(n131_adj_1351));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_13 (.A0(n131_adj_1289), .B0(n13022), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1288), .B1(n13022), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12351), .COUT(n12352), .S0(n128_adj_1350), 
          .S1(n125_adj_1349));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_15 (.A0(n125_adj_1287), .B0(n13022), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1286), .B1(n13022), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12352), .COUT(n12353), .S0(n122_adj_1348), 
          .S1(n119_adj_1347));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_17 (.A0(n119_adj_1285), .B0(n13022), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1284), .B1(n13022), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12353), .COUT(n12354), .S0(n116_adj_1346), 
          .S1(n113_adj_1345));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_19 (.A0(n113_adj_1283), .B0(n13022), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1282), .B1(n13022), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12354), .COUT(n12355), .S0(n110_adj_1344), 
          .S1(n107_adj_1343));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_21 (.A0(n107_adj_1281), .B0(n13022), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1280), .B1(n13022), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12355), .COUT(n12356), .S0(n104_adj_1342), 
          .S1(n101_adj_1341));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_23 (.A0(n101_adj_1279), .B0(n13022), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1278), .B1(n13022), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12356), .COUT(n12357), .S0(n98_adj_1340), 
          .S1(n95_adj_1339));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_25 (.A0(n95_adj_1277), .B0(n13022), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1276), .B1(n13022), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12357), .COUT(n12358), .S0(n92_adj_1338), 
          .S1(n89_adj_1337));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_27 (.A0(n89_adj_1275), .B0(n13022), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1274), .B1(n13022), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12358), .COUT(n12359), .S0(n86_adj_1336), 
          .S1(n83_adj_1335));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_29 (.A0(n83_adj_1273), .B0(n13022), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1272), .B1(n13022), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12359), .COUT(n12360), .S0(n80_adj_1334), 
          .S1(n77_adj_1333));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_31 (.A0(n77_adj_1271), .B0(n13022), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1270), .B1(n13022), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12360), .COUT(n12361), .S0(n74_adj_1332), 
          .S1(n71_adj_1331));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_465_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_465_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_465_add_4_33 (.A0(n1067), .B0(n13022), .C0(n71_adj_1269), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12361), .S0(n68_adj_1330));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_465_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_465_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_465_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_465_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13022), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12362), .S1(n161_adj_1393));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_462_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_3 (.A0(n161_adj_791), .B0(n13022), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1329), .B1(n13022), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12362), .COUT(n12363), .S0(n158_adj_1392), 
          .S1(n155_adj_1391));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_5 (.A0(n155_adj_1328), .B0(n13022), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1327), .B1(n13022), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12363), .COUT(n12364), .S0(n152_adj_1390), 
          .S1(n149_adj_1389));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_7 (.A0(n149_adj_1326), .B0(n13022), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1325), .B1(n13022), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12364), .COUT(n12365), .S0(n146_adj_1388), 
          .S1(n143_adj_1387));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_9 (.A0(n143_adj_1324), .B0(n13022), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1323), .B1(n13022), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12365), .COUT(n12366), .S0(n140_adj_1386), 
          .S1(n137_adj_1385));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_11 (.A0(n137_adj_1322), .B0(n13022), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1321), .B1(n13022), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12366), .COUT(n12367), .S0(n134_adj_1384), 
          .S1(n131_adj_1383));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_13 (.A0(n131_adj_1320), .B0(n13022), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1319), .B1(n13022), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12367), .COUT(n12368), .S0(n128_adj_1382), 
          .S1(n125_adj_1381));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_15 (.A0(n125_adj_1318), .B0(n13022), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1317), .B1(n13022), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12368), .COUT(n12369), .S0(n122_adj_1380), 
          .S1(n119_adj_1379));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_17 (.A0(n119_adj_1316), .B0(n13022), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1315), .B1(n13022), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12369), .COUT(n12370), .S0(n116_adj_1378), 
          .S1(n113_adj_1377));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_19 (.A0(n113_adj_1314), .B0(n13022), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1313), .B1(n13022), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12370), .COUT(n12371), .S0(n110_adj_1376), 
          .S1(n107_adj_1375));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_21 (.A0(n107_adj_1312), .B0(n13022), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1311), .B1(n13022), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12371), .COUT(n12372), .S0(n104_adj_1374), 
          .S1(n101_adj_1373));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_23 (.A0(n101_adj_1310), .B0(n13022), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1309), .B1(n13022), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12372), .COUT(n12373), .S0(n98_adj_1372), 
          .S1(n95_adj_1371));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_25 (.A0(n95_adj_1308), .B0(n13022), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1307), .B1(n13022), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12373), .COUT(n12374), .S0(n92_adj_1370), 
          .S1(n89_adj_1369));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_27 (.A0(n89_adj_1306), .B0(n13022), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1305), .B1(n13022), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12374), .COUT(n12375), .S0(n86_adj_1368), 
          .S1(n83_adj_1367));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_29 (.A0(n83_adj_1304), .B0(n13022), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1303), .B1(n13022), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12375), .COUT(n12376), .S0(n80_adj_1366), 
          .S1(n77_adj_1365));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_31 (.A0(n77_adj_1302), .B0(n13022), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1301), .B1(n13022), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12376), .COUT(n12377), .S0(n74_adj_1364), 
          .S1(n71_adj_1363));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_462_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_462_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_462_add_4_33 (.A0(n1067), .B0(n13022), .C0(n71_adj_1300), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12377), .S0(n68_adj_1362));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_462_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_462_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_462_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_462_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13021), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12378), .S1(n161_adj_1425));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_459_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_3 (.A0(n161_adj_1361), .B0(n13021), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1360), .B1(n13021), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12378), .COUT(n12379), .S0(n158_adj_1424), 
          .S1(n155_adj_1423));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_5 (.A0(n155_adj_1359), .B0(n13021), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1358), .B1(n13021), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12379), .COUT(n12380), .S0(n152_adj_1422), 
          .S1(n149_adj_1421));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_7 (.A0(n149_adj_1357), .B0(n13021), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1356), .B1(n13021), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12380), .COUT(n12381), .S0(n146_adj_1420), 
          .S1(n143_adj_1419));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_9 (.A0(n143_adj_1355), .B0(n13021), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1354), .B1(n13021), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12381), .COUT(n12382), .S0(n140_adj_1418), 
          .S1(n137_adj_1417));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_11 (.A0(n137_adj_1353), .B0(n13021), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1352), .B1(n13021), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12382), .COUT(n12383), .S0(n134_adj_1416), 
          .S1(n131_adj_1415));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_13 (.A0(n131_adj_1351), .B0(n13021), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1350), .B1(n13021), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12383), .COUT(n12384), .S0(n128_adj_1414), 
          .S1(n125_adj_1413));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_15 (.A0(n125_adj_1349), .B0(n13021), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1348), .B1(n13021), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12384), .COUT(n12385), .S0(n122_adj_1412), 
          .S1(n119_adj_1411));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_17 (.A0(n119_adj_1347), .B0(n13021), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1346), .B1(n13021), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12385), .COUT(n12386), .S0(n116_adj_1410), 
          .S1(n113_adj_1409));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_19 (.A0(n113_adj_1345), .B0(n13021), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1344), .B1(n13021), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12386), .COUT(n12387), .S0(n110_adj_1408), 
          .S1(n107_adj_1407));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_21 (.A0(n107_adj_1343), .B0(n13021), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1342), .B1(n13021), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12387), .COUT(n12388), .S0(n104_adj_1406), 
          .S1(n101_adj_1405));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_23 (.A0(n101_adj_1341), .B0(n13021), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1340), .B1(n13021), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12388), .COUT(n12389), .S0(n98_adj_1404), 
          .S1(n95_adj_1403));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_25 (.A0(n95_adj_1339), .B0(n13021), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1338), .B1(n13021), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12389), .COUT(n12390), .S0(n92_adj_1402), 
          .S1(n89_adj_1401));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_27 (.A0(n89_adj_1337), .B0(n13021), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1336), .B1(n13021), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12390), .COUT(n12391), .S0(n86_adj_1400), 
          .S1(n83_adj_1399));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_29 (.A0(n83_adj_1335), .B0(n13021), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1334), .B1(n13021), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12391), .COUT(n12392), .S0(n80_adj_1398), 
          .S1(n77_adj_1397));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_31 (.A0(n77_adj_1333), .B0(n13021), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1332), .B1(n13021), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12392), .COUT(n12393), .S0(n74_adj_1396), 
          .S1(n71_adj_1395));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_459_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_459_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_459_add_4_33 (.A0(n1067), .B0(n13021), .C0(n71_adj_1331), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12393), .S0(n68_adj_1394));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_459_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_459_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_459_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_459_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13021), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12394), .S1(n161_adj_1457));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_456_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_3 (.A0(n161_adj_1393), .B0(n13021), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1392), .B1(n13021), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12394), .COUT(n12395), .S0(n158_adj_1456), 
          .S1(n155_adj_1455));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_5 (.A0(n155_adj_1391), .B0(n13021), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1390), .B1(n13021), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12395), .COUT(n12396), .S0(n152_adj_1454), 
          .S1(n149_adj_1453));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_7 (.A0(n149_adj_1389), .B0(n13021), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1388), .B1(n13021), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12396), .COUT(n12397), .S0(n146_adj_1452), 
          .S1(n143_adj_1451));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_9 (.A0(n143_adj_1387), .B0(n13021), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1386), .B1(n13021), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12397), .COUT(n12398), .S0(n140_adj_1450), 
          .S1(n137_adj_1449));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_11 (.A0(n137_adj_1385), .B0(n13021), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1384), .B1(n13021), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12398), .COUT(n12399), .S0(n134_adj_1448), 
          .S1(n131_adj_1447));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_13 (.A0(n131_adj_1383), .B0(n13021), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1382), .B1(n13021), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12399), .COUT(n12400), .S0(n128_adj_1446), 
          .S1(n125_adj_1445));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_15 (.A0(n125_adj_1381), .B0(n13021), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1380), .B1(n13021), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12400), .COUT(n12401), .S0(n122_adj_1444), 
          .S1(n119_adj_1443));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_17 (.A0(n119_adj_1379), .B0(n13021), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1378), .B1(n13021), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12401), .COUT(n12402), .S0(n116_adj_1442), 
          .S1(n113_adj_1441));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_19 (.A0(n113_adj_1377), .B0(n13021), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1376), .B1(n13021), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12402), .COUT(n12403), .S0(n110_adj_1440), 
          .S1(n107_adj_1439));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_21 (.A0(n107_adj_1375), .B0(n13021), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1374), .B1(n13021), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12403), .COUT(n12404), .S0(n104_adj_1438), 
          .S1(n101_adj_1437));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_23 (.A0(n101_adj_1373), .B0(n13021), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1372), .B1(n13021), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12404), .COUT(n12405), .S0(n98_adj_1436), 
          .S1(n95_adj_1435));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_25 (.A0(n95_adj_1371), .B0(n13021), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1370), .B1(n13021), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12405), .COUT(n12406), .S0(n92_adj_1434), 
          .S1(n89_adj_1433));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_27 (.A0(n89_adj_1369), .B0(n13021), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1368), .B1(n13021), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12406), .COUT(n12407), .S0(n86_adj_1432), 
          .S1(n83_adj_1431));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_29 (.A0(n83_adj_1367), .B0(n13021), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1366), .B1(n13021), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12407), .COUT(n12408), .S0(n80_adj_1430), 
          .S1(n77_adj_1429));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_31 (.A0(n77_adj_1365), .B0(n13021), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1364), .B1(n13021), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12408), .COUT(n12409), .S0(n74_adj_1428), 
          .S1(n71_adj_1427));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_456_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_456_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_456_add_4_33 (.A0(n1067), .B0(n13021), .C0(n71_adj_1363), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12409), .S0(n68_adj_1426));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_456_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_456_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_456_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_456_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13020), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12410), .S1(n161_adj_1489));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_453_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_3 (.A0(n161_adj_1425), .B0(n13020), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1424), .B1(n13020), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12410), .COUT(n12411), .S0(n158_adj_1488), 
          .S1(n155_adj_1487));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_5 (.A0(n155_adj_1423), .B0(n13020), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1422), .B1(n13020), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12411), .COUT(n12412), .S0(n152_adj_1486), 
          .S1(n149_adj_1485));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_7 (.A0(n149_adj_1421), .B0(n13020), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1420), .B1(n13020), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12412), .COUT(n12413), .S0(n146_adj_1484), 
          .S1(n143_adj_1483));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_9 (.A0(n143_adj_1419), .B0(n13020), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1418), .B1(n13020), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12413), .COUT(n12414), .S0(n140_adj_1482), 
          .S1(n137_adj_1481));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_11 (.A0(n137_adj_1417), .B0(n13020), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1416), .B1(n13020), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12414), .COUT(n12415), .S0(n134_adj_1480), 
          .S1(n131_adj_1479));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_13 (.A0(n131_adj_1415), .B0(n13020), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1414), .B1(n13020), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12415), .COUT(n12416), .S0(n128_adj_1478), 
          .S1(n125_adj_1477));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_15 (.A0(n125_adj_1413), .B0(n13020), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1412), .B1(n13020), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12416), .COUT(n12417), .S0(n122_adj_1476), 
          .S1(n119_adj_1475));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_17 (.A0(n119_adj_1411), .B0(n13020), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1410), .B1(n13020), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12417), .COUT(n12418), .S0(n116_adj_1474), 
          .S1(n113_adj_1473));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_19 (.A0(n113_adj_1409), .B0(n13020), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1408), .B1(n13020), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12418), .COUT(n12419), .S0(n110_adj_1472), 
          .S1(n107_adj_1471));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_21 (.A0(n107_adj_1407), .B0(n13020), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1406), .B1(n13020), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12419), .COUT(n12420), .S0(n104_adj_1470), 
          .S1(n101_adj_1469));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_23 (.A0(n101_adj_1405), .B0(n13020), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1404), .B1(n13020), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12420), .COUT(n12421), .S0(n98_adj_1468), 
          .S1(n95_adj_1467));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_25 (.A0(n95_adj_1403), .B0(n13020), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1402), .B1(n13020), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12421), .COUT(n12422), .S0(n92_adj_1466), 
          .S1(n89_adj_1465));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_27 (.A0(n89_adj_1401), .B0(n13020), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1400), .B1(n13020), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12422), .COUT(n12423), .S0(n86_adj_1464), 
          .S1(n83_adj_1463));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_29 (.A0(n83_adj_1399), .B0(n13020), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1398), .B1(n13020), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12423), .COUT(n12424), .S0(n80_adj_1462), 
          .S1(n77_adj_1461));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_31 (.A0(n77_adj_1397), .B0(n13020), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1396), .B1(n13020), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12424), .COUT(n12425), .S0(n74_adj_1460), 
          .S1(n71_adj_1459));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_453_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_453_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_453_add_4_33 (.A0(n1067), .B0(n13020), .C0(n71_adj_1395), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12425), .S0(n68_adj_1458));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_453_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_453_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_453_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_453_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13020), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12426), .S1(n161_adj_1521));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_450_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_3 (.A0(n161_adj_1457), .B0(n13020), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1456), .B1(n13020), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12426), .COUT(n12427), .S0(n158_adj_1520), 
          .S1(n155_adj_1519));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_5 (.A0(n155_adj_1455), .B0(n13020), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1454), .B1(n13020), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12427), .COUT(n12428), .S0(n152_adj_1518), 
          .S1(n149_adj_1517));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_7 (.A0(n149_adj_1453), .B0(n13020), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1452), .B1(n13020), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12428), .COUT(n12429), .S0(n146_adj_1516), 
          .S1(n143_adj_1515));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_9 (.A0(n143_adj_1451), .B0(n13020), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1450), .B1(n13020), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12429), .COUT(n12430), .S0(n140_adj_1514), 
          .S1(n137_adj_1513));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_11 (.A0(n137_adj_1449), .B0(n13020), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1448), .B1(n13020), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12430), .COUT(n12431), .S0(n134_adj_1512), 
          .S1(n131_adj_1511));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_13 (.A0(n131_adj_1447), .B0(n13020), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1446), .B1(n13020), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12431), .COUT(n12432), .S0(n128_adj_1510), 
          .S1(n125_adj_1509));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_15 (.A0(n125_adj_1445), .B0(n13020), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1444), .B1(n13020), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12432), .COUT(n12433), .S0(n122_adj_1508), 
          .S1(n119_adj_1507));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_17 (.A0(n119_adj_1443), .B0(n13020), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1442), .B1(n13020), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12433), .COUT(n12434), .S0(n116_adj_1506), 
          .S1(n113_adj_1505));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_19 (.A0(n113_adj_1441), .B0(n13020), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1440), .B1(n13020), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12434), .COUT(n12435), .S0(n110_adj_1504), 
          .S1(n107_adj_1503));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_21 (.A0(n107_adj_1439), .B0(n13020), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1438), .B1(n13020), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12435), .COUT(n12436), .S0(n104_adj_1502), 
          .S1(n101_adj_1501));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_23 (.A0(n101_adj_1437), .B0(n13020), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1436), .B1(n13020), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12436), .COUT(n12437), .S0(n98_adj_1500), 
          .S1(n95_adj_1499));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_25 (.A0(n95_adj_1435), .B0(n13020), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1434), .B1(n13020), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12437), .COUT(n12438), .S0(n92_adj_1498), 
          .S1(n89_adj_1497));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_27 (.A0(n89_adj_1433), .B0(n13020), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1432), .B1(n13020), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12438), .COUT(n12439), .S0(n86_adj_1496), 
          .S1(n83_adj_1495));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_29 (.A0(n83_adj_1431), .B0(n13020), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1430), .B1(n13020), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12439), .COUT(n12440), .S0(n80_adj_1494), 
          .S1(n77_adj_1493));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_31 (.A0(n77_adj_1429), .B0(n13020), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1428), .B1(n13020), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12440), .COUT(n12441), .S0(n74_adj_1492), 
          .S1(n71_adj_1491));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_450_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_450_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_450_add_4_33 (.A0(n1067), .B0(n13020), .C0(n71_adj_1427), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12441), .S0(n68_adj_1490));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_450_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_450_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_450_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_450_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13019), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12442), .S1(n161_adj_1553));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_447_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_3 (.A0(n161_adj_1489), .B0(n13019), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1488), .B1(n13019), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12442), .COUT(n12443), .S0(n158_adj_1552), 
          .S1(n155_adj_1551));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_5 (.A0(n155_adj_1487), .B0(n13019), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1486), .B1(n13019), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12443), .COUT(n12444), .S0(n152_adj_1550), 
          .S1(n149_adj_1549));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_7 (.A0(n149_adj_1485), .B0(n13019), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1484), .B1(n13019), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12444), .COUT(n12445), .S0(n146_adj_1548), 
          .S1(n143_adj_1547));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_9 (.A0(n143_adj_1483), .B0(n13019), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1482), .B1(n13019), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12445), .COUT(n12446), .S0(n140_adj_1546), 
          .S1(n137_adj_1545));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_11 (.A0(n137_adj_1481), .B0(n13019), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1480), .B1(n13019), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12446), .COUT(n12447), .S0(n134_adj_1544), 
          .S1(n131_adj_1543));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_13 (.A0(n131_adj_1479), .B0(n13019), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1478), .B1(n13019), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12447), .COUT(n12448), .S0(n128_adj_1542), 
          .S1(n125_adj_1541));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_15 (.A0(n125_adj_1477), .B0(n13019), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1476), .B1(n13019), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12448), .COUT(n12449), .S0(n122_adj_1540), 
          .S1(n119_adj_1539));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_17 (.A0(n119_adj_1475), .B0(n13019), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1474), .B1(n13019), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12449), .COUT(n12450), .S0(n116_adj_1538), 
          .S1(n113_adj_1537));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_19 (.A0(n113_adj_1473), .B0(n13019), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1472), .B1(n13019), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12450), .COUT(n12451), .S0(n110_adj_1536), 
          .S1(n107_adj_1535));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_21 (.A0(n107_adj_1471), .B0(n13019), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1470), .B1(n13019), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12451), .COUT(n12452), .S0(n104_adj_1534), 
          .S1(n101_adj_1533));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_23 (.A0(n101_adj_1469), .B0(n13019), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1468), .B1(n13019), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12452), .COUT(n12453), .S0(n98_adj_1532), 
          .S1(n95_adj_1531));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_25 (.A0(n95_adj_1467), .B0(n13019), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1466), .B1(n13019), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12453), .COUT(n12454), .S0(n92_adj_1530), 
          .S1(n89_adj_1529));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_27 (.A0(n89_adj_1465), .B0(n13019), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1464), .B1(n13019), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12454), .COUT(n12455), .S0(n86_adj_1528), 
          .S1(n83_adj_1527));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_29 (.A0(n83_adj_1463), .B0(n13019), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1462), .B1(n13019), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12455), .COUT(n12456), .S0(n80_adj_1526), 
          .S1(n77_adj_1525));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_31 (.A0(n77_adj_1461), .B0(n13019), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1460), .B1(n13019), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12456), .COUT(n12457), .S0(n74_adj_1524), 
          .S1(n71_adj_1523));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_447_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_447_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_447_add_4_33 (.A0(n1067), .B0(n13019), .C0(n71_adj_1459), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12457), .S0(n68_adj_1522));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_447_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_447_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_447_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_447_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28_31__N_65[0]), .B1(det_q4_28_31__N_33[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n12458), .S1(det_q4_28_31__N_1[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_417_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_4 (.A0(det_q4_28_31__N_65[1]), .B0(det_q4_28_31__N_33[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[2]), .B1(det_q4_28_31__N_33[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12458), .COUT(n12459), .S0(det_q4_28_31__N_1[1]), 
          .S1(det_q4_28_31__N_1[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_6 (.A0(det_q4_28_31__N_65[3]), .B0(det_q4_28_31__N_33[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[4]), .B1(det_q4_28_31__N_33[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12459), .COUT(n12460), .S0(det_q4_28_31__N_1[3]), 
          .S1(det_q4_28_31__N_1[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_8 (.A0(det_q4_28_31__N_65[5]), .B0(det_q4_28_31__N_33[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[6]), .B1(det_q4_28_31__N_33[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12460), .COUT(n12461), .S0(det_q4_28_31__N_1[5]), 
          .S1(det_q4_28_31__N_1[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_10 (.A0(det_q4_28_31__N_65[7]), .B0(det_q4_28_31__N_33[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[8]), .B1(det_q4_28_31__N_33[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12461), .COUT(n12462), .S0(det_q4_28_31__N_1[7]), 
          .S1(det_q4_28_31__N_1[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_12 (.A0(det_q4_28_31__N_65[9]), .B0(det_q4_28_31__N_33[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[10]), .B1(det_q4_28_31__N_33[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12462), .COUT(n12463), .S0(det_q4_28_31__N_1[9]), 
          .S1(det_q4_28_31__N_1[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_14 (.A0(det_q4_28_31__N_65[11]), .B0(det_q4_28_31__N_33[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[12]), .B1(det_q4_28_31__N_33[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12463), .COUT(n12464), .S0(det_q4_28_31__N_1[11]), 
          .S1(det_q4_28_31__N_1[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_16 (.A0(det_q4_28_31__N_65[13]), .B0(det_q4_28_31__N_33[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[14]), .B1(det_q4_28_31__N_33[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12464), .COUT(n12465), .S0(det_q4_28_31__N_1[13]), 
          .S1(det_q4_28_31__N_1[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_18 (.A0(det_q4_28_31__N_65[15]), .B0(det_q4_28_31__N_33[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[16]), .B1(det_q4_28_31__N_33[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12465), .COUT(n12466), .S0(det_q4_28_31__N_1[15]), 
          .S1(det_q4_28_31__N_1[16]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_20 (.A0(det_q4_28_31__N_65[17]), .B0(det_q4_28_31__N_33[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[18]), .B1(det_q4_28_31__N_33[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12466), .COUT(n12467), .S0(det_q4_28_31__N_1[17]), 
          .S1(det_q4_28_31__N_1[18]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_22 (.A0(det_q4_28_31__N_65[19]), .B0(det_q4_28_31__N_33[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[20]), .B1(det_q4_28_31__N_33[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12467), .COUT(n12468), .S0(det_q4_28_31__N_1[19]), 
          .S1(det_q4_28_31__N_1[20]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_24 (.A0(det_q4_28_31__N_65[21]), .B0(det_q4_28_31__N_33[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[22]), .B1(det_q4_28_31__N_33[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12468), .COUT(n12469), .S0(det_q4_28_31__N_1[21]), 
          .S1(det_q4_28_31__N_1[22]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_26 (.A0(det_q4_28_31__N_65[23]), .B0(det_q4_28_31__N_33[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[24]), .B1(det_q4_28_31__N_33[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12469), .COUT(n12470), .S0(det_q4_28_31__N_1[23]), 
          .S1(det_q4_28_31__N_1[24]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_28 (.A0(det_q4_28_31__N_65[25]), .B0(det_q4_28_31__N_33[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[26]), .B1(det_q4_28_31__N_33[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12470), .COUT(n12471), .S0(det_q4_28_31__N_1[25]), 
          .S1(det_q4_28_31__N_1[26]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_30 (.A0(det_q4_28_31__N_65[27]), .B0(det_q4_28_31__N_33[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[28]), .B1(det_q4_28_31__N_33[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12471), .COUT(n12472), .S0(det_q4_28_31__N_1[27]), 
          .S1(det_q4_28_31__N_1[28]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_32 (.A0(det_q4_28_31__N_65[29]), .B0(det_q4_28_31__N_33[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(det_q4_28_31__N_65[30]), .B1(det_q4_28_31__N_33[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n12472), .COUT(n12473), .S0(det_q4_28_31__N_1[29]), 
          .S1(det_q4_28_31__N_1[30]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_417_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_417_add_4_34 (.A0(det_q4_28_31__N_65[31]), .B0(det_q4_28_31__N_33[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12473), .S0(det_q4_28_31__N_1[31]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(43[26:43])
    defparam _add_1_417_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_417_add_4_34.INIT1 = 16'h0000;
    defparam _add_1_417_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_417_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13028), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12474), .S1(n161_adj_1585));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_501_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_3 (.A0(n161_adj_1905), .B0(n13028), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1904), .B1(n13028), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12474), .COUT(n12475), .S0(n158_adj_1584), 
          .S1(n155_adj_1583));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_5 (.A0(n155_adj_1903), .B0(n13028), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1902), .B1(n13028), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12475), .COUT(n12476), .S0(n152_adj_1582), 
          .S1(n149_adj_1581));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_7 (.A0(n149_adj_1901), .B0(n13028), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1900), .B1(n13028), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12476), .COUT(n12477), .S0(n146_adj_1580), 
          .S1(n143_adj_1579));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_9 (.A0(n143_adj_1899), .B0(n13028), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1898), .B1(n13028), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12477), .COUT(n12478), .S0(n140_adj_1578), 
          .S1(n137_adj_1577));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_11 (.A0(n137_adj_1897), .B0(n13028), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1896), .B1(n13028), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12478), .COUT(n12479), .S0(n134_adj_1576), 
          .S1(n131_adj_1575));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_13 (.A0(n131_adj_1895), .B0(n13028), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1894), .B1(n13028), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12479), .COUT(n12480), .S0(n128_adj_1574), 
          .S1(n125_adj_1573));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_15 (.A0(n125_adj_1893), .B0(n13028), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1892), .B1(n13028), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12480), .COUT(n12481), .S0(n122_adj_1572), 
          .S1(n119_adj_1571));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_17 (.A0(n119_adj_1891), .B0(n13028), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1890), .B1(n13028), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12481), .COUT(n12482), .S0(n116_adj_1570), 
          .S1(n113_adj_1569));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_19 (.A0(n113_adj_1889), .B0(n13028), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1888), .B1(n13028), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12482), .COUT(n12483), .S0(n110_adj_1568), 
          .S1(n107_adj_1567));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_21 (.A0(n107_adj_1887), .B0(n13028), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1886), .B1(n13028), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12483), .COUT(n12484), .S0(n104_adj_1566), 
          .S1(n101_adj_1565));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_23 (.A0(n101_adj_1885), .B0(n13028), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1884), .B1(n13028), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12484), .COUT(n12485), .S0(n98_adj_1564), 
          .S1(n95_adj_1563));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_25 (.A0(n95_adj_1883), .B0(n13028), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1882), .B1(n13028), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12485), .COUT(n12486), .S0(n92_adj_1562), 
          .S1(n89_adj_1561));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_27 (.A0(n89_adj_1881), .B0(n13028), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1880), .B1(n13028), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12486), .COUT(n12487), .S0(n86_adj_1560), 
          .S1(n83_adj_1559));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_29 (.A0(n83_adj_1879), .B0(n13028), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1878), .B1(n13028), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12487), .COUT(n12488), .S0(n80_adj_1558), 
          .S1(n77_adj_1557));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_31 (.A0(n77_adj_1877), .B0(n13028), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1876), .B1(n13028), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12488), .COUT(n12489), .S0(n74_adj_1556), 
          .S1(n71_adj_1555));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_501_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_501_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_501_add_4_33 (.A0(n1067), .B0(n13028), .C0(n71_adj_1875), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12489), .S0(n68_adj_1554));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_501_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_501_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_501_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_501_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n1536), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12493));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_426_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_426_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_3 (.A0(det_q4_28[0]), .B0(n1536), .C0(n161_adj_1776), 
          .D0(n2070), .A1(n161_adj_1841), .B1(n1536), .C1(n158_adj_1775), 
          .D1(n2069), .CIN(n12493), .COUT(n12494), .S0(n161_adj_1616), 
          .S1(n158_adj_1615));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_3.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_3.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_5 (.A0(n158_adj_1840), .B0(n1536), .C0(n155_adj_1774), 
          .D0(n2068), .A1(n155_adj_1839), .B1(n1536), .C1(n152_adj_1773), 
          .D1(n2067), .CIN(n12494), .COUT(n12495), .S0(n155_adj_1614), 
          .S1(n152_adj_1613));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_5.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_5.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_7 (.A0(n152_adj_1838), .B0(n1536), .C0(n149_adj_1772), 
          .D0(n2066), .A1(n149_adj_1837), .B1(n1536), .C1(n146_adj_1771), 
          .D1(n2065), .CIN(n12495), .COUT(n12496), .S0(n149_adj_1612), 
          .S1(n146_adj_1611));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_7.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_7.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_9 (.A0(n146_adj_1836), .B0(n1536), .C0(n143_adj_1770), 
          .D0(n2064), .A1(n143_adj_1835), .B1(n1536), .C1(n140_adj_1769), 
          .D1(n2063), .CIN(n12496), .COUT(n12497), .S0(n143_adj_1610), 
          .S1(n140_adj_1609));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_9.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_9.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_11 (.A0(n140_adj_1834), .B0(n1536), .C0(n137_adj_1768), 
          .D0(n2062), .A1(n137_adj_1833), .B1(n1536), .C1(n134_adj_1767), 
          .D1(n2061), .CIN(n12497), .COUT(n12498), .S0(n137_adj_1608), 
          .S1(n134_adj_1607));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_11.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_11.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_13 (.A0(n134_adj_1832), .B0(n1536), .C0(n131_adj_1766), 
          .D0(n2060), .A1(n131_adj_1831), .B1(n1536), .C1(n128_adj_1765), 
          .D1(n2059), .CIN(n12498), .COUT(n12499), .S0(n131_adj_1606), 
          .S1(n128_adj_1605));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_13.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_13.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_15 (.A0(n128_adj_1830), .B0(n1536), .C0(n125_adj_1764), 
          .D0(n2058), .A1(n125_adj_1829), .B1(n1536), .C1(n122_adj_1763), 
          .D1(n2057), .CIN(n12499), .COUT(n12500), .S0(n125_adj_1604), 
          .S1(n122_adj_1603));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_15.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_15.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_17 (.A0(n122_adj_1828), .B0(n1536), .C0(n119_adj_1762), 
          .D0(n2056), .A1(n119_adj_1827), .B1(n1536), .C1(n116_adj_1761), 
          .D1(n2055), .CIN(n12500), .COUT(n12501), .S0(n119_adj_1602), 
          .S1(n116_adj_1601));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_17.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_17.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_19 (.A0(n116_adj_1826), .B0(n1536), .C0(n113_adj_1760), 
          .D0(n2054), .A1(n113_adj_1825), .B1(n1536), .C1(n110_adj_1759), 
          .D1(n2053), .CIN(n12501), .COUT(n12502), .S0(n113_adj_1600), 
          .S1(n110_adj_1599));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_19.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_19.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_21 (.A0(n110_adj_1824), .B0(n1536), .C0(n107_adj_1758), 
          .D0(n2052), .A1(n107_adj_1823), .B1(n1536), .C1(n104_adj_1757), 
          .D1(n2051), .CIN(n12502), .COUT(n12503), .S0(n107_adj_1598), 
          .S1(n104_adj_1597));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_21.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_21.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_23 (.A0(n104_adj_1822), .B0(n1536), .C0(n101_adj_1756), 
          .D0(n2050), .A1(n101_adj_1821), .B1(n1536), .C1(n98_adj_1755), 
          .D1(n2049), .CIN(n12503), .COUT(n12504), .S0(n101_adj_1596), 
          .S1(n98_adj_1595));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_23.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_23.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_25 (.A0(n98_adj_1820), .B0(n1536), .C0(n95_adj_1754), 
          .D0(n2048), .A1(n95_adj_1819), .B1(n1536), .C1(n92_adj_1753), 
          .D1(n2047), .CIN(n12504), .COUT(n12505), .S0(n95_adj_1594), 
          .S1(n92_adj_1593));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_25.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_25.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_27 (.A0(n92_adj_1818), .B0(n1536), .C0(n89_adj_1752), 
          .D0(n2046), .A1(n89_adj_1817), .B1(n1536), .C1(n86_adj_1751), 
          .D1(n2045), .CIN(n12505), .COUT(n12506), .S0(n89_adj_1592), 
          .S1(n86_adj_1591));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_27.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_27.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_29 (.A0(n86_adj_1816), .B0(n1536), .C0(n83_adj_1750), 
          .D0(n2044), .A1(n83_adj_1815), .B1(n1536), .C1(n80_adj_1749), 
          .D1(n2043), .CIN(n12506), .COUT(n12507), .S0(n83_adj_1590), 
          .S1(n80_adj_1589));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_29.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_29.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_31 (.A0(n80_adj_1814), .B0(n1536), .C0(n77_adj_1748), 
          .D0(n2042), .A1(n77_adj_1813), .B1(n1536), .C1(n74_adj_1747), 
          .D1(n2041), .CIN(n12507), .COUT(n12508), .S0(n77_adj_1588), 
          .S1(n74_adj_1587));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_31.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_31.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_426_add_4_33 (.A0(n74_adj_1812), .B0(n1536), .C0(n71_adj_1746), 
          .D0(n2040), .A1(n71_adj_1811), .B1(n1536), .C1(n68_adj_1745), 
          .D1(n2039), .CIN(n12508), .S0(n71_adj_1586), .S1(n2072));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_426_add_4_33.INIT0 = 16'h74b8;
    defparam _add_1_426_add_4_33.INIT1 = 16'h74b8;
    defparam _add_1_426_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_426_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13018), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12510), .S1(n161_adj_1648));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_438_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_3 (.A0(n161_adj_2129), .B0(n13018), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_2128), .B1(n13018), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12510), .COUT(n12511), .S0(n158_adj_1647), 
          .S1(n155_adj_1646));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_5 (.A0(n155_adj_2127), .B0(n13018), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_2126), .B1(n13018), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12511), .COUT(n12512), .S0(n152_adj_1645), 
          .S1(n149_adj_1644));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_7 (.A0(n149_adj_2125), .B0(n13018), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_2124), .B1(n13018), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12512), .COUT(n12513), .S0(n146_adj_1643), 
          .S1(n143_adj_1642));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_9 (.A0(n143_adj_2123), .B0(n13018), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_2122), .B1(n13018), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12513), .COUT(n12514), .S0(n140_adj_1641), 
          .S1(n137_adj_1640));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_11 (.A0(n137_adj_2121), .B0(n13018), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_2120), .B1(n13018), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12514), .COUT(n12515), .S0(n134_adj_1639), 
          .S1(n131_adj_1638));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_13 (.A0(n131_adj_2119), .B0(n13018), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_2118), .B1(n13018), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12515), .COUT(n12516), .S0(n128_adj_1637), 
          .S1(n125_adj_1636));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_15 (.A0(n125_adj_2117), .B0(n13018), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_2116), .B1(n13018), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12516), .COUT(n12517), .S0(n122_adj_1635), 
          .S1(n119_adj_1634));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_17 (.A0(n119_adj_2115), .B0(n13018), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_2114), .B1(n13018), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12517), .COUT(n12518), .S0(n116_adj_1633), 
          .S1(n113_adj_1632));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_19 (.A0(n113_adj_2113), .B0(n13018), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_2112), .B1(n13018), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12518), .COUT(n12519), .S0(n110_adj_1631), 
          .S1(n107_adj_1630));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_21 (.A0(n107_adj_2111), .B0(n13018), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_2110), .B1(n13018), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12519), .COUT(n12520), .S0(n104_adj_1629), 
          .S1(n101_adj_1628));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_23 (.A0(n101_adj_2109), .B0(n13018), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_2108), .B1(n13018), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12520), .COUT(n12521), .S0(n98_adj_1627), 
          .S1(n95_adj_1626));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_25 (.A0(n95_adj_2107), .B0(n13018), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_2106), .B1(n13018), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12521), .COUT(n12522), .S0(n92_adj_1625), 
          .S1(n89_adj_1624));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_27 (.A0(n89_adj_2105), .B0(n13018), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_2104), .B1(n13018), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12522), .COUT(n12523), .S0(n86_adj_1623), 
          .S1(n83_adj_1622));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_29 (.A0(n83_adj_2103), .B0(n13018), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_2102), .B1(n13018), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12523), .COUT(n12524), .S0(n80_adj_1621), 
          .S1(n77_adj_1620));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_31 (.A0(n77_adj_2101), .B0(n13018), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_2100), .B1(n13018), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12524), .COUT(n12525), .S0(n74_adj_1619), 
          .S1(n71_adj_1618));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_438_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_438_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_438_add_4_33 (.A0(n1067), .B0(n13018), .C0(n71_adj_2099), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12525), .S0(n68_adj_1617));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_438_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_438_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_438_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_438_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13009), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12526), .S1(n161_adj_1680));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_573_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_3 (.A0(n161_adj_1809), .B0(n13009), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1808), .B1(n13009), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12526), .COUT(n12527), .S0(n158_adj_1679), 
          .S1(n155_adj_1678));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_5 (.A0(n155_adj_1807), .B0(n13009), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1806), .B1(n13009), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12527), .COUT(n12528), .S0(n152_adj_1677), 
          .S1(n149_adj_1676));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_7 (.A0(n149_adj_1805), .B0(n13009), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1804), .B1(n13009), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12528), .COUT(n12529), .S0(n146_adj_1675), 
          .S1(n143_adj_1674));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_9 (.A0(n143_adj_1803), .B0(n13009), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1802), .B1(n13009), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12529), .COUT(n12530), .S0(n140_adj_1673), 
          .S1(n137_adj_1672));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_11 (.A0(n137_adj_1801), .B0(n13009), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1800), .B1(n13009), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12530), .COUT(n12531), .S0(n134_adj_1671), 
          .S1(n131_adj_1670));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_13 (.A0(n131_adj_1799), .B0(n13009), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1798), .B1(n13009), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12531), .COUT(n12532), .S0(n128_adj_1669), 
          .S1(n125_adj_1668));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_15 (.A0(n125_adj_1797), .B0(n13009), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1796), .B1(n13009), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12532), .COUT(n12533), .S0(n122_adj_1667), 
          .S1(n119_adj_1666));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_17 (.A0(n119_adj_1795), .B0(n13009), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1794), .B1(n13009), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12533), .COUT(n12534), .S0(n116_adj_1665), 
          .S1(n113_adj_1664));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_19 (.A0(n113_adj_1793), .B0(n13009), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1792), .B1(n13009), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12534), .COUT(n12535), .S0(n110_adj_1663), 
          .S1(n107_adj_1662));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_21 (.A0(n107_adj_1791), .B0(n13009), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1790), .B1(n13009), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12535), .COUT(n12536), .S0(n104_adj_1661), 
          .S1(n101_adj_1660));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_23 (.A0(n101_adj_1789), .B0(n13009), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1788), .B1(n13009), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12536), .COUT(n12537), .S0(n98_adj_1659), 
          .S1(n95_adj_1658));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_25 (.A0(n95_adj_1787), .B0(n13009), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1786), .B1(n13009), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12537), .COUT(n12538), .S0(n92_adj_1657), 
          .S1(n89_adj_1656));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_27 (.A0(n89_adj_1785), .B0(n13009), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1784), .B1(n13009), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12538), .COUT(n12539), .S0(n86_adj_1655), 
          .S1(n83_adj_1654));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_29 (.A0(n83_adj_1783), .B0(n13009), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1782), .B1(n13009), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12539), .COUT(n12540), .S0(n80_adj_1653), 
          .S1(n77_adj_1652));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_31 (.A0(n77_adj_1781), .B0(n13009), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1780), .B1(n13009), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12540), .COUT(n12541), .S0(n74_adj_1651), 
          .S1(n71_adj_1650));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_573_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_573_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_573_add_4_33 (.A0(n1067), .B0(n13009), .C0(n71_adj_1779), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12541), .S0(n68_adj_1649));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_573_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_573_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_573_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_573_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13009), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12542), .S1(n161_adj_1712));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_570_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_3 (.A0(n161_adj_1873), .B0(n13009), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1872), .B1(n13009), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12542), .COUT(n12543), .S0(n158_adj_1711), 
          .S1(n155_adj_1710));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_5 (.A0(n155_adj_1871), .B0(n13009), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1870), .B1(n13009), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12543), .COUT(n12544), .S0(n152_adj_1709), 
          .S1(n149_adj_1708));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_7 (.A0(n149_adj_1869), .B0(n13009), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1868), .B1(n13009), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12544), .COUT(n12545), .S0(n146_adj_1707), 
          .S1(n143_adj_1706));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_9 (.A0(n143_adj_1867), .B0(n13009), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1866), .B1(n13009), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12545), .COUT(n12546), .S0(n140_adj_1705), 
          .S1(n137_adj_1704));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_11 (.A0(n137_adj_1865), .B0(n13009), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1864), .B1(n13009), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12546), .COUT(n12547), .S0(n134_adj_1703), 
          .S1(n131_adj_1702));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_13 (.A0(n131_adj_1863), .B0(n13009), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1862), .B1(n13009), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12547), .COUT(n12548), .S0(n128_adj_1701), 
          .S1(n125_adj_1700));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_15 (.A0(n125_adj_1861), .B0(n13009), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1860), .B1(n13009), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12548), .COUT(n12549), .S0(n122_adj_1699), 
          .S1(n119_adj_1698));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_17 (.A0(n119_adj_1859), .B0(n13009), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1858), .B1(n13009), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12549), .COUT(n12550), .S0(n116_adj_1697), 
          .S1(n113_adj_1696));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_19 (.A0(n113_adj_1857), .B0(n13009), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1856), .B1(n13009), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12550), .COUT(n12551), .S0(n110_adj_1695), 
          .S1(n107_adj_1694));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_21 (.A0(n107_adj_1855), .B0(n13009), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1854), .B1(n13009), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12551), .COUT(n12552), .S0(n104_adj_1693), 
          .S1(n101_adj_1692));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_23 (.A0(n101_adj_1853), .B0(n13009), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1852), .B1(n13009), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12552), .COUT(n12553), .S0(n98_adj_1691), 
          .S1(n95_adj_1690));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_25 (.A0(n95_adj_1851), .B0(n13009), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1850), .B1(n13009), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12553), .COUT(n12554), .S0(n92_adj_1689), 
          .S1(n89_adj_1688));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_27 (.A0(n89_adj_1849), .B0(n13009), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1848), .B1(n13009), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12554), .COUT(n12555), .S0(n86_adj_1687), 
          .S1(n83_adj_1686));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_29 (.A0(n83_adj_1847), .B0(n13009), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1846), .B1(n13009), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12555), .COUT(n12556), .S0(n80_adj_1685), 
          .S1(n77_adj_1684));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_31 (.A0(n77_adj_1845), .B0(n13009), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1844), .B1(n13009), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12556), .COUT(n12557), .S0(n74_adj_1683), 
          .S1(n71_adj_1682));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_570_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_570_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_570_add_4_33 (.A0(n1067), .B0(n13009), .C0(n71_adj_1843), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12557), .S0(n68_adj_1681));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_570_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_570_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_570_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_570_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13028), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12558), .S1(n161_adj_1744));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_498_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_3 (.A0(n161_adj_2097), .B0(n13028), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_2096), .B1(n13028), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12558), .COUT(n12559), .S0(n158_adj_1743), 
          .S1(n155_adj_1742));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_5 (.A0(n155_adj_2095), .B0(n13028), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_2094), .B1(n13028), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12559), .COUT(n12560), .S0(n152_adj_1741), 
          .S1(n149_adj_1740));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_7 (.A0(n149_adj_2093), .B0(n13028), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_2092), .B1(n13028), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12560), .COUT(n12561), .S0(n146_adj_1739), 
          .S1(n143_adj_1738));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_9 (.A0(n143_adj_2091), .B0(n13028), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_2090), .B1(n13028), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12561), .COUT(n12562), .S0(n140_adj_1737), 
          .S1(n137_adj_1736));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_11 (.A0(n137_adj_2089), .B0(n13028), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_2088), .B1(n13028), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12562), .COUT(n12563), .S0(n134_adj_1735), 
          .S1(n131_adj_1734));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_13 (.A0(n131_adj_2087), .B0(n13028), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_2086), .B1(n13028), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12563), .COUT(n12564), .S0(n128_adj_1733), 
          .S1(n125_adj_1732));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_15 (.A0(n125_adj_2085), .B0(n13028), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_2084), .B1(n13028), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12564), .COUT(n12565), .S0(n122_adj_1731), 
          .S1(n119_adj_1730));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_17 (.A0(n119_adj_2083), .B0(n13028), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_2082), .B1(n13028), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12565), .COUT(n12566), .S0(n116_adj_1729), 
          .S1(n113_adj_1728));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_19 (.A0(n113_adj_2081), .B0(n13028), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_2080), .B1(n13028), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12566), .COUT(n12567), .S0(n110_adj_1727), 
          .S1(n107_adj_1726));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_21 (.A0(n107_adj_2079), .B0(n13028), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_2078), .B1(n13028), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12567), .COUT(n12568), .S0(n104_adj_1725), 
          .S1(n101_adj_1724));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_23 (.A0(n101_adj_2077), .B0(n13028), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_2076), .B1(n13028), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12568), .COUT(n12569), .S0(n98_adj_1723), 
          .S1(n95_adj_1722));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_25 (.A0(n95_adj_2075), .B0(n13028), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_2074), .B1(n13028), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12569), .COUT(n12570), .S0(n92_adj_1721), 
          .S1(n89_adj_1720));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_27 (.A0(n89_adj_2073), .B0(n13028), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_2072), .B1(n13028), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12570), .COUT(n12571), .S0(n86_adj_1719), 
          .S1(n83_adj_1718));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_29 (.A0(n83_adj_2071), .B0(n13028), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_2070), .B1(n13028), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12571), .COUT(n12572), .S0(n80_adj_1717), 
          .S1(n77_adj_1716));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_31 (.A0(n77_adj_2069), .B0(n13028), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_2068), .B1(n13028), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12572), .COUT(n12573), .S0(n74_adj_1715), 
          .S1(n71_adj_1714));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_498_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_498_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_498_add_4_33 (.A0(n1067), .B0(n13028), .C0(n71_adj_2067), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12573), .S0(n68_adj_1713));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_498_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_498_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_498_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_498_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13016), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12574), .S1(n161_adj_1776));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_429_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_3 (.A0(n161_adj_249), .B0(n13016), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_248), .B1(n13016), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12574), .COUT(n12575), .S0(n158_adj_1775), 
          .S1(n155_adj_1774));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_5 (.A0(n155_adj_247), .B0(n13016), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_246), .B1(n13016), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12575), .COUT(n12576), .S0(n152_adj_1773), 
          .S1(n149_adj_1772));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_7 (.A0(n149_adj_245), .B0(n13016), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_244), .B1(n13016), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12576), .COUT(n12577), .S0(n146_adj_1771), 
          .S1(n143_adj_1770));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_9 (.A0(n143_adj_243), .B0(n13016), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_242), .B1(n13016), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12577), .COUT(n12578), .S0(n140_adj_1769), 
          .S1(n137_adj_1768));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_11 (.A0(n137_adj_241), .B0(n13016), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_240), .B1(n13016), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12578), .COUT(n12579), .S0(n134_adj_1767), 
          .S1(n131_adj_1766));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_13 (.A0(n131_adj_239), .B0(n13016), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_238), .B1(n13016), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12579), .COUT(n12580), .S0(n128_adj_1765), 
          .S1(n125_adj_1764));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_15 (.A0(n125_adj_237), .B0(n13016), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_236), .B1(n13016), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12580), .COUT(n12581), .S0(n122_adj_1763), 
          .S1(n119_adj_1762));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_17 (.A0(n119_adj_235), .B0(n13016), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_234), .B1(n13016), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12581), .COUT(n12582), .S0(n116_adj_1761), 
          .S1(n113_adj_1760));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_19 (.A0(n113_adj_233), .B0(n13016), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_232), .B1(n13016), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12582), .COUT(n12583), .S0(n110_adj_1759), 
          .S1(n107_adj_1758));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_21 (.A0(n107_adj_231), .B0(n13016), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_230), .B1(n13016), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12583), .COUT(n12584), .S0(n104_adj_1757), 
          .S1(n101_adj_1756));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_23 (.A0(n101_adj_229), .B0(n13016), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_228), .B1(n13016), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12584), .COUT(n12585), .S0(n98_adj_1755), 
          .S1(n95_adj_1754));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_25 (.A0(n95_adj_227), .B0(n13016), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_226), .B1(n13016), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12585), .COUT(n12586), .S0(n92_adj_1753), 
          .S1(n89_adj_1752));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_27 (.A0(n89_adj_225), .B0(n13016), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_224), .B1(n13016), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12586), .COUT(n12587), .S0(n86_adj_1751), 
          .S1(n83_adj_1750));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_29 (.A0(n83_adj_223), .B0(n13016), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_222), .B1(n13016), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12587), .COUT(n12588), .S0(n80_adj_1749), 
          .S1(n77_adj_1748));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_31 (.A0(n77_adj_221), .B0(n13016), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_220), .B1(n13016), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12588), .COUT(n12589), .S0(n74_adj_1747), 
          .S1(n71_adj_1746));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_429_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_429_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_429_add_4_33 (.A0(n1067), .B0(n13016), .C0(n71_adj_219), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12589), .S0(n68_adj_1745));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_429_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_429_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_429_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_429_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_2 (.A0(n1098), .B0(det_q4_28[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n1097), .B1(n161_adj_281), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12590));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_423_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_4 (.A0(n1096), .B0(n158_adj_280), .C0(GND_net), 
          .D0(VCC_net), .A1(n1095), .B1(n155_adj_279), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12590), .COUT(n12591));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_6 (.A0(n1094), .B0(n152_adj_278), .C0(GND_net), 
          .D0(VCC_net), .A1(n1093), .B1(n149_adj_277), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12591), .COUT(n12592));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_8 (.A0(n1092), .B0(n146_adj_276), .C0(GND_net), 
          .D0(VCC_net), .A1(n1091), .B1(n143_adj_275), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12592), .COUT(n12593));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_10 (.A0(n1090), .B0(n140_adj_274), .C0(GND_net), 
          .D0(VCC_net), .A1(n1089), .B1(n137_adj_273), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12593), .COUT(n12594));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_12 (.A0(n1088), .B0(n134_adj_272), .C0(GND_net), 
          .D0(VCC_net), .A1(n1087), .B1(n131_adj_271), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12594), .COUT(n12595));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_14 (.A0(n1086), .B0(n128_adj_270), .C0(GND_net), 
          .D0(VCC_net), .A1(n1085), .B1(n125_adj_269), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12595), .COUT(n12596));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_16 (.A0(n1084), .B0(n122_adj_268), .C0(GND_net), 
          .D0(VCC_net), .A1(n1083), .B1(n119_adj_267), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12596), .COUT(n12597));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_18 (.A0(n1082), .B0(n116_adj_266), .C0(GND_net), 
          .D0(VCC_net), .A1(n1081), .B1(n113_adj_265), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12597), .COUT(n12598));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_20 (.A0(n1080), .B0(n110_adj_264), .C0(GND_net), 
          .D0(VCC_net), .A1(n1079), .B1(n107_adj_263), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12598), .COUT(n12599));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_22 (.A0(n1078), .B0(n104_adj_262), .C0(GND_net), 
          .D0(VCC_net), .A1(n1077), .B1(n101_adj_261), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12599), .COUT(n12600));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_24 (.A0(n1076), .B0(n98_adj_260), .C0(GND_net), 
          .D0(VCC_net), .A1(n1075), .B1(n95_adj_259), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12600), .COUT(n12601));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_26 (.A0(n1074), .B0(n92_adj_258), .C0(GND_net), 
          .D0(VCC_net), .A1(n1073), .B1(n89_adj_257), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12601), .COUT(n12602));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_28 (.A0(n1072), .B0(n86_adj_256), .C0(GND_net), 
          .D0(VCC_net), .A1(n1071), .B1(n83_adj_255), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12602), .COUT(n12603));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_30 (.A0(n1070), .B0(n80_adj_254), .C0(GND_net), 
          .D0(VCC_net), .A1(n1069), .B1(n77_adj_253), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12603), .COUT(n12604));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_423_add_4_32 (.A0(n1068), .B0(n74_adj_252), .C0(GND_net), 
          .D0(VCC_net), .A1(n1067), .B1(n71_adj_251), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12604), .S1(n68_adj_1777));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_423_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_423_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_423_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_423_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13010), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12606), .S1(n161_adj_1809));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_567_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_3 (.A0(n161_adj_1969), .B0(n13010), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1968), .B1(n13010), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12606), .COUT(n12607), .S0(n158_adj_1808), 
          .S1(n155_adj_1807));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_5 (.A0(n155_adj_1967), .B0(n13010), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1966), .B1(n13010), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12607), .COUT(n12608), .S0(n152_adj_1806), 
          .S1(n149_adj_1805));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_7 (.A0(n149_adj_1965), .B0(n13010), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1964), .B1(n13010), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12608), .COUT(n12609), .S0(n146_adj_1804), 
          .S1(n143_adj_1803));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_9 (.A0(n143_adj_1963), .B0(n13010), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1962), .B1(n13010), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12609), .COUT(n12610), .S0(n140_adj_1802), 
          .S1(n137_adj_1801));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_11 (.A0(n137_adj_1961), .B0(n13010), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1960), .B1(n13010), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12610), .COUT(n12611), .S0(n134_adj_1800), 
          .S1(n131_adj_1799));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_13 (.A0(n131_adj_1959), .B0(n13010), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1958), .B1(n13010), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12611), .COUT(n12612), .S0(n128_adj_1798), 
          .S1(n125_adj_1797));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_15 (.A0(n125_adj_1957), .B0(n13010), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1956), .B1(n13010), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12612), .COUT(n12613), .S0(n122_adj_1796), 
          .S1(n119_adj_1795));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_17 (.A0(n119_adj_1955), .B0(n13010), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1954), .B1(n13010), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12613), .COUT(n12614), .S0(n116_adj_1794), 
          .S1(n113_adj_1793));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_19 (.A0(n113_adj_1953), .B0(n13010), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1952), .B1(n13010), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12614), .COUT(n12615), .S0(n110_adj_1792), 
          .S1(n107_adj_1791));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_21 (.A0(n107_adj_1951), .B0(n13010), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1950), .B1(n13010), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12615), .COUT(n12616), .S0(n104_adj_1790), 
          .S1(n101_adj_1789));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_23 (.A0(n101_adj_1949), .B0(n13010), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1948), .B1(n13010), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12616), .COUT(n12617), .S0(n98_adj_1788), 
          .S1(n95_adj_1787));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_25 (.A0(n95_adj_1947), .B0(n13010), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1946), .B1(n13010), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12617), .COUT(n12618), .S0(n92_adj_1786), 
          .S1(n89_adj_1785));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_27 (.A0(n89_adj_1945), .B0(n13010), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1944), .B1(n13010), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12618), .COUT(n12619), .S0(n86_adj_1784), 
          .S1(n83_adj_1783));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_29 (.A0(n83_adj_1943), .B0(n13010), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1942), .B1(n13010), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12619), .COUT(n12620), .S0(n80_adj_1782), 
          .S1(n77_adj_1781));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_31 (.A0(n77_adj_1941), .B0(n13010), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1940), .B1(n13010), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12620), .COUT(n12621), .S0(n74_adj_1780), 
          .S1(n71_adj_1779));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_567_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_567_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_567_add_4_33 (.A0(n1067), .B0(n13010), .C0(n71_adj_1939), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12621), .S0(n68_adj_1778));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_567_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_567_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_567_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_567_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13017), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12622), .S1(n161_adj_1841));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_432_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_3 (.A0(n161_adj_1648), .B0(n13017), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1647), .B1(n13017), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12622), .COUT(n12623), .S0(n158_adj_1840), 
          .S1(n155_adj_1839));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_5 (.A0(n155_adj_1646), .B0(n13017), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1645), .B1(n13017), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12623), .COUT(n12624), .S0(n152_adj_1838), 
          .S1(n149_adj_1837));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_7 (.A0(n149_adj_1644), .B0(n13017), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1643), .B1(n13017), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12624), .COUT(n12625), .S0(n146_adj_1836), 
          .S1(n143_adj_1835));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_9 (.A0(n143_adj_1642), .B0(n13017), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1641), .B1(n13017), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12625), .COUT(n12626), .S0(n140_adj_1834), 
          .S1(n137_adj_1833));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_11 (.A0(n137_adj_1640), .B0(n13017), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1639), .B1(n13017), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12626), .COUT(n12627), .S0(n134_adj_1832), 
          .S1(n131_adj_1831));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_13 (.A0(n131_adj_1638), .B0(n13017), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1637), .B1(n13017), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12627), .COUT(n12628), .S0(n128_adj_1830), 
          .S1(n125_adj_1829));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_15 (.A0(n125_adj_1636), .B0(n13017), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1635), .B1(n13017), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12628), .COUT(n12629), .S0(n122_adj_1828), 
          .S1(n119_adj_1827));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_17 (.A0(n119_adj_1634), .B0(n13017), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1633), .B1(n13017), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12629), .COUT(n12630), .S0(n116_adj_1826), 
          .S1(n113_adj_1825));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_19 (.A0(n113_adj_1632), .B0(n13017), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1631), .B1(n13017), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12630), .COUT(n12631), .S0(n110_adj_1824), 
          .S1(n107_adj_1823));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_21 (.A0(n107_adj_1630), .B0(n13017), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1629), .B1(n13017), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12631), .COUT(n12632), .S0(n104_adj_1822), 
          .S1(n101_adj_1821));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_23 (.A0(n101_adj_1628), .B0(n13017), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1627), .B1(n13017), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12632), .COUT(n12633), .S0(n98_adj_1820), 
          .S1(n95_adj_1819));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_25 (.A0(n95_adj_1626), .B0(n13017), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1625), .B1(n13017), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12633), .COUT(n12634), .S0(n92_adj_1818), 
          .S1(n89_adj_1817));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_27 (.A0(n89_adj_1624), .B0(n13017), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1623), .B1(n13017), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12634), .COUT(n12635), .S0(n86_adj_1816), 
          .S1(n83_adj_1815));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_29 (.A0(n83_adj_1622), .B0(n13017), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1621), .B1(n13017), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12635), .COUT(n12636), .S0(n80_adj_1814), 
          .S1(n77_adj_1813));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_31 (.A0(n77_adj_1620), .B0(n13017), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1619), .B1(n13017), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12636), .COUT(n12637), .S0(n74_adj_1812), 
          .S1(n71_adj_1811));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_432_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_432_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_432_add_4_33 (.A0(n1067), .B0(n13017), .C0(n71_adj_1618), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12637), .S0(n68_adj_1810));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_432_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_432_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_432_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_432_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13010), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12638), .S1(n161_adj_1873));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_564_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_3 (.A0(n161_adj_2001), .B0(n13010), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_2000), .B1(n13010), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12638), .COUT(n12639), .S0(n158_adj_1872), 
          .S1(n155_adj_1871));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_5 (.A0(n155_adj_1999), .B0(n13010), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1998), .B1(n13010), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12639), .COUT(n12640), .S0(n152_adj_1870), 
          .S1(n149_adj_1869));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_7 (.A0(n149_adj_1997), .B0(n13010), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1996), .B1(n13010), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12640), .COUT(n12641), .S0(n146_adj_1868), 
          .S1(n143_adj_1867));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_9 (.A0(n143_adj_1995), .B0(n13010), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1994), .B1(n13010), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12641), .COUT(n12642), .S0(n140_adj_1866), 
          .S1(n137_adj_1865));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_11 (.A0(n137_adj_1993), .B0(n13010), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1992), .B1(n13010), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12642), .COUT(n12643), .S0(n134_adj_1864), 
          .S1(n131_adj_1863));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_13 (.A0(n131_adj_1991), .B0(n13010), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1990), .B1(n13010), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12643), .COUT(n12644), .S0(n128_adj_1862), 
          .S1(n125_adj_1861));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_15 (.A0(n125_adj_1989), .B0(n13010), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1988), .B1(n13010), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12644), .COUT(n12645), .S0(n122_adj_1860), 
          .S1(n119_adj_1859));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_17 (.A0(n119_adj_1987), .B0(n13010), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1986), .B1(n13010), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12645), .COUT(n12646), .S0(n116_adj_1858), 
          .S1(n113_adj_1857));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_19 (.A0(n113_adj_1985), .B0(n13010), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1984), .B1(n13010), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12646), .COUT(n12647), .S0(n110_adj_1856), 
          .S1(n107_adj_1855));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_21 (.A0(n107_adj_1983), .B0(n13010), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1982), .B1(n13010), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12647), .COUT(n12648), .S0(n104_adj_1854), 
          .S1(n101_adj_1853));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_23 (.A0(n101_adj_1981), .B0(n13010), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1980), .B1(n13010), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12648), .COUT(n12649), .S0(n98_adj_1852), 
          .S1(n95_adj_1851));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_25 (.A0(n95_adj_1979), .B0(n13010), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1978), .B1(n13010), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12649), .COUT(n12650), .S0(n92_adj_1850), 
          .S1(n89_adj_1849));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_27 (.A0(n89_adj_1977), .B0(n13010), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1976), .B1(n13010), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12650), .COUT(n12651), .S0(n86_adj_1848), 
          .S1(n83_adj_1847));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_29 (.A0(n83_adj_1975), .B0(n13010), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1974), .B1(n13010), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12651), .COUT(n12652), .S0(n80_adj_1846), 
          .S1(n77_adj_1845));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_31 (.A0(n77_adj_1973), .B0(n13010), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1972), .B1(n13010), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12652), .COUT(n12653), .S0(n74_adj_1844), 
          .S1(n71_adj_1843));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_564_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_564_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_564_add_4_33 (.A0(n1067), .B0(n13010), .C0(n71_adj_1971), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12653), .S0(n68_adj_1842));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_564_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_564_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_564_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_564_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[1]), .B1(det_q4_28[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12654), .S1(n161_adj_1905));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_495_add_4_1.INIT1 = 16'h999a;
    defparam _add_1_495_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_3 (.A0(det_q4_28[2]), .B0(n1064), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[3]), .B1(n1063), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12654), .COUT(n12655), .S0(n158_adj_1904), 
          .S1(n155_adj_1903));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_3.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_5 (.A0(det_q4_28[4]), .B0(n1062), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[5]), .B1(n1061), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12655), .COUT(n12656), .S0(n152_adj_1902), 
          .S1(n149_adj_1901));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_5.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_5.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_7 (.A0(det_q4_28[6]), .B0(n1060), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[7]), .B1(n1059), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12656), .COUT(n12657), .S0(n146_adj_1900), 
          .S1(n143_adj_1899));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_7.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_7.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_9 (.A0(det_q4_28[8]), .B0(n1058), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[9]), .B1(n1057), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12657), .COUT(n12658), .S0(n140_adj_1898), 
          .S1(n137_adj_1897));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_9.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_9.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_11 (.A0(det_q4_28[10]), .B0(n1056), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[11]), .B1(n1055), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12658), .COUT(n12659), .S0(n134_adj_1896), 
          .S1(n131_adj_1895));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_11.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_11.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_13 (.A0(det_q4_28[12]), .B0(n1054), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[13]), .B1(n1053), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12659), .COUT(n12660), .S0(n128_adj_1894), 
          .S1(n125_adj_1893));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_13.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_13.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_15 (.A0(det_q4_28[14]), .B0(n1052), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[15]), .B1(n1051), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12660), .COUT(n12661), .S0(n122_adj_1892), 
          .S1(n119_adj_1891));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_15.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_15.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_17 (.A0(det_q4_28[16]), .B0(n1050), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[17]), .B1(n1049), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12661), .COUT(n12662), .S0(n116_adj_1890), 
          .S1(n113_adj_1889));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_17.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_17.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_19 (.A0(det_q4_28[18]), .B0(n1048), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[19]), .B1(n1047), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12662), .COUT(n12663), .S0(n110_adj_1888), 
          .S1(n107_adj_1887));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_19.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_19.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_21 (.A0(det_q4_28[20]), .B0(n1046), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[21]), .B1(n1045), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12663), .COUT(n12664), .S0(n104_adj_1886), 
          .S1(n101_adj_1885));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_21.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_21.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_23 (.A0(det_q4_28[22]), .B0(n1044), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[23]), .B1(n1043), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12664), .COUT(n12665), .S0(n98_adj_1884), 
          .S1(n95_adj_1883));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_23.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_23.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_25 (.A0(det_q4_28[24]), .B0(n1042), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[25]), .B1(n1041), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12665), .COUT(n12666), .S0(n92_adj_1882), 
          .S1(n89_adj_1881));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_25.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_25.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_27 (.A0(det_q4_28[26]), .B0(n1040), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[27]), .B1(n1039), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12666), .COUT(n12667), .S0(n86_adj_1880), 
          .S1(n83_adj_1879));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_27.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_27.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_29 (.A0(det_q4_28[28]), .B0(n1038), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[29]), .B1(n1037), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12667), .COUT(n12668), .S0(n80_adj_1878), 
          .S1(n77_adj_1877));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_29.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_29.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_31 (.A0(det_q4_28[30]), .B0(n1036), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[31]), .B1(n1035), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12668), .COUT(n12669), .S0(n74_adj_1876), 
          .S1(n71_adj_1875));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_31.INIT0 = 16'h666a;
    defparam _add_1_495_add_4_31.INIT1 = 16'h666a;
    defparam _add_1_495_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_495_add_4_33 (.A0(n1034), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12669), .S0(n68_adj_1874));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_495_add_4_33.INIT0 = 16'haaa0;
    defparam _add_1_495_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_495_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_495_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13018), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12670), .S1(n161_adj_1937));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_441_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_3 (.A0(n161_adj_1553), .B0(n13018), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1552), .B1(n13018), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12670), .COUT(n12671), .S0(n158_adj_1936), 
          .S1(n155_adj_1935));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_5 (.A0(n155_adj_1551), .B0(n13018), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1550), .B1(n13018), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12671), .COUT(n12672), .S0(n152_adj_1934), 
          .S1(n149_adj_1933));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_7 (.A0(n149_adj_1549), .B0(n13018), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1548), .B1(n13018), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12672), .COUT(n12673), .S0(n146_adj_1932), 
          .S1(n143_adj_1931));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_9 (.A0(n143_adj_1547), .B0(n13018), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1546), .B1(n13018), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12673), .COUT(n12674), .S0(n140_adj_1930), 
          .S1(n137_adj_1929));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_11 (.A0(n137_adj_1545), .B0(n13018), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1544), .B1(n13018), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12674), .COUT(n12675), .S0(n134_adj_1928), 
          .S1(n131_adj_1927));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_13 (.A0(n131_adj_1543), .B0(n13018), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1542), .B1(n13018), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12675), .COUT(n12676), .S0(n128_adj_1926), 
          .S1(n125_adj_1925));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_15 (.A0(n125_adj_1541), .B0(n13018), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1540), .B1(n13018), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12676), .COUT(n12677), .S0(n122_adj_1924), 
          .S1(n119_adj_1923));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_17 (.A0(n119_adj_1539), .B0(n13018), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1538), .B1(n13018), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12677), .COUT(n12678), .S0(n116_adj_1922), 
          .S1(n113_adj_1921));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_19 (.A0(n113_adj_1537), .B0(n13018), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1536), .B1(n13018), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12678), .COUT(n12679), .S0(n110_adj_1920), 
          .S1(n107_adj_1919));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_21 (.A0(n107_adj_1535), .B0(n13018), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1534), .B1(n13018), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12679), .COUT(n12680), .S0(n104_adj_1918), 
          .S1(n101_adj_1917));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_23 (.A0(n101_adj_1533), .B0(n13018), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1532), .B1(n13018), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12680), .COUT(n12681), .S0(n98_adj_1916), 
          .S1(n95_adj_1915));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_25 (.A0(n95_adj_1531), .B0(n13018), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1530), .B1(n13018), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12681), .COUT(n12682), .S0(n92_adj_1914), 
          .S1(n89_adj_1913));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_27 (.A0(n89_adj_1529), .B0(n13018), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1528), .B1(n13018), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12682), .COUT(n12683), .S0(n86_adj_1912), 
          .S1(n83_adj_1911));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_29 (.A0(n83_adj_1527), .B0(n13018), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1526), .B1(n13018), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12683), .COUT(n12684), .S0(n80_adj_1910), 
          .S1(n77_adj_1909));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_31 (.A0(n77_adj_1525), .B0(n13018), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1524), .B1(n13018), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12684), .COUT(n12685), .S0(n74_adj_1908), 
          .S1(n71_adj_1907));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_441_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_441_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_441_add_4_33 (.A0(n1067), .B0(n13018), .C0(n71_adj_1523), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12685), .S0(n68_adj_1906));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_441_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_441_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_441_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_441_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13011), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12686), .S1(n161_adj_1969));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_561_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_3 (.A0(n161_adj_2033), .B0(n13011), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_2032), .B1(n13011), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12686), .COUT(n12687), .S0(n158_adj_1968), 
          .S1(n155_adj_1967));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_5 (.A0(n155_adj_2031), .B0(n13011), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_2030), .B1(n13011), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12687), .COUT(n12688), .S0(n152_adj_1966), 
          .S1(n149_adj_1965));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_7 (.A0(n149_adj_2029), .B0(n13011), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_2028), .B1(n13011), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12688), .COUT(n12689), .S0(n146_adj_1964), 
          .S1(n143_adj_1963));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_9 (.A0(n143_adj_2027), .B0(n13011), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_2026), .B1(n13011), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12689), .COUT(n12690), .S0(n140_adj_1962), 
          .S1(n137_adj_1961));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_11 (.A0(n137_adj_2025), .B0(n13011), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_2024), .B1(n13011), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12690), .COUT(n12691), .S0(n134_adj_1960), 
          .S1(n131_adj_1959));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_13 (.A0(n131_adj_2023), .B0(n13011), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_2022), .B1(n13011), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12691), .COUT(n12692), .S0(n128_adj_1958), 
          .S1(n125_adj_1957));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_15 (.A0(n125_adj_2021), .B0(n13011), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_2020), .B1(n13011), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12692), .COUT(n12693), .S0(n122_adj_1956), 
          .S1(n119_adj_1955));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_17 (.A0(n119_adj_2019), .B0(n13011), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_2018), .B1(n13011), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12693), .COUT(n12694), .S0(n116_adj_1954), 
          .S1(n113_adj_1953));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_19 (.A0(n113_adj_2017), .B0(n13011), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_2016), .B1(n13011), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12694), .COUT(n12695), .S0(n110_adj_1952), 
          .S1(n107_adj_1951));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_21 (.A0(n107_adj_2015), .B0(n13011), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_2014), .B1(n13011), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12695), .COUT(n12696), .S0(n104_adj_1950), 
          .S1(n101_adj_1949));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_23 (.A0(n101_adj_2013), .B0(n13011), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_2012), .B1(n13011), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12696), .COUT(n12697), .S0(n98_adj_1948), 
          .S1(n95_adj_1947));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_25 (.A0(n95_adj_2011), .B0(n13011), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_2010), .B1(n13011), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12697), .COUT(n12698), .S0(n92_adj_1946), 
          .S1(n89_adj_1945));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_27 (.A0(n89_adj_2009), .B0(n13011), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_2008), .B1(n13011), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12698), .COUT(n12699), .S0(n86_adj_1944), 
          .S1(n83_adj_1943));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_29 (.A0(n83_adj_2007), .B0(n13011), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_2006), .B1(n13011), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12699), .COUT(n12700), .S0(n80_adj_1942), 
          .S1(n77_adj_1941));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_31 (.A0(n77_adj_2005), .B0(n13011), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_2004), .B1(n13011), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12700), .COUT(n12701), .S0(n74_adj_1940), 
          .S1(n71_adj_1939));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_561_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_561_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_561_add_4_33 (.A0(n1067), .B0(n13011), .C0(n71_adj_2003), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12701), .S0(n68_adj_1938));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_561_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_561_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_561_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_561_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13011), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12702), .S1(n161_adj_2001));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_558_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_3 (.A0(n161_adj_2065), .B0(n13011), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_2064), .B1(n13011), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12702), .COUT(n12703), .S0(n158_adj_2000), 
          .S1(n155_adj_1999));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_5 (.A0(n155_adj_2063), .B0(n13011), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_2062), .B1(n13011), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12703), .COUT(n12704), .S0(n152_adj_1998), 
          .S1(n149_adj_1997));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_7 (.A0(n149_adj_2061), .B0(n13011), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_2060), .B1(n13011), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12704), .COUT(n12705), .S0(n146_adj_1996), 
          .S1(n143_adj_1995));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_9 (.A0(n143_adj_2059), .B0(n13011), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_2058), .B1(n13011), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12705), .COUT(n12706), .S0(n140_adj_1994), 
          .S1(n137_adj_1993));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_11 (.A0(n137_adj_2057), .B0(n13011), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_2056), .B1(n13011), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12706), .COUT(n12707), .S0(n134_adj_1992), 
          .S1(n131_adj_1991));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_13 (.A0(n131_adj_2055), .B0(n13011), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_2054), .B1(n13011), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12707), .COUT(n12708), .S0(n128_adj_1990), 
          .S1(n125_adj_1989));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_15 (.A0(n125_adj_2053), .B0(n13011), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_2052), .B1(n13011), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12708), .COUT(n12709), .S0(n122_adj_1988), 
          .S1(n119_adj_1987));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_17 (.A0(n119_adj_2051), .B0(n13011), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_2050), .B1(n13011), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12709), .COUT(n12710), .S0(n116_adj_1986), 
          .S1(n113_adj_1985));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_19 (.A0(n113_adj_2049), .B0(n13011), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_2048), .B1(n13011), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12710), .COUT(n12711), .S0(n110_adj_1984), 
          .S1(n107_adj_1983));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_21 (.A0(n107_adj_2047), .B0(n13011), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_2046), .B1(n13011), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12711), .COUT(n12712), .S0(n104_adj_1982), 
          .S1(n101_adj_1981));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_23 (.A0(n101_adj_2045), .B0(n13011), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_2044), .B1(n13011), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12712), .COUT(n12713), .S0(n98_adj_1980), 
          .S1(n95_adj_1979));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_25 (.A0(n95_adj_2043), .B0(n13011), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_2042), .B1(n13011), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12713), .COUT(n12714), .S0(n92_adj_1978), 
          .S1(n89_adj_1977));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_27 (.A0(n89_adj_2041), .B0(n13011), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_2040), .B1(n13011), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12714), .COUT(n12715), .S0(n86_adj_1976), 
          .S1(n83_adj_1975));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_29 (.A0(n83_adj_2039), .B0(n13011), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_2038), .B1(n13011), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12715), .COUT(n12716), .S0(n80_adj_1974), 
          .S1(n77_adj_1973));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_31 (.A0(n77_adj_2037), .B0(n13011), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_2036), .B1(n13011), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12716), .COUT(n12717), .S0(n74_adj_1972), 
          .S1(n71_adj_1971));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_558_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_558_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_558_add_4_33 (.A0(n1067), .B0(n13011), .C0(n71_adj_2035), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12717), .S0(n68_adj_1970));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_558_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_558_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_558_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_558_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[1]), .B1(det_q4_28[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12718), .S1(n1098));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_492_add_4_1.INIT1 = 16'h6665;
    defparam _add_1_492_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_3 (.A0(det_q4_28[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12718), .COUT(n12719), .S0(n1097), .S1(n1096));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_5 (.A0(det_q4_28[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12719), .COUT(n12720), .S0(n1095), .S1(n1094));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_7 (.A0(det_q4_28[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12720), .COUT(n12721), .S0(n1093), .S1(n1092));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_9 (.A0(det_q4_28[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12721), .COUT(n12722), .S0(n1091), .S1(n1090));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_11 (.A0(det_q4_28[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12722), .COUT(n12723), .S0(n1089), .S1(n1088));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_13 (.A0(det_q4_28[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12723), .COUT(n12724), .S0(n1087), .S1(n1086));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_13.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_15 (.A0(det_q4_28[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12724), .COUT(n12725), .S0(n1085), .S1(n1084));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_15.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_15.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_17 (.A0(det_q4_28[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12725), .COUT(n12726), .S0(n1083), .S1(n1082));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_17.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_17.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_19 (.A0(det_q4_28[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12726), .COUT(n12727), .S0(n1081), .S1(n1080));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_19.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_19.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_21 (.A0(det_q4_28[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12727), .COUT(n12728), .S0(n1079), .S1(n1078));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_21.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_21.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_23 (.A0(det_q4_28[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12728), .COUT(n12729), .S0(n1077), .S1(n1076));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_23.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_23.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_25 (.A0(det_q4_28[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12729), .COUT(n12730), .S0(n1075), .S1(n1074));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_25.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_25.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_27 (.A0(det_q4_28[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12730), .COUT(n12731), .S0(n1073), .S1(n1072));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_27.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_27.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_29 (.A0(det_q4_28[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12731), .COUT(n12732), .S0(n1071), .S1(n1070));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_29.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_29.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_31 (.A0(det_q4_28[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12732), .COUT(n12733), .S0(n1069), .S1(n1068));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_31.INIT0 = 16'h5555;
    defparam _add_1_492_add_4_31.INIT1 = 16'h5555;
    defparam _add_1_492_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_492_add_4_33 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12733), .S0(n1067));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_492_add_4_33.INIT0 = 16'hffff;
    defparam _add_1_492_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_492_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_492_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n12734), .S1(b_s[0]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_411_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_411_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_3 (.A0(b_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12734), .COUT(n12735), .S0(b_s[1]), .S1(b_s[2]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_5 (.A0(b_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12735), .COUT(n12736), .S0(b_s[3]), .S1(b_s[4]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_7 (.A0(b_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12736), .COUT(n12737), .S0(b_s[5]), .S1(b_s[6]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_9 (.A0(b_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n12737), .COUT(n12738), .S0(b_s[7]), .S1(b_s[8]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_11 (.A0(b_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12738), .COUT(n12739), .S0(b_s[9]), .S1(b_s[10]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_13 (.A0(b_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12739), .COUT(n12740), .S0(b_s[11]), .S1(b_s[12]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_13.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_15 (.A0(b_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12740), .COUT(n12741), .S0(b_s[13]), .S1(b_s[14]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_15.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_15.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_411_add_4_17 (.A0(b_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(b_reg[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n12741), .S0(b_s[15]), .S1(b_s[16]));   // d:/rtl_fpga/projeto_final/inverter/inverter.v(79[30:58])
    defparam _add_1_411_add_4_17.INIT0 = 16'h5555;
    defparam _add_1_411_add_4_17.INIT1 = 16'h5555;
    defparam _add_1_411_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_411_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13012), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12743), .S1(n161_adj_2033));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_555_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_3 (.A0(n161_adj_663), .B0(n13012), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_662), .B1(n13012), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12743), .COUT(n12744), .S0(n158_adj_2032), 
          .S1(n155_adj_2031));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_5 (.A0(n155_adj_661), .B0(n13012), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_660), .B1(n13012), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12744), .COUT(n12745), .S0(n152_adj_2030), 
          .S1(n149_adj_2029));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_7 (.A0(n149_adj_659), .B0(n13012), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_658), .B1(n13012), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12745), .COUT(n12746), .S0(n146_adj_2028), 
          .S1(n143_adj_2027));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_9 (.A0(n143_adj_657), .B0(n13012), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_656), .B1(n13012), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12746), .COUT(n12747), .S0(n140_adj_2026), 
          .S1(n137_adj_2025));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_11 (.A0(n137_adj_655), .B0(n13012), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_654), .B1(n13012), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12747), .COUT(n12748), .S0(n134_adj_2024), 
          .S1(n131_adj_2023));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_13 (.A0(n131_adj_653), .B0(n13012), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_652), .B1(n13012), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12748), .COUT(n12749), .S0(n128_adj_2022), 
          .S1(n125_adj_2021));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_15 (.A0(n125_adj_651), .B0(n13012), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_650), .B1(n13012), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12749), .COUT(n12750), .S0(n122_adj_2020), 
          .S1(n119_adj_2019));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_17 (.A0(n119_adj_649), .B0(n13012), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_648), .B1(n13012), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12750), .COUT(n12751), .S0(n116_adj_2018), 
          .S1(n113_adj_2017));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_19 (.A0(n113_adj_647), .B0(n13012), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_646), .B1(n13012), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12751), .COUT(n12752), .S0(n110_adj_2016), 
          .S1(n107_adj_2015));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_21 (.A0(n107_adj_645), .B0(n13012), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_644), .B1(n13012), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12752), .COUT(n12753), .S0(n104_adj_2014), 
          .S1(n101_adj_2013));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_23 (.A0(n101_adj_643), .B0(n13012), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_642), .B1(n13012), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12753), .COUT(n12754), .S0(n98_adj_2012), 
          .S1(n95_adj_2011));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_25 (.A0(n95_adj_641), .B0(n13012), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_640), .B1(n13012), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12754), .COUT(n12755), .S0(n92_adj_2010), 
          .S1(n89_adj_2009));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_27 (.A0(n89_adj_639), .B0(n13012), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_638), .B1(n13012), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12755), .COUT(n12756), .S0(n86_adj_2008), 
          .S1(n83_adj_2007));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_29 (.A0(n83_adj_637), .B0(n13012), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_636), .B1(n13012), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12756), .COUT(n12757), .S0(n80_adj_2006), 
          .S1(n77_adj_2005));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_31 (.A0(n77_adj_635), .B0(n13012), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_634), .B1(n13012), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12757), .COUT(n12758), .S0(n74_adj_2004), 
          .S1(n71_adj_2003));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_555_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_555_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_555_add_4_33 (.A0(n1067), .B0(n13012), .C0(n71_adj_633), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12758), .S0(n68_adj_2002));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_555_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_555_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_555_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_555_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13012), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12759), .S1(n161_adj_2065));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_552_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_3 (.A0(n161_adj_695), .B0(n13012), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_694), .B1(n13012), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12759), .COUT(n12760), .S0(n158_adj_2064), 
          .S1(n155_adj_2063));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_5 (.A0(n155_adj_693), .B0(n13012), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_692), .B1(n13012), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12760), .COUT(n12761), .S0(n152_adj_2062), 
          .S1(n149_adj_2061));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_7 (.A0(n149_adj_691), .B0(n13012), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_690), .B1(n13012), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12761), .COUT(n12762), .S0(n146_adj_2060), 
          .S1(n143_adj_2059));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_9 (.A0(n143_adj_689), .B0(n13012), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_688), .B1(n13012), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12762), .COUT(n12763), .S0(n140_adj_2058), 
          .S1(n137_adj_2057));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_11 (.A0(n137_adj_687), .B0(n13012), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_686), .B1(n13012), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12763), .COUT(n12764), .S0(n134_adj_2056), 
          .S1(n131_adj_2055));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_13 (.A0(n131_adj_685), .B0(n13012), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_684), .B1(n13012), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12764), .COUT(n12765), .S0(n128_adj_2054), 
          .S1(n125_adj_2053));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_15 (.A0(n125_adj_683), .B0(n13012), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_682), .B1(n13012), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12765), .COUT(n12766), .S0(n122_adj_2052), 
          .S1(n119_adj_2051));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_17 (.A0(n119_adj_681), .B0(n13012), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_680), .B1(n13012), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12766), .COUT(n12767), .S0(n116_adj_2050), 
          .S1(n113_adj_2049));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_19 (.A0(n113_adj_679), .B0(n13012), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_678), .B1(n13012), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12767), .COUT(n12768), .S0(n110_adj_2048), 
          .S1(n107_adj_2047));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_21 (.A0(n107_adj_677), .B0(n13012), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_676), .B1(n13012), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12768), .COUT(n12769), .S0(n104_adj_2046), 
          .S1(n101_adj_2045));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_23 (.A0(n101_adj_675), .B0(n13012), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_674), .B1(n13012), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12769), .COUT(n12770), .S0(n98_adj_2044), 
          .S1(n95_adj_2043));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_25 (.A0(n95_adj_673), .B0(n13012), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_672), .B1(n13012), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12770), .COUT(n12771), .S0(n92_adj_2042), 
          .S1(n89_adj_2041));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_27 (.A0(n89_adj_671), .B0(n13012), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_670), .B1(n13012), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12771), .COUT(n12772), .S0(n86_adj_2040), 
          .S1(n83_adj_2039));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_29 (.A0(n83_adj_669), .B0(n13012), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_668), .B1(n13012), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12772), .COUT(n12773), .S0(n80_adj_2038), 
          .S1(n77_adj_2037));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_31 (.A0(n77_adj_667), .B0(n13012), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_666), .B1(n13012), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12773), .COUT(n12774), .S0(n74_adj_2036), 
          .S1(n71_adj_2035));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_552_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_552_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_552_add_4_33 (.A0(n1067), .B0(n13012), .C0(n71_adj_665), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12774), .S0(n68_adj_2034));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_552_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_552_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_552_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_552_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n1098), .B1(det_q4_28[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n12775), .S1(n161_adj_2097));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_414_add_4_1.INIT1 = 16'h999a;
    defparam _add_1_414_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_3 (.A0(n1097), .B0(n1064), .C0(GND_net), .D0(VCC_net), 
          .A1(n1096), .B1(n1063), .C1(GND_net), .D1(VCC_net), .CIN(n12775), 
          .COUT(n12776), .S0(n158_adj_2096), .S1(n155_adj_2095));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_3.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_5 (.A0(n1095), .B0(n1062), .C0(GND_net), .D0(VCC_net), 
          .A1(n1094), .B1(n1061), .C1(GND_net), .D1(VCC_net), .CIN(n12776), 
          .COUT(n12777), .S0(n152_adj_2094), .S1(n149_adj_2093));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_5.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_5.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_7 (.A0(n1093), .B0(n1060), .C0(GND_net), .D0(VCC_net), 
          .A1(n1092), .B1(n1059), .C1(GND_net), .D1(VCC_net), .CIN(n12777), 
          .COUT(n12778), .S0(n146_adj_2092), .S1(n143_adj_2091));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_7.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_7.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_9 (.A0(n1091), .B0(n1058), .C0(GND_net), .D0(VCC_net), 
          .A1(n1090), .B1(n1057), .C1(GND_net), .D1(VCC_net), .CIN(n12778), 
          .COUT(n12779), .S0(n140_adj_2090), .S1(n137_adj_2089));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_9.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_9.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_11 (.A0(n1089), .B0(n1056), .C0(GND_net), .D0(VCC_net), 
          .A1(n1088), .B1(n1055), .C1(GND_net), .D1(VCC_net), .CIN(n12779), 
          .COUT(n12780), .S0(n134_adj_2088), .S1(n131_adj_2087));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_11.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_11.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_13 (.A0(n1087), .B0(n1054), .C0(GND_net), .D0(VCC_net), 
          .A1(n1086), .B1(n1053), .C1(GND_net), .D1(VCC_net), .CIN(n12780), 
          .COUT(n12781), .S0(n128_adj_2086), .S1(n125_adj_2085));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_13.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_13.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_15 (.A0(n1085), .B0(n1052), .C0(GND_net), .D0(VCC_net), 
          .A1(n1084), .B1(n1051), .C1(GND_net), .D1(VCC_net), .CIN(n12781), 
          .COUT(n12782), .S0(n122_adj_2084), .S1(n119_adj_2083));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_15.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_15.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_17 (.A0(n1083), .B0(n1050), .C0(GND_net), .D0(VCC_net), 
          .A1(n1082), .B1(n1049), .C1(GND_net), .D1(VCC_net), .CIN(n12782), 
          .COUT(n12783), .S0(n116_adj_2082), .S1(n113_adj_2081));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_17.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_17.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_19 (.A0(n1081), .B0(n1048), .C0(GND_net), .D0(VCC_net), 
          .A1(n1080), .B1(n1047), .C1(GND_net), .D1(VCC_net), .CIN(n12783), 
          .COUT(n12784), .S0(n110_adj_2080), .S1(n107_adj_2079));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_19.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_19.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_21 (.A0(n1079), .B0(n1046), .C0(GND_net), .D0(VCC_net), 
          .A1(n1078), .B1(n1045), .C1(GND_net), .D1(VCC_net), .CIN(n12784), 
          .COUT(n12785), .S0(n104_adj_2078), .S1(n101_adj_2077));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_21.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_21.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_23 (.A0(n1077), .B0(n1044), .C0(GND_net), .D0(VCC_net), 
          .A1(n1076), .B1(n1043), .C1(GND_net), .D1(VCC_net), .CIN(n12785), 
          .COUT(n12786), .S0(n98_adj_2076), .S1(n95_adj_2075));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_23.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_23.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_25 (.A0(n1075), .B0(n1042), .C0(GND_net), .D0(VCC_net), 
          .A1(n1074), .B1(n1041), .C1(GND_net), .D1(VCC_net), .CIN(n12786), 
          .COUT(n12787), .S0(n92_adj_2074), .S1(n89_adj_2073));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_25.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_25.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_27 (.A0(n1073), .B0(n1040), .C0(GND_net), .D0(VCC_net), 
          .A1(n1072), .B1(n1039), .C1(GND_net), .D1(VCC_net), .CIN(n12787), 
          .COUT(n12788), .S0(n86_adj_2072), .S1(n83_adj_2071));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_27.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_27.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_29 (.A0(n1071), .B0(n1038), .C0(GND_net), .D0(VCC_net), 
          .A1(n1070), .B1(n1037), .C1(GND_net), .D1(VCC_net), .CIN(n12788), 
          .COUT(n12789), .S0(n80_adj_2070), .S1(n77_adj_2069));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_29.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_29.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_31 (.A0(n1069), .B0(n1036), .C0(GND_net), .D0(VCC_net), 
          .A1(n1068), .B1(n1035), .C1(GND_net), .D1(VCC_net), .CIN(n12789), 
          .COUT(n12790), .S0(n74_adj_2068), .S1(n71_adj_2067));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_31.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_31.INIT1 = 16'h666a;
    defparam _add_1_414_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_414_add_4_33 (.A0(n1067), .B0(n1034), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12790), 
          .S0(n68_adj_2066));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_414_add_4_33.INIT0 = 16'h666a;
    defparam _add_1_414_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_414_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_414_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(det_q4_28[0]), .B1(n13019), .C1(det_q4_28[1]), 
          .D1(n1098), .COUT(n12791), .S1(n161_adj_2129));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_444_add_4_1.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_3 (.A0(n161_adj_1521), .B0(n13019), .C0(det_q4_28[2]), 
          .D0(n1097), .A1(n158_adj_1520), .B1(n13019), .C1(det_q4_28[3]), 
          .D1(n1096), .CIN(n12791), .COUT(n12792), .S0(n158_adj_2128), 
          .S1(n155_adj_2127));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_3.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_5 (.A0(n155_adj_1519), .B0(n13019), .C0(det_q4_28[4]), 
          .D0(n1095), .A1(n152_adj_1518), .B1(n13019), .C1(det_q4_28[5]), 
          .D1(n1094), .CIN(n12792), .COUT(n12793), .S0(n152_adj_2126), 
          .S1(n149_adj_2125));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_7 (.A0(n149_adj_1517), .B0(n13019), .C0(det_q4_28[6]), 
          .D0(n1093), .A1(n146_adj_1516), .B1(n13019), .C1(det_q4_28[7]), 
          .D1(n1092), .CIN(n12793), .COUT(n12794), .S0(n146_adj_2124), 
          .S1(n143_adj_2123));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_9 (.A0(n143_adj_1515), .B0(n13019), .C0(det_q4_28[8]), 
          .D0(n1091), .A1(n140_adj_1514), .B1(n13019), .C1(det_q4_28[9]), 
          .D1(n1090), .CIN(n12794), .COUT(n12795), .S0(n140_adj_2122), 
          .S1(n137_adj_2121));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_11 (.A0(n137_adj_1513), .B0(n13019), .C0(det_q4_28[10]), 
          .D0(n1089), .A1(n134_adj_1512), .B1(n13019), .C1(det_q4_28[11]), 
          .D1(n1088), .CIN(n12795), .COUT(n12796), .S0(n134_adj_2120), 
          .S1(n131_adj_2119));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_13 (.A0(n131_adj_1511), .B0(n13019), .C0(det_q4_28[12]), 
          .D0(n1087), .A1(n128_adj_1510), .B1(n13019), .C1(det_q4_28[13]), 
          .D1(n1086), .CIN(n12796), .COUT(n12797), .S0(n128_adj_2118), 
          .S1(n125_adj_2117));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_13.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_13.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_15 (.A0(n125_adj_1509), .B0(n13019), .C0(det_q4_28[14]), 
          .D0(n1085), .A1(n122_adj_1508), .B1(n13019), .C1(det_q4_28[15]), 
          .D1(n1084), .CIN(n12797), .COUT(n12798), .S0(n122_adj_2116), 
          .S1(n119_adj_2115));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_15.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_15.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_17 (.A0(n119_adj_1507), .B0(n13019), .C0(det_q4_28[16]), 
          .D0(n1083), .A1(n116_adj_1506), .B1(n13019), .C1(det_q4_28[17]), 
          .D1(n1082), .CIN(n12798), .COUT(n12799), .S0(n116_adj_2114), 
          .S1(n113_adj_2113));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_17.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_17.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_19 (.A0(n113_adj_1505), .B0(n13019), .C0(det_q4_28[18]), 
          .D0(n1081), .A1(n110_adj_1504), .B1(n13019), .C1(det_q4_28[19]), 
          .D1(n1080), .CIN(n12799), .COUT(n12800), .S0(n110_adj_2112), 
          .S1(n107_adj_2111));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_19.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_19.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_21 (.A0(n107_adj_1503), .B0(n13019), .C0(det_q4_28[20]), 
          .D0(n1079), .A1(n104_adj_1502), .B1(n13019), .C1(det_q4_28[21]), 
          .D1(n1078), .CIN(n12800), .COUT(n12801), .S0(n104_adj_2110), 
          .S1(n101_adj_2109));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_21.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_21.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_23 (.A0(n101_adj_1501), .B0(n13019), .C0(det_q4_28[22]), 
          .D0(n1077), .A1(n98_adj_1500), .B1(n13019), .C1(det_q4_28[23]), 
          .D1(n1076), .CIN(n12801), .COUT(n12802), .S0(n98_adj_2108), 
          .S1(n95_adj_2107));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_23.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_23.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_25 (.A0(n95_adj_1499), .B0(n13019), .C0(det_q4_28[24]), 
          .D0(n1075), .A1(n92_adj_1498), .B1(n13019), .C1(det_q4_28[25]), 
          .D1(n1074), .CIN(n12802), .COUT(n12803), .S0(n92_adj_2106), 
          .S1(n89_adj_2105));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_25.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_25.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_27 (.A0(n89_adj_1497), .B0(n13019), .C0(det_q4_28[26]), 
          .D0(n1073), .A1(n86_adj_1496), .B1(n13019), .C1(det_q4_28[27]), 
          .D1(n1072), .CIN(n12803), .COUT(n12804), .S0(n86_adj_2104), 
          .S1(n83_adj_2103));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_27.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_27.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_29 (.A0(n83_adj_1495), .B0(n13019), .C0(det_q4_28[28]), 
          .D0(n1071), .A1(n80_adj_1494), .B1(n13019), .C1(det_q4_28[29]), 
          .D1(n1070), .CIN(n12804), .COUT(n12805), .S0(n80_adj_2102), 
          .S1(n77_adj_2101));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_29.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_29.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_31 (.A0(n77_adj_1493), .B0(n13019), .C0(det_q4_28[30]), 
          .D0(n1069), .A1(n74_adj_1492), .B1(n13019), .C1(det_q4_28[31]), 
          .D1(n1068), .CIN(n12805), .COUT(n12806), .S0(n74_adj_2100), 
          .S1(n71_adj_2099));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_31.INIT0 = 16'h596a;
    defparam _add_1_444_add_4_31.INIT1 = 16'h596a;
    defparam _add_1_444_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_444_add_4_33 (.A0(n1067), .B0(n13019), .C0(n71_adj_1491), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12806), .S0(n68_adj_2098));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam _add_1_444_add_4_33.INIT0 = 16'hd2d2;
    defparam _add_1_444_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_444_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_444_add_4_33.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module reciprocal_q16_16
//

module reciprocal_q16_16 (error_recip, clk_c, det_zero, n1081, det_q4_28, 
            n13023, n1517, n1080, n1516, n1079, n1515, n1078, 
            n1514, n1077, n1513, n1076, n1512, n1075, n1511, n1092, 
            n13016, n2064, n1091, n2063, n1074, n1510, n1073, 
            n1509, n1072, n1508, n1071, n1507, n1070, n1506, n1090, 
            n2062, n1069, n1505, n1068, n1504, n1098, n2070, n1097, 
            n2069, n1089, n2061, n1096, n2068, n1095, n2067, n1094, 
            n2066, n1088, n2060, n1087, n2059, n1086, n2058, n1085, 
            n2057, n1084, n2056, n1083, n2055, n1082, n2054, n2053, 
            n2052, n2051, n2050, n2049, n2048, n2047, n2046, n2045, 
            n2044, n2043, n2042, n2041, n2040, n1093, n2065, n3077, 
            n3110, n1067, n13015, n2241, n2243, n2242, n2245, 
            n2244, n2247, n2246, n2249, n2248, n2251, n2250, n2253, 
            n2252, n2255, n2254, n2257, n2256, n2259, n2258, n2261, 
            n2260, n2263, n2262, n2265, n2264, n2267, n2266, n2269, 
            n2268, n2271, n2270, n13004, n3075, n3074, n3073, 
            n3072, n3071, n3070, n3069, n3068, n3067, n3066, n3065, 
            n3064, n3063, n3062, n3061, n3060, n3059, n3058, n3057, 
            n3056, n3055, n3054, n3053, n3052, n3051, n3050, n3049, 
            n3048, n1536, n39, n68, n68_adj_1, n68_adj_2, n64, 
            n63, n62, n3047, n3046, n3045, n1534, n1533, n1532, 
            n1531, n1530, n1529, n1528, n1527, n1526, n1525, n1524, 
            n1523, n1522, n1521, n2273, n50, n2139, n48, n2072, 
            n47, GND_net, n1520, n1519, n1518, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output error_recip;
    input clk_c;
    output det_zero;
    input n1081;
    input [31:0]det_q4_28;
    input n13023;
    output n1517;
    input n1080;
    output n1516;
    input n1079;
    output n1515;
    input n1078;
    output n1514;
    input n1077;
    output n1513;
    input n1076;
    output n1512;
    input n1075;
    output n1511;
    input n1092;
    input n13016;
    output n2064;
    input n1091;
    output n2063;
    input n1074;
    output n1510;
    input n1073;
    output n1509;
    input n1072;
    output n1508;
    input n1071;
    output n1507;
    input n1070;
    output n1506;
    input n1090;
    output n2062;
    input n1069;
    output n1505;
    input n1068;
    output n1504;
    input n1098;
    output n2070;
    input n1097;
    output n2069;
    input n1089;
    output n2061;
    input n1096;
    output n2068;
    input n1095;
    output n2067;
    input n1094;
    output n2066;
    input n1088;
    output n2060;
    input n1087;
    output n2059;
    input n1086;
    output n2058;
    input n1085;
    output n2057;
    input n1084;
    output n2056;
    input n1083;
    output n2055;
    input n1082;
    output n2054;
    output n2053;
    output n2052;
    output n2051;
    output n2050;
    output n2049;
    output n2048;
    output n2047;
    output n2046;
    output n2045;
    output n2044;
    output n2043;
    output n2042;
    output n2041;
    output n2040;
    input n1093;
    output n2065;
    input n3077;
    output [31:0]n3110;
    input n1067;
    input n13015;
    output n2241;
    output n2243;
    output n2242;
    output n2245;
    output n2244;
    output n2247;
    output n2246;
    output n2249;
    output n2248;
    output n2251;
    output n2250;
    output n2253;
    output n2252;
    output n2255;
    output n2254;
    output n2257;
    output n2256;
    output n2259;
    output n2258;
    output n2261;
    output n2260;
    output n2263;
    output n2262;
    output n2265;
    output n2264;
    output n2267;
    output n2266;
    output n2269;
    output n2268;
    output n2271;
    output n2270;
    input n13004;
    output n3075;
    output n3074;
    output n3073;
    output n3072;
    output n3071;
    output n3070;
    output n3069;
    output n3068;
    output n3067;
    output n3066;
    output n3065;
    output n3064;
    output n3063;
    output n3062;
    output n3061;
    output n3060;
    output n3059;
    output n3058;
    output n3057;
    output n3056;
    output n3055;
    output n3054;
    output n3053;
    output n3052;
    output n3051;
    output n3050;
    output n3049;
    output n3048;
    input n1536;
    output n39;
    input n68;
    input n68_adj_1;
    input n68_adj_2;
    output n64;
    output n63;
    output n62;
    output n3047;
    output n3046;
    output n3045;
    output n1534;
    output n1533;
    output n1532;
    output n1531;
    output n1530;
    output n1529;
    output n1528;
    output n1527;
    output n1526;
    output n1525;
    output n1524;
    output n1523;
    output n1522;
    output n1521;
    input n2273;
    output n50;
    input n2139;
    output n48;
    input n2072;
    output n47;
    input GND_net;
    output n1520;
    output n1519;
    output n1518;
    input VCC_net;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // d:/rtl_fpga/projeto_final/inverter/inverter.v(16[20:23])
    
    wire n12843, n12842, n12841, n12840;
    
    FD1S3AX error_10 (.D(det_zero), .CK(clk_c), .Q(error_recip)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=23, LSE_RCOL=6, LSE_LLINE=61, LSE_RLINE=67 */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(24[18] 31[12])
    defparam error_10.GSR = "ENABLED";
    LUT4 mux_51_i18_3_lut (.A(n1081), .B(det_q4_28[18]), .C(n13023), .Z(n1517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i18_3_lut.init = 16'hcaca;
    LUT4 mux_51_i19_3_lut (.A(n1080), .B(det_q4_28[19]), .C(n13023), .Z(n1516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i19_3_lut.init = 16'hcaca;
    LUT4 mux_51_i20_3_lut (.A(n1079), .B(det_q4_28[20]), .C(n13023), .Z(n1515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i20_3_lut.init = 16'hcaca;
    LUT4 mux_51_i21_3_lut (.A(n1078), .B(det_q4_28[21]), .C(n13023), .Z(n1514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i21_3_lut.init = 16'hcaca;
    LUT4 mux_51_i22_3_lut (.A(n1077), .B(det_q4_28[22]), .C(n13023), .Z(n1513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i22_3_lut.init = 16'hcaca;
    LUT4 mux_51_i23_3_lut (.A(n1076), .B(det_q4_28[23]), .C(n13023), .Z(n1512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i23_3_lut.init = 16'hcaca;
    LUT4 mux_51_i24_3_lut (.A(n1075), .B(det_q4_28[24]), .C(n13023), .Z(n1511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i24_3_lut.init = 16'hcaca;
    LUT4 mux_67_i7_3_lut (.A(n1092), .B(det_q4_28[7]), .C(n13016), .Z(n2064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i7_3_lut.init = 16'hcaca;
    LUT4 mux_67_i8_3_lut (.A(n1091), .B(det_q4_28[8]), .C(n13016), .Z(n2063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i8_3_lut.init = 16'hcaca;
    LUT4 mux_51_i25_3_lut (.A(n1074), .B(det_q4_28[25]), .C(n13023), .Z(n1510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i25_3_lut.init = 16'hcaca;
    LUT4 mux_51_i26_3_lut (.A(n1073), .B(det_q4_28[26]), .C(n13023), .Z(n1509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i26_3_lut.init = 16'hcaca;
    LUT4 mux_51_i27_3_lut (.A(n1072), .B(det_q4_28[27]), .C(n13023), .Z(n1508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i27_3_lut.init = 16'hcaca;
    LUT4 mux_51_i28_3_lut (.A(n1071), .B(det_q4_28[28]), .C(n13023), .Z(n1507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i28_3_lut.init = 16'hcaca;
    LUT4 mux_51_i29_3_lut (.A(n1070), .B(det_q4_28[29]), .C(n13023), .Z(n1506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i29_3_lut.init = 16'hcaca;
    LUT4 mux_67_i9_3_lut (.A(n1090), .B(det_q4_28[9]), .C(n13016), .Z(n2062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i9_3_lut.init = 16'hcaca;
    LUT4 mux_51_i30_3_lut (.A(n1069), .B(det_q4_28[30]), .C(n13023), .Z(n1505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i30_3_lut.init = 16'hcaca;
    LUT4 mux_51_i31_3_lut (.A(n1068), .B(det_q4_28[31]), .C(n13023), .Z(n1504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i31_3_lut.init = 16'hcaca;
    LUT4 mux_67_i1_3_lut (.A(n1098), .B(det_q4_28[1]), .C(n13016), .Z(n2070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i1_3_lut.init = 16'hcaca;
    LUT4 mux_67_i2_3_lut (.A(n1097), .B(det_q4_28[2]), .C(n13016), .Z(n2069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i2_3_lut.init = 16'hcaca;
    LUT4 mux_67_i10_3_lut (.A(n1089), .B(det_q4_28[10]), .C(n13016), .Z(n2061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i10_3_lut.init = 16'hcaca;
    LUT4 mux_67_i3_3_lut (.A(n1096), .B(det_q4_28[3]), .C(n13016), .Z(n2068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i3_3_lut.init = 16'hcaca;
    LUT4 mux_67_i4_3_lut (.A(n1095), .B(det_q4_28[4]), .C(n13016), .Z(n2067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i4_3_lut.init = 16'hcaca;
    LUT4 mux_67_i5_3_lut (.A(n1094), .B(det_q4_28[5]), .C(n13016), .Z(n2066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i5_3_lut.init = 16'hcaca;
    LUT4 mux_67_i11_3_lut (.A(n1088), .B(det_q4_28[11]), .C(n13016), .Z(n2060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i11_3_lut.init = 16'hcaca;
    LUT4 mux_67_i12_3_lut (.A(n1087), .B(det_q4_28[12]), .C(n13016), .Z(n2059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i12_3_lut.init = 16'hcaca;
    LUT4 mux_67_i13_3_lut (.A(n1086), .B(det_q4_28[13]), .C(n13016), .Z(n2058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i13_3_lut.init = 16'hcaca;
    LUT4 mux_67_i14_3_lut (.A(n1085), .B(det_q4_28[14]), .C(n13016), .Z(n2057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i14_3_lut.init = 16'hcaca;
    LUT4 mux_67_i15_3_lut (.A(n1084), .B(det_q4_28[15]), .C(n13016), .Z(n2056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i15_3_lut.init = 16'hcaca;
    LUT4 mux_67_i16_3_lut (.A(n1083), .B(det_q4_28[16]), .C(n13016), .Z(n2055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i16_3_lut.init = 16'hcaca;
    LUT4 mux_67_i17_3_lut (.A(n1082), .B(det_q4_28[17]), .C(n13016), .Z(n2054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i17_3_lut.init = 16'hcaca;
    LUT4 mux_67_i18_3_lut (.A(n1081), .B(det_q4_28[18]), .C(n13016), .Z(n2053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i18_3_lut.init = 16'hcaca;
    LUT4 mux_67_i19_3_lut (.A(n1080), .B(det_q4_28[19]), .C(n13016), .Z(n2052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i19_3_lut.init = 16'hcaca;
    LUT4 mux_67_i20_3_lut (.A(n1079), .B(det_q4_28[20]), .C(n13016), .Z(n2051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i20_3_lut.init = 16'hcaca;
    LUT4 mux_67_i21_3_lut (.A(n1078), .B(det_q4_28[21]), .C(n13016), .Z(n2050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i21_3_lut.init = 16'hcaca;
    LUT4 mux_67_i22_3_lut (.A(n1077), .B(det_q4_28[22]), .C(n13016), .Z(n2049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i22_3_lut.init = 16'hcaca;
    LUT4 mux_67_i23_3_lut (.A(n1076), .B(det_q4_28[23]), .C(n13016), .Z(n2048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i23_3_lut.init = 16'hcaca;
    LUT4 mux_67_i24_3_lut (.A(n1075), .B(det_q4_28[24]), .C(n13016), .Z(n2047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i24_3_lut.init = 16'hcaca;
    LUT4 mux_67_i25_3_lut (.A(n1074), .B(det_q4_28[25]), .C(n13016), .Z(n2046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i25_3_lut.init = 16'hcaca;
    LUT4 mux_67_i26_3_lut (.A(n1073), .B(det_q4_28[26]), .C(n13016), .Z(n2045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i26_3_lut.init = 16'hcaca;
    LUT4 mux_67_i27_3_lut (.A(n1072), .B(det_q4_28[27]), .C(n13016), .Z(n2044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i27_3_lut.init = 16'hcaca;
    LUT4 mux_67_i28_3_lut (.A(n1071), .B(det_q4_28[28]), .C(n13016), .Z(n2043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i28_3_lut.init = 16'hcaca;
    LUT4 mux_67_i29_3_lut (.A(n1070), .B(det_q4_28[29]), .C(n13016), .Z(n2042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i29_3_lut.init = 16'hcaca;
    LUT4 mux_67_i30_3_lut (.A(n1069), .B(det_q4_28[30]), .C(n13016), .Z(n2041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i30_3_lut.init = 16'hcaca;
    LUT4 mux_67_i31_3_lut (.A(n1068), .B(det_q4_28[31]), .C(n13016), .Z(n2040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i31_3_lut.init = 16'hcaca;
    LUT4 mux_67_i6_3_lut (.A(n1093), .B(det_q4_28[6]), .C(n13016), .Z(n2065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_67_i6_3_lut.init = 16'hcaca;
    LUT4 mux_99_i31_3_lut (.A(n1068), .B(det_q4_28[31]), .C(n3077), .Z(n3110[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i31_3_lut.init = 16'hcaca;
    LUT4 i809_2_lut (.A(n1067), .B(n3077), .Z(n3110[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam i809_2_lut.init = 16'h2222;
    LUT4 mux_99_i29_3_lut (.A(n1070), .B(det_q4_28[29]), .C(n3077), .Z(n3110[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i29_3_lut.init = 16'hcaca;
    LUT4 mux_99_i30_3_lut (.A(n1069), .B(det_q4_28[30]), .C(n3077), .Z(n3110[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i30_3_lut.init = 16'hcaca;
    LUT4 mux_99_i27_3_lut (.A(n1072), .B(det_q4_28[27]), .C(n3077), .Z(n3110[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i27_3_lut.init = 16'hcaca;
    LUT4 mux_99_i28_3_lut (.A(n1071), .B(det_q4_28[28]), .C(n3077), .Z(n3110[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i28_3_lut.init = 16'hcaca;
    LUT4 mux_99_i25_3_lut (.A(n1074), .B(det_q4_28[25]), .C(n3077), .Z(n3110[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i25_3_lut.init = 16'hcaca;
    LUT4 mux_99_i26_3_lut (.A(n1073), .B(det_q4_28[26]), .C(n3077), .Z(n3110[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i26_3_lut.init = 16'hcaca;
    LUT4 mux_99_i23_3_lut (.A(n1076), .B(det_q4_28[23]), .C(n3077), .Z(n3110[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i23_3_lut.init = 16'hcaca;
    LUT4 mux_99_i24_3_lut (.A(n1075), .B(det_q4_28[24]), .C(n3077), .Z(n3110[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i24_3_lut.init = 16'hcaca;
    LUT4 mux_99_i21_3_lut (.A(n1078), .B(det_q4_28[21]), .C(n3077), .Z(n3110[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i21_3_lut.init = 16'hcaca;
    LUT4 mux_99_i22_3_lut (.A(n1077), .B(det_q4_28[22]), .C(n3077), .Z(n3110[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i22_3_lut.init = 16'hcaca;
    LUT4 mux_99_i19_3_lut (.A(n1080), .B(det_q4_28[19]), .C(n3077), .Z(n3110[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i19_3_lut.init = 16'hcaca;
    LUT4 mux_99_i20_3_lut (.A(n1079), .B(det_q4_28[20]), .C(n3077), .Z(n3110[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i20_3_lut.init = 16'hcaca;
    LUT4 mux_99_i17_3_lut (.A(n1082), .B(det_q4_28[17]), .C(n3077), .Z(n3110[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i17_3_lut.init = 16'hcaca;
    LUT4 mux_99_i18_3_lut (.A(n1081), .B(det_q4_28[18]), .C(n3077), .Z(n3110[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i18_3_lut.init = 16'hcaca;
    LUT4 mux_99_i15_3_lut (.A(n1084), .B(det_q4_28[15]), .C(n3077), .Z(n3110[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i15_3_lut.init = 16'hcaca;
    LUT4 mux_99_i16_3_lut (.A(n1083), .B(det_q4_28[16]), .C(n3077), .Z(n3110[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i16_3_lut.init = 16'hcaca;
    LUT4 mux_99_i13_3_lut (.A(n1086), .B(det_q4_28[13]), .C(n3077), .Z(n3110[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i13_3_lut.init = 16'hcaca;
    LUT4 mux_99_i14_3_lut (.A(n1085), .B(det_q4_28[14]), .C(n3077), .Z(n3110[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i14_3_lut.init = 16'hcaca;
    LUT4 mux_99_i11_3_lut (.A(n1088), .B(det_q4_28[11]), .C(n3077), .Z(n3110[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i11_3_lut.init = 16'hcaca;
    LUT4 mux_99_i12_3_lut (.A(n1087), .B(det_q4_28[12]), .C(n3077), .Z(n3110[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i12_3_lut.init = 16'hcaca;
    LUT4 mux_99_i9_3_lut (.A(n1090), .B(det_q4_28[9]), .C(n3077), .Z(n3110[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i9_3_lut.init = 16'hcaca;
    LUT4 mux_99_i10_3_lut (.A(n1089), .B(det_q4_28[10]), .C(n3077), .Z(n3110[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i10_3_lut.init = 16'hcaca;
    LUT4 mux_99_i7_3_lut (.A(n1092), .B(det_q4_28[7]), .C(n3077), .Z(n3110[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i7_3_lut.init = 16'hcaca;
    LUT4 mux_99_i8_3_lut (.A(n1091), .B(det_q4_28[8]), .C(n3077), .Z(n3110[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i8_3_lut.init = 16'hcaca;
    LUT4 mux_99_i5_3_lut (.A(n1094), .B(det_q4_28[5]), .C(n3077), .Z(n3110[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i5_3_lut.init = 16'hcaca;
    LUT4 mux_99_i6_3_lut (.A(n1093), .B(det_q4_28[6]), .C(n3077), .Z(n3110[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i6_3_lut.init = 16'hcaca;
    LUT4 mux_99_i3_3_lut (.A(n1096), .B(det_q4_28[3]), .C(n3077), .Z(n3110[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i3_3_lut.init = 16'hcaca;
    LUT4 mux_99_i4_3_lut (.A(n1095), .B(det_q4_28[4]), .C(n3077), .Z(n3110[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i4_3_lut.init = 16'hcaca;
    LUT4 mux_99_i1_3_lut (.A(n1098), .B(det_q4_28[1]), .C(n3077), .Z(n3110[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i1_3_lut.init = 16'hcaca;
    LUT4 mux_99_i2_3_lut (.A(n1097), .B(det_q4_28[2]), .C(n3077), .Z(n3110[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_99_i2_3_lut.init = 16'hcaca;
    LUT4 mux_73_i31_3_lut (.A(n1068), .B(det_q4_28[31]), .C(n13015), .Z(n2241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i31_3_lut.init = 16'hcaca;
    LUT4 mux_73_i29_3_lut (.A(n1070), .B(det_q4_28[29]), .C(n13015), .Z(n2243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i29_3_lut.init = 16'hcaca;
    LUT4 mux_73_i30_3_lut (.A(n1069), .B(det_q4_28[30]), .C(n13015), .Z(n2242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i30_3_lut.init = 16'hcaca;
    LUT4 mux_73_i27_3_lut (.A(n1072), .B(det_q4_28[27]), .C(n13015), .Z(n2245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i27_3_lut.init = 16'hcaca;
    LUT4 mux_73_i28_3_lut (.A(n1071), .B(det_q4_28[28]), .C(n13015), .Z(n2244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i28_3_lut.init = 16'hcaca;
    LUT4 mux_73_i25_3_lut (.A(n1074), .B(det_q4_28[25]), .C(n13015), .Z(n2247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i25_3_lut.init = 16'hcaca;
    LUT4 mux_73_i26_3_lut (.A(n1073), .B(det_q4_28[26]), .C(n13015), .Z(n2246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i26_3_lut.init = 16'hcaca;
    LUT4 mux_73_i23_3_lut (.A(n1076), .B(det_q4_28[23]), .C(n13015), .Z(n2249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i23_3_lut.init = 16'hcaca;
    LUT4 mux_73_i24_3_lut (.A(n1075), .B(det_q4_28[24]), .C(n13015), .Z(n2248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i24_3_lut.init = 16'hcaca;
    LUT4 mux_73_i21_3_lut (.A(n1078), .B(det_q4_28[21]), .C(n13015), .Z(n2251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i21_3_lut.init = 16'hcaca;
    LUT4 mux_73_i22_3_lut (.A(n1077), .B(det_q4_28[22]), .C(n13015), .Z(n2250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i22_3_lut.init = 16'hcaca;
    LUT4 mux_73_i19_3_lut (.A(n1080), .B(det_q4_28[19]), .C(n13015), .Z(n2253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i19_3_lut.init = 16'hcaca;
    LUT4 mux_73_i20_3_lut (.A(n1079), .B(det_q4_28[20]), .C(n13015), .Z(n2252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i20_3_lut.init = 16'hcaca;
    LUT4 mux_73_i17_3_lut (.A(n1082), .B(det_q4_28[17]), .C(n13015), .Z(n2255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i17_3_lut.init = 16'hcaca;
    LUT4 mux_73_i18_3_lut (.A(n1081), .B(det_q4_28[18]), .C(n13015), .Z(n2254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i18_3_lut.init = 16'hcaca;
    LUT4 mux_73_i15_3_lut (.A(n1084), .B(det_q4_28[15]), .C(n13015), .Z(n2257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i15_3_lut.init = 16'hcaca;
    LUT4 mux_73_i16_3_lut (.A(n1083), .B(det_q4_28[16]), .C(n13015), .Z(n2256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i16_3_lut.init = 16'hcaca;
    LUT4 mux_73_i13_3_lut (.A(n1086), .B(det_q4_28[13]), .C(n13015), .Z(n2259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i13_3_lut.init = 16'hcaca;
    LUT4 mux_73_i14_3_lut (.A(n1085), .B(det_q4_28[14]), .C(n13015), .Z(n2258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i14_3_lut.init = 16'hcaca;
    LUT4 mux_73_i11_3_lut (.A(n1088), .B(det_q4_28[11]), .C(n13015), .Z(n2261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i11_3_lut.init = 16'hcaca;
    LUT4 mux_73_i12_3_lut (.A(n1087), .B(det_q4_28[12]), .C(n13015), .Z(n2260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i12_3_lut.init = 16'hcaca;
    LUT4 mux_73_i9_3_lut (.A(n1090), .B(det_q4_28[9]), .C(n13015), .Z(n2263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i9_3_lut.init = 16'hcaca;
    LUT4 mux_73_i10_3_lut (.A(n1089), .B(det_q4_28[10]), .C(n13015), .Z(n2262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i10_3_lut.init = 16'hcaca;
    LUT4 mux_73_i7_3_lut (.A(n1092), .B(det_q4_28[7]), .C(n13015), .Z(n2265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i7_3_lut.init = 16'hcaca;
    LUT4 mux_73_i8_3_lut (.A(n1091), .B(det_q4_28[8]), .C(n13015), .Z(n2264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i8_3_lut.init = 16'hcaca;
    LUT4 mux_73_i5_3_lut (.A(n1094), .B(det_q4_28[5]), .C(n13015), .Z(n2267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i5_3_lut.init = 16'hcaca;
    LUT4 mux_73_i6_3_lut (.A(n1093), .B(det_q4_28[6]), .C(n13015), .Z(n2266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i6_3_lut.init = 16'hcaca;
    LUT4 mux_73_i3_3_lut (.A(n1096), .B(det_q4_28[3]), .C(n13015), .Z(n2269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i3_3_lut.init = 16'hcaca;
    LUT4 mux_73_i4_3_lut (.A(n1095), .B(det_q4_28[4]), .C(n13015), .Z(n2268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i4_3_lut.init = 16'hcaca;
    LUT4 mux_73_i1_3_lut (.A(n1098), .B(det_q4_28[1]), .C(n13015), .Z(n2271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i1_3_lut.init = 16'hcaca;
    LUT4 mux_73_i2_3_lut (.A(n1097), .B(det_q4_28[2]), .C(n13015), .Z(n2270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_73_i2_3_lut.init = 16'hcaca;
    LUT4 mux_97_i1_3_lut (.A(n1098), .B(det_q4_28[1]), .C(n13004), .Z(n3075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i1_3_lut.init = 16'hcaca;
    LUT4 mux_97_i2_3_lut (.A(n1097), .B(det_q4_28[2]), .C(n13004), .Z(n3074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i2_3_lut.init = 16'hcaca;
    LUT4 mux_97_i3_3_lut (.A(n1096), .B(det_q4_28[3]), .C(n13004), .Z(n3073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i3_3_lut.init = 16'hcaca;
    LUT4 mux_97_i4_3_lut (.A(n1095), .B(det_q4_28[4]), .C(n13004), .Z(n3072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i4_3_lut.init = 16'hcaca;
    LUT4 mux_97_i5_3_lut (.A(n1094), .B(det_q4_28[5]), .C(n13004), .Z(n3071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i5_3_lut.init = 16'hcaca;
    LUT4 mux_97_i6_3_lut (.A(n1093), .B(det_q4_28[6]), .C(n13004), .Z(n3070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i6_3_lut.init = 16'hcaca;
    LUT4 mux_97_i7_3_lut (.A(n1092), .B(det_q4_28[7]), .C(n13004), .Z(n3069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i7_3_lut.init = 16'hcaca;
    LUT4 mux_97_i8_3_lut (.A(n1091), .B(det_q4_28[8]), .C(n13004), .Z(n3068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i8_3_lut.init = 16'hcaca;
    LUT4 mux_97_i9_3_lut (.A(n1090), .B(det_q4_28[9]), .C(n13004), .Z(n3067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i9_3_lut.init = 16'hcaca;
    LUT4 mux_97_i10_3_lut (.A(n1089), .B(det_q4_28[10]), .C(n13004), .Z(n3066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i10_3_lut.init = 16'hcaca;
    LUT4 mux_97_i11_3_lut (.A(n1088), .B(det_q4_28[11]), .C(n13004), .Z(n3065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i11_3_lut.init = 16'hcaca;
    LUT4 mux_97_i12_3_lut (.A(n1087), .B(det_q4_28[12]), .C(n13004), .Z(n3064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i12_3_lut.init = 16'hcaca;
    LUT4 mux_97_i13_3_lut (.A(n1086), .B(det_q4_28[13]), .C(n13004), .Z(n3063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i13_3_lut.init = 16'hcaca;
    LUT4 mux_97_i14_3_lut (.A(n1085), .B(det_q4_28[14]), .C(n13004), .Z(n3062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i14_3_lut.init = 16'hcaca;
    LUT4 mux_97_i15_3_lut (.A(n1084), .B(det_q4_28[15]), .C(n13004), .Z(n3061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i15_3_lut.init = 16'hcaca;
    LUT4 mux_97_i16_3_lut (.A(n1083), .B(det_q4_28[16]), .C(n13004), .Z(n3060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i16_3_lut.init = 16'hcaca;
    LUT4 mux_97_i17_3_lut (.A(n1082), .B(det_q4_28[17]), .C(n13004), .Z(n3059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i17_3_lut.init = 16'hcaca;
    LUT4 mux_97_i18_3_lut (.A(n1081), .B(det_q4_28[18]), .C(n13004), .Z(n3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i18_3_lut.init = 16'hcaca;
    LUT4 mux_97_i19_3_lut (.A(n1080), .B(det_q4_28[19]), .C(n13004), .Z(n3057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i19_3_lut.init = 16'hcaca;
    LUT4 mux_97_i20_3_lut (.A(n1079), .B(det_q4_28[20]), .C(n13004), .Z(n3056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i20_3_lut.init = 16'hcaca;
    LUT4 mux_97_i21_3_lut (.A(n1078), .B(det_q4_28[21]), .C(n13004), .Z(n3055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i21_3_lut.init = 16'hcaca;
    LUT4 mux_97_i22_3_lut (.A(n1077), .B(det_q4_28[22]), .C(n13004), .Z(n3054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i22_3_lut.init = 16'hcaca;
    LUT4 mux_97_i23_3_lut (.A(n1076), .B(det_q4_28[23]), .C(n13004), .Z(n3053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i23_3_lut.init = 16'hcaca;
    LUT4 mux_97_i24_3_lut (.A(n1075), .B(det_q4_28[24]), .C(n13004), .Z(n3052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i24_3_lut.init = 16'hcaca;
    LUT4 mux_97_i25_3_lut (.A(n1074), .B(det_q4_28[25]), .C(n13004), .Z(n3051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i25_3_lut.init = 16'hcaca;
    LUT4 mux_97_i26_3_lut (.A(n1073), .B(det_q4_28[26]), .C(n13004), .Z(n3050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i26_3_lut.init = 16'hcaca;
    LUT4 mux_97_i27_3_lut (.A(n1072), .B(det_q4_28[27]), .C(n13004), .Z(n3049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i27_3_lut.init = 16'hcaca;
    LUT4 mux_97_i28_3_lut (.A(n1071), .B(det_q4_28[28]), .C(n13004), .Z(n3048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i28_3_lut.init = 16'hcaca;
    LUT4 i1386_2_lut (.A(n1536), .B(det_zero), .Z(n39)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1386_2_lut.init = 16'h1111;
    LUT4 i1449_4_lut (.A(n68), .B(det_zero), .C(n68_adj_1), .D(n68_adj_2), 
         .Z(n64)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+(C (D))))) */ ;
    defparam i1449_4_lut.init = 16'h0311;
    LUT4 i1422_2_lut (.A(n68_adj_2), .B(det_zero), .Z(n63)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1422_2_lut.init = 16'h1111;
    LUT4 i1425_2_lut (.A(n3077), .B(det_zero), .Z(n62)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1425_2_lut.init = 16'h1111;
    LUT4 mux_97_i29_3_lut (.A(n1070), .B(det_q4_28[29]), .C(n13004), .Z(n3047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i29_3_lut.init = 16'hcaca;
    LUT4 mux_97_i30_3_lut (.A(n1069), .B(det_q4_28[30]), .C(n13004), .Z(n3046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i30_3_lut.init = 16'hcaca;
    LUT4 mux_97_i31_3_lut (.A(n1068), .B(det_q4_28[31]), .C(n13004), .Z(n3045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_97_i31_3_lut.init = 16'hcaca;
    LUT4 mux_51_i1_3_lut (.A(n1098), .B(det_q4_28[1]), .C(n13023), .Z(n1534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i1_3_lut.init = 16'hcaca;
    LUT4 mux_51_i2_3_lut (.A(n1097), .B(det_q4_28[2]), .C(n13023), .Z(n1533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i2_3_lut.init = 16'hcaca;
    LUT4 mux_51_i3_3_lut (.A(n1096), .B(det_q4_28[3]), .C(n13023), .Z(n1532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i3_3_lut.init = 16'hcaca;
    LUT4 mux_51_i4_3_lut (.A(n1095), .B(det_q4_28[4]), .C(n13023), .Z(n1531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i4_3_lut.init = 16'hcaca;
    LUT4 mux_51_i5_3_lut (.A(n1094), .B(det_q4_28[5]), .C(n13023), .Z(n1530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i5_3_lut.init = 16'hcaca;
    LUT4 mux_51_i6_3_lut (.A(n1093), .B(det_q4_28[6]), .C(n13023), .Z(n1529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i6_3_lut.init = 16'hcaca;
    LUT4 mux_51_i7_3_lut (.A(n1092), .B(det_q4_28[7]), .C(n13023), .Z(n1528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i7_3_lut.init = 16'hcaca;
    LUT4 mux_51_i8_3_lut (.A(n1091), .B(det_q4_28[8]), .C(n13023), .Z(n1527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i8_3_lut.init = 16'hcaca;
    LUT4 mux_51_i9_3_lut (.A(n1090), .B(det_q4_28[9]), .C(n13023), .Z(n1526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i9_3_lut.init = 16'hcaca;
    LUT4 mux_51_i10_3_lut (.A(n1089), .B(det_q4_28[10]), .C(n13023), .Z(n1525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i10_3_lut.init = 16'hcaca;
    LUT4 mux_51_i11_3_lut (.A(n1088), .B(det_q4_28[11]), .C(n13023), .Z(n1524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i11_3_lut.init = 16'hcaca;
    LUT4 mux_51_i12_3_lut (.A(n1087), .B(det_q4_28[12]), .C(n13023), .Z(n1523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i12_3_lut.init = 16'hcaca;
    LUT4 mux_51_i13_3_lut (.A(n1086), .B(det_q4_28[13]), .C(n13023), .Z(n1522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i13_3_lut.init = 16'hcaca;
    LUT4 mux_51_i14_3_lut (.A(n1085), .B(det_q4_28[14]), .C(n13023), .Z(n1521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i14_3_lut.init = 16'hcaca;
    LUT4 i1419_2_lut (.A(n2273), .B(det_zero), .Z(n50)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1419_2_lut.init = 16'h1111;
    LUT4 i1383_2_lut (.A(n2139), .B(det_zero), .Z(n48)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1383_2_lut.init = 16'h1111;
    LUT4 i1410_2_lut (.A(n2072), .B(det_zero), .Z(n47)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1410_2_lut.init = 16'h1111;
    CCU2C equal_1287_32 (.A0(det_q4_28[11]), .B0(det_q4_28[16]), .C0(det_q4_28[21]), 
          .D0(det_q4_28[24]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12843), .S1(det_zero));
    defparam equal_1287_32.INIT0 = 16'h0001;
    defparam equal_1287_32.INIT1 = 16'h0000;
    defparam equal_1287_32.INJECT1_0 = "YES";
    defparam equal_1287_32.INJECT1_1 = "NO";
    LUT4 mux_51_i15_3_lut (.A(n1084), .B(det_q4_28[15]), .C(n13023), .Z(n1520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i15_3_lut.init = 16'hcaca;
    CCU2C equal_1287_31 (.A0(det_q4_28[6]), .B0(det_q4_28[31]), .C0(det_q4_28[17]), 
          .D0(det_q4_28[1]), .A1(det_q4_28[4]), .B1(det_q4_28[9]), .C1(det_q4_28[26]), 
          .D1(det_q4_28[12]), .CIN(n12842), .COUT(n12843));
    defparam equal_1287_31.INIT0 = 16'h0001;
    defparam equal_1287_31.INIT1 = 16'h0001;
    defparam equal_1287_31.INJECT1_0 = "YES";
    defparam equal_1287_31.INJECT1_1 = "YES";
    LUT4 mux_51_i16_3_lut (.A(n1083), .B(det_q4_28[16]), .C(n13023), .Z(n1519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i16_3_lut.init = 16'hcaca;
    CCU2C equal_1287_29 (.A0(det_q4_28[15]), .B0(det_q4_28[20]), .C0(det_q4_28[5]), 
          .D0(det_q4_28[22]), .A1(det_q4_28[14]), .B1(det_q4_28[3]), .C1(det_q4_28[13]), 
          .D1(det_q4_28[23]), .CIN(n12841), .COUT(n12842));
    defparam equal_1287_29.INIT0 = 16'h0001;
    defparam equal_1287_29.INIT1 = 16'h0001;
    defparam equal_1287_29.INJECT1_0 = "YES";
    defparam equal_1287_29.INJECT1_1 = "YES";
    LUT4 mux_51_i17_3_lut (.A(n1082), .B(det_q4_28[17]), .C(n13023), .Z(n1518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam mux_51_i17_3_lut.init = 16'hcaca;
    CCU2C equal_1287_27 (.A0(det_q4_28[18]), .B0(det_q4_28[28]), .C0(det_q4_28[2]), 
          .D0(det_q4_28[10]), .A1(det_q4_28[19]), .B1(det_q4_28[7]), .C1(det_q4_28[30]), 
          .D1(det_q4_28[29]), .CIN(n12840), .COUT(n12841));
    defparam equal_1287_27.INIT0 = 16'h0001;
    defparam equal_1287_27.INIT1 = 16'h0001;
    defparam equal_1287_27.INJECT1_0 = "YES";
    defparam equal_1287_27.INJECT1_1 = "YES";
    CCU2C equal_1287_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(det_q4_28[0]), .B1(det_q4_28[27]), .C1(det_q4_28[25]), .D1(det_q4_28[8]), 
          .COUT(n12840));   // d:/rtl_fpga/projeto_final/inverter/reciprocal_q16_16.v(29[24:39])
    defparam equal_1287_0.INIT0 = 16'h000F;
    defparam equal_1287_0.INIT1 = 16'h0001;
    defparam equal_1287_0.INJECT1_0 = "NO";
    defparam equal_1287_0.INJECT1_1 = "YES";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

